module biu32_axi(rstn, clk, write_req, write_ack, write_data, write_sz, write_msk
		, read_req, read_ack, read_data, read_sz, Daddr, code_req, code_ack
		, code_data, code_addr, code_wreq, code_wack, code_wdata, readio_req
		, writeio_req, readio_ack, writeio_ack, writeio_data, readio_data
		, io_add, axi_AW, axi_AWVALID, axi_AWREADY, axi_AWBURST, axi_AWLEN
		, axi_AWSIZE, axi_W, axi_WVALID, axi_WREADY, axi_WSTRB, axi_WLAST
		, axi_AR, axi_ARVALID, axi_ARREADY, axi_ARBURST, axi_ARLEN, axi_ARSIZE
		, axi_R, axi_RVALID, axi_RREADY, axi_RLAST, axi_io_AW, axi_io_AWVALID
		, axi_io_AWREADY, axi_io_AWBURST, axi_io_AWLEN, axi_io_AWSIZE, axi_io_W
		, axi_io_WVALID, axi_io_WREADY, axi_io_WSTRB, axi_io_WLAST, axi_io_AR
		, axi_io_ARVALID, axi_io_ARREADY, axi_io_ARBURST, axi_io_ARLEN, axi_io_ARSIZE
		, axi_io_R, axi_io_RVALID, axi_io_RREADY, axi_io_RLAST, busy, outstanding
		);

	input rstn;
	input clk;
	input write_req;
	output write_ack;
	input [31:0] write_data;
	input [1:0] write_sz;
	input [3:0] write_msk;
	input read_req;
	output read_ack;
	output [31:0] read_data;
	input [1:0] read_sz;
	input [31:0] Daddr;
	input code_req;
	output code_ack;
	output [127:0] code_data;
	input [31:0] code_addr;
	input code_wreq;
	output code_wack;
	input [31:0] code_wdata;
	input readio_req;
	input writeio_req;
	output readio_ack;
	output writeio_ack;
	input [31:0] writeio_data;
	output [31:0] readio_data;
	input [31:0] io_add;
	output [31:0] axi_AW;
	output axi_AWVALID;
	input axi_AWREADY;
	output [1:0] axi_AWBURST;
	output [7:0] axi_AWLEN;
	output [2:0] axi_AWSIZE;
	output [31:0] axi_W;
	output axi_WVALID;
	input axi_WREADY;
	output [3:0] axi_WSTRB;
	output axi_WLAST;
	output [31:0] axi_AR;
	output axi_ARVALID;
	input axi_ARREADY;
	output [1:0] axi_ARBURST;
	output [7:0] axi_ARLEN;
	output [2:0] axi_ARSIZE;
	input [31:0] axi_R;
	input axi_RVALID;
	output axi_RREADY;
	input axi_RLAST;
	output [31:0] axi_io_AW;
	output axi_io_AWVALID;
	input axi_io_AWREADY;
	output [1:0] axi_io_AWBURST;
	output [7:0] axi_io_AWLEN;
	output [2:0] axi_io_AWSIZE;
	output [31:0] axi_io_W;
	output axi_io_WVALID;
	input axi_io_WREADY;
	output [3:0] axi_io_WSTRB;
	output axi_io_WLAST;
	output [31:0] axi_io_AR;
	output axi_io_ARVALID;
	input axi_io_ARREADY;
	output [1:0] axi_io_ARBURST;
	output [7:0] axi_io_ARLEN;
	output [2:0] axi_io_ARSIZE;
	input [31:0] axi_io_R;
	input axi_io_RVALID;
	output axi_io_RREADY;
	input axi_io_RLAST;
	output busy;
	input outstanding;

	wire [1:0] A4;
	wire [4:0] fsm;
	wire [4:0] burst_idx;
	wire [9:0] cacheA;
	wire [149:0] cacheQ;
	wire [149:0] cacheD;
	wire [15:0] cacheM;



	notech_inv i_15188(.A(n_63355), .Z(n_63356));
	notech_inv i_15187(.A(n_63348), .Z(n_63355));
	notech_inv i_15186(.A(n_63353), .Z(n_63354));
	notech_inv i_15185(.A(n_63340), .Z(n_63353));
	notech_inv i_15184(.A(n_63351), .Z(n_63352));
	notech_inv i_15183(.A(n_63336), .Z(n_63351));
	notech_inv i_15182(.A(n_63349), .Z(n_63350));
	notech_inv i_15181(.A(n_63334), .Z(n_63349));
	notech_inv i_15180(.A(n_63347), .Z(n_63348));
	notech_inv i_15179(.A(n_63332), .Z(n_63347));
	notech_inv i_15178(.A(n_63345), .Z(n_63346));
	notech_inv i_15177(.A(n_63324), .Z(n_63345));
	notech_inv i_15176(.A(n_63343), .Z(n_63344));
	notech_inv i_15175(.A(n_63322), .Z(n_63343));
	notech_inv i_15174(.A(n_63341), .Z(n_63342));
	notech_inv i_15173(.A(n_63320), .Z(n_63341));
	notech_inv i_15172(.A(n_63339), .Z(n_63340));
	notech_inv i_15171(.A(n_63318), .Z(n_63339));
	notech_inv i_15170(.A(n_63337), .Z(n_63338));
	notech_inv i_15169(.A(n_63316), .Z(n_63337));
	notech_inv i_15168(.A(n_63335), .Z(n_63336));
	notech_inv i_15167(.A(n_63314), .Z(n_63335));
	notech_inv i_15166(.A(n_63333), .Z(n_63334));
	notech_inv i_15165(.A(n_63312), .Z(n_63333));
	notech_inv i_15164(.A(n_63331), .Z(n_63332));
	notech_inv i_15163(.A(n_63350), .Z(n_63331));
	notech_inv i_15162(.A(n_63329), .Z(n_63330));
	notech_inv i_15161(.A(n_63306), .Z(n_63329));
	notech_inv i_15160(.A(n_63327), .Z(n_63328));
	notech_inv i_15159(.A(n_63302), .Z(n_63327));
	notech_inv i_15158(.A(n_63325), .Z(n_63326));
	notech_inv i_15157(.A(n_63300), .Z(n_63325));
	notech_inv i_15156(.A(n_63323), .Z(n_63324));
	notech_inv i_15155(.A(n_63326), .Z(n_63323));
	notech_inv i_15154(.A(n_63321), .Z(n_63322));
	notech_inv i_15153(.A(n_63296), .Z(n_63321));
	notech_inv i_15152(.A(n_63319), .Z(n_63320));
	notech_inv i_15151(.A(n_63294), .Z(n_63319));
	notech_inv i_15150(.A(n_63317), .Z(n_63318));
	notech_inv i_15149(.A(n_63342), .Z(n_63317));
	notech_inv i_15148(.A(n_63315), .Z(n_63316));
	notech_inv i_15147(.A(n_63292), .Z(n_63315));
	notech_inv i_15146(.A(n_63313), .Z(n_63314));
	notech_inv i_15145(.A(n_63338), .Z(n_63313));
	notech_inv i_15144(.A(n_63311), .Z(n_63312));
	notech_inv i_15143(.A(n_63352), .Z(n_63311));
	notech_inv i_15142(.A(n_63309), .Z(n_63310));
	notech_inv i_15141(.A(n_63288), .Z(n_63309));
	notech_inv i_15140(.A(n_63307), .Z(n_63308));
	notech_inv i_15139(.A(n_63286), .Z(n_63307));
	notech_inv i_15138(.A(n_63305), .Z(n_63306));
	notech_inv i_15137(.A(n_63308), .Z(n_63305));
	notech_inv i_15136(.A(n_63303), .Z(n_63304));
	notech_inv i_15135(.A(n_63284), .Z(n_63303));
	notech_inv i_15134(.A(n_63301), .Z(n_63302));
	notech_inv i_15133(.A(n_63304), .Z(n_63301));
	notech_inv i_15132(.A(n_63299), .Z(n_63300));
	notech_inv i_15131(.A(n_63328), .Z(n_63299));
	notech_inv i_15130(.A(n_63297), .Z(n_63298));
	notech_inv i_15129(.A(n_63282), .Z(n_63297));
	notech_inv i_15128(.A(n_63295), .Z(n_63296));
	notech_inv i_15127(.A(n_63298), .Z(n_63295));
	notech_inv i_15126(.A(n_63293), .Z(n_63294));
	notech_inv i_15125(.A(n_63344), .Z(n_63293));
	notech_inv i_15124(.A(n_63291), .Z(n_63292));
	notech_inv i_15123(.A(n_63354), .Z(n_63291));
	notech_inv i_15122(.A(n_63289), .Z(n_63290));
	notech_inv i_15121(.A(clk), .Z(n_63289));
	notech_inv i_15120(.A(n_63287), .Z(n_63288));
	notech_inv i_15119(.A(n_63290), .Z(n_63287));
	notech_inv i_15118(.A(n_63285), .Z(n_63286));
	notech_inv i_15117(.A(n_63310), .Z(n_63285));
	notech_inv i_15116(.A(n_63283), .Z(n_63284));
	notech_inv i_15115(.A(n_63330), .Z(n_63283));
	notech_inv i_15114(.A(n_63281), .Z(n_63282));
	notech_inv i_15113(.A(n_63346), .Z(n_63281));
	notech_inv i_14669(.A(n_62814), .Z(n_62826));
	notech_inv i_14668(.A(n_62814), .Z(n_62825));
	notech_inv i_14663(.A(n_62814), .Z(n_62820));
	notech_inv i_14658(.A(n_62814), .Z(n_62815));
	notech_inv i_14657(.A(n_2008), .Z(n_62814));
	notech_inv i_14654(.A(n_62798), .Z(n_62810));
	notech_inv i_14653(.A(n_62798), .Z(n_62809));
	notech_inv i_14648(.A(n_62798), .Z(n_62804));
	notech_inv i_14643(.A(n_62798), .Z(n_62799));
	notech_inv i_14642(.A(n_1996), .Z(n_62798));
	notech_inv i_14638(.A(n_62787), .Z(n_62793));
	notech_inv i_14633(.A(n_62787), .Z(n_62788));
	notech_inv i_14632(.A(n_968), .Z(n_62787));
	notech_inv i_14629(.A(n_62771), .Z(n_62783));
	notech_inv i_14628(.A(n_62771), .Z(n_62782));
	notech_inv i_14623(.A(n_62771), .Z(n_62777));
	notech_inv i_14618(.A(n_62771), .Z(n_62772));
	notech_inv i_14617(.A(n_972), .Z(n_62771));
	notech_inv i_14589(.A(n_62733), .Z(n_62739));
	notech_inv i_14584(.A(n_62733), .Z(n_62734));
	notech_inv i_14583(.A(n_2004), .Z(n_62733));
	notech_inv i_14582(.A(n_62711), .Z(n_62731));
	notech_inv i_14581(.A(n_62711), .Z(n_62730));
	notech_inv i_14580(.A(n_62711), .Z(n_62729));
	notech_inv i_14579(.A(n_62711), .Z(n_62728));
	notech_inv i_14578(.A(n_62711), .Z(n_62727));
	notech_inv i_14577(.A(n_62711), .Z(n_62726));
	notech_inv i_14575(.A(n_62711), .Z(n_62724));
	notech_inv i_14574(.A(n_62711), .Z(n_62723));
	notech_inv i_14573(.A(n_62711), .Z(n_62722));
	notech_inv i_14572(.A(n_62711), .Z(n_62721));
	notech_inv i_14571(.A(n_62711), .Z(n_62720));
	notech_inv i_14570(.A(n_62711), .Z(n_62719));
	notech_inv i_14568(.A(n_62711), .Z(n_62717));
	notech_inv i_14567(.A(n_62711), .Z(n_62716));
	notech_inv i_14566(.A(n_62711), .Z(n_62715));
	notech_inv i_14565(.A(n_62711), .Z(n_62714));
	notech_inv i_14564(.A(n_62711), .Z(n_62713));
	notech_inv i_14563(.A(n_62711), .Z(n_62712));
	notech_inv i_14562(.A(rstn), .Z(n_62711));
	notech_inv i_14014(.A(n_62169), .Z(n_62170));
	notech_inv i_14013(.A(n_2033), .Z(n_62169));
	notech_inv i_14006(.A(n_62160), .Z(n_62161));
	notech_inv i_14005(.A(n_2010), .Z(n_62160));
	notech_inv i_13996(.A(n_62149), .Z(n_62150));
	notech_inv i_13995(.A(n_1067), .Z(n_62149));
	notech_inv i_13988(.A(n_62140), .Z(n_62141));
	notech_inv i_13987(.A(n_1061), .Z(n_62140));
	notech_inv i_13980(.A(n_62131), .Z(n_62132));
	notech_inv i_13979(.A(n_2023), .Z(n_62131));
	notech_inv i_13972(.A(n_62122), .Z(n_62123));
	notech_inv i_13971(.A(n_8212), .Z(n_62122));
	notech_inv i_13964(.A(n_62113), .Z(n_62114));
	notech_inv i_13963(.A(n_8233), .Z(n_62113));
	notech_inv i_13956(.A(n_62100), .Z(n_62105));
	notech_inv i_13952(.A(n_62100), .Z(n_62101));
	notech_inv i_13951(.A(\nbus_11662[0] ), .Z(n_62100));
	notech_inv i_13408(.A(n_61571), .Z(n_61573));
	notech_inv i_13407(.A(n_61571), .Z(code_data[0]));
	notech_inv i_13406(.A(\nbus_14547[0] ), .Z(n_61571));
	notech_inv i_12771(.A(n_60808), .Z(n_60809));
	notech_inv i_12770(.A(n_1277), .Z(n_60808));
	notech_inv i_12761(.A(n_60797), .Z(n_60798));
	notech_inv i_12760(.A(n_1375), .Z(n_60797));
	notech_inv i_12753(.A(n_60784), .Z(n_60789));
	notech_inv i_12749(.A(n_60784), .Z(n_60785));
	notech_inv i_12748(.A(A4[1]), .Z(n_60784));
	notech_inv i_12744(.A(n_60765), .Z(n_60779));
	notech_inv i_12743(.A(n_60765), .Z(n_60778));
	notech_inv i_12737(.A(n_60765), .Z(n_60772));
	notech_inv i_12731(.A(n_60765), .Z(n_60766));
	notech_inv i_12730(.A(n_2072), .Z(n_60765));
	notech_inv i_12728(.A(n_60749), .Z(n_60762));
	notech_inv i_12726(.A(n_60749), .Z(n_60760));
	notech_inv i_12722(.A(n_60749), .Z(n_60756));
	notech_inv i_12721(.A(n_60749), .Z(n_60755));
	notech_inv i_12716(.A(n_60749), .Z(n_60750));
	notech_inv i_12715(.A(A4[0]), .Z(n_60749));
	notech_inv i_12711(.A(n_60730), .Z(n_60744));
	notech_inv i_12710(.A(n_60730), .Z(n_60743));
	notech_inv i_12704(.A(n_60730), .Z(n_60737));
	notech_inv i_12698(.A(n_60730), .Z(n_60731));
	notech_inv i_12697(.A(n_2074), .Z(n_60730));
	notech_inv i_12695(.A(n_60755), .Z(n_60727));
	notech_inv i_12693(.A(n_60755), .Z(n_60725));
	notech_inv i_12690(.A(n_60755), .Z(n_60722));
	notech_inv i_12688(.A(n_60755), .Z(n_60720));
	notech_inv i_12685(.A(n_60755), .Z(n_60717));
	notech_inv i_12683(.A(n_60755), .Z(n_60715));
	notech_inv i_12673(.A(n_60703), .Z(n_60704));
	notech_inv i_12672(.A(n_1377), .Z(n_60703));
	notech_inv i_12663(.A(n_60692), .Z(n_60693));
	notech_inv i_12662(.A(n_1474), .Z(n_60692));
	notech_inv i_12653(.A(n_60681), .Z(n_60682));
	notech_inv i_12652(.A(n_1476), .Z(n_60681));
	notech_inv i_12643(.A(n_60670), .Z(n_60671));
	notech_inv i_12642(.A(n_1573), .Z(n_60670));
	notech_inv i_12633(.A(n_60659), .Z(n_60660));
	notech_inv i_12632(.A(n_1575), .Z(n_60659));
	notech_inv i_12623(.A(n_60648), .Z(n_60649));
	notech_inv i_12622(.A(n_1703), .Z(n_60648));
	notech_inv i_12613(.A(n_60637), .Z(n_60638));
	notech_inv i_12612(.A(n_1705), .Z(n_60637));
	notech_inv i_9884(.A(n_57732), .Z(n_57733));
	notech_inv i_9883(.A(\nbus_11667[0] ), .Z(n_57732));
	notech_inv i_8247(.A(n_56051), .Z(n_56052));
	notech_inv i_8246(.A(\nbus_11671[0] ), .Z(n_56051));
	notech_inv i_7933(.A(n_55689), .Z(n_55690));
	notech_inv i_7932(.A(\nbus_11667[96] ), .Z(n_55689));
	notech_inv i_7923(.A(n_55678), .Z(n_55679));
	notech_inv i_7922(.A(\nbus_11667[32] ), .Z(n_55678));
	notech_inv i_7913(.A(n_55667), .Z(n_55668));
	notech_inv i_7912(.A(\nbus_11667[64] ), .Z(n_55667));
	notech_inv i_7774(.A(n_55485), .Z(n_55486));
	notech_inv i_7773(.A(n_2244), .Z(n_55485));
	notech_inv i_7764(.A(n_55474), .Z(n_55475));
	notech_inv i_7763(.A(n_2239), .Z(n_55474));
	notech_inv i_7756(.A(n_55421), .Z(n_55422));
	notech_inv i_7755(.A(n_2237), .Z(n_55421));
	notech_ao4 i_56360(.A(n_1061), .B(n_8394), .C(n_2010), .D(n_8432), .Z(n_986
		));
	notech_ao4 i_56366(.A(n_1061), .B(n_8395), .C(n_2010), .D(n_8433), .Z(n_983
		));
	notech_ao4 i_56372(.A(n_1061), .B(n_8396), .C(n_2010), .D(n_8434), .Z(n_980
		));
	notech_and4 i_57606(.A(n_62825), .B(n_62739), .C(n_973), .D(n_976), .Z(n_977
		));
	notech_nand3 i_151(.A(axi_RVALID), .B(axi_RLAST), .C(n_22714), .Z(n_976)
		);
	notech_ao3 i_58535(.A(n_62782), .B(n_973), .C(n_974), .Z(n_975));
	notech_and2 i_147(.A(axi_WREADY), .B(n_25047), .Z(n_974));
	notech_and2 i_45(.A(n_1215), .B(n_2010), .Z(n_973));
	notech_and3 i_50(.A(n_62825), .B(n_62793), .C(n_8323), .Z(n_972));
	notech_nor2 i_137(.A(code_ack), .B(n_8564), .Z(n_971));
	notech_nor2 i_136(.A(read_ack), .B(n_8565), .Z(n_970));
	notech_nao3 i_64(.A(n_8325), .B(n_8328), .C(n_2000), .Z(busy));
	notech_and2 i_11(.A(n_62809), .B(n_8225), .Z(n_968));
	notech_xor2 i_132(.A(burst_idx[4]), .B(n_2027), .Z(n_967));
	notech_xor2 i_131(.A(burst_idx[3]), .B(n_2026), .Z(n_966));
	notech_xor2 i_130(.A(burst_idx[2]), .B(n_2025), .Z(n_965));
	notech_nand2 i_127(.A(n_1215), .B(n_8323), .Z(n_963));
	notech_xor2 i_1880680(.A(axi_AR[14]), .B(cacheQ[128]), .Z(n_960));
	notech_xor2 i_1980681(.A(axi_AR[15]), .B(cacheQ[129]), .Z(n_959));
	notech_xor2 i_20(.A(axi_AR[16]), .B(cacheQ[130]), .Z(n_958));
	notech_xor2 i_2180682(.A(axi_AR[17]), .B(cacheQ[131]), .Z(n_957));
	notech_xor2 i_2280683(.A(axi_AR[18]), .B(cacheQ[132]), .Z(n_956));
	notech_xor2 i_2380684(.A(axi_AR[19]), .B(cacheQ[133]), .Z(n_955));
	notech_xor2 i_24(.A(axi_AR[20]), .B(cacheQ[134]), .Z(n_954));
	notech_xor2 i_25(.A(axi_AR[21]), .B(cacheQ[135]), .Z(n_953));
	notech_xor2 i_2680685(.A(axi_AR[22]), .B(cacheQ[136]), .Z(n_952));
	notech_xor2 i_2780686(.A(axi_AR[23]), .B(cacheQ[137]), .Z(n_951));
	notech_xor2 i_28(.A(axi_AR[24]), .B(cacheQ[138]), .Z(n_950));
	notech_xor2 i_2980687(.A(axi_AR[25]), .B(cacheQ[139]), .Z(n_949));
	notech_xor2 i_3080688(.A(axi_AR[26]), .B(cacheQ[140]), .Z(n_948));
	notech_xor2 i_3180689(.A(axi_AR[27]), .B(cacheQ[141]), .Z(n_947));
	notech_xor2 i_3280690(.A(axi_AR[28]), .B(cacheQ[142]), .Z(n_946));
	notech_xor2 i_3380691(.A(axi_AR[29]), .B(cacheQ[143]), .Z(n_945));
	notech_xor2 i_3480692(.A(axi_AR[30]), .B(cacheQ[144]), .Z(n_944));
	notech_xor2 i_3580693(.A(axi_AR[31]), .B(cacheQ[145]), .Z(n_943));
	notech_or4 i_4780703(.A(n_960), .B(n_959), .C(n_958), .D(n_957), .Z(n_934
		));
	notech_or4 i_4880704(.A(n_956), .B(n_955), .C(n_954), .D(n_953), .Z(n_933
		));
	notech_or4 i_4980705(.A(n_952), .B(n_951), .C(n_950), .D(n_949), .Z(n_932
		));
	notech_or4 i_5080706(.A(n_948), .B(n_947), .C(n_946), .D(n_945), .Z(n_931
		));
	notech_or4 i_5580709(.A(n_934), .B(n_933), .C(n_932), .D(n_931), .Z(n_928
		));
	notech_xor2 i_1880729(.A(cacheQ[128]), .B(axi_AW[14]), .Z(n_926));
	notech_xor2 i_1980730(.A(cacheQ[129]), .B(axi_AW[15]), .Z(n_925));
	notech_xor2 i_2080731(.A(cacheQ[130]), .B(axi_AW[16]), .Z(n_924));
	notech_xor2 i_2180732(.A(cacheQ[131]), .B(axi_AW[17]), .Z(n_923));
	notech_xor2 i_2280733(.A(cacheQ[132]), .B(axi_AW[18]), .Z(n_922));
	notech_xor2 i_2380734(.A(cacheQ[133]), .B(axi_AW[19]), .Z(n_921));
	notech_xor2 i_2480735(.A(cacheQ[134]), .B(axi_AW[20]), .Z(n_920));
	notech_xor2 i_2580736(.A(cacheQ[135]), .B(axi_AW[21]), .Z(n_919));
	notech_xor2 i_2680737(.A(cacheQ[136]), .B(axi_AW[22]), .Z(n_918));
	notech_xor2 i_2780738(.A(cacheQ[137]), .B(axi_AW[23]), .Z(n_917));
	notech_xor2 i_2880739(.A(cacheQ[138]), .B(axi_AW[24]), .Z(n_916));
	notech_xor2 i_2980740(.A(cacheQ[139]), .B(axi_AW[25]), .Z(n_915));
	notech_xor2 i_3080741(.A(cacheQ[140]), .B(axi_AW[26]), .Z(n_914));
	notech_xor2 i_3180742(.A(cacheQ[141]), .B(axi_AW[27]), .Z(n_913));
	notech_xor2 i_3280743(.A(cacheQ[142]), .B(axi_AW[28]), .Z(n_912));
	notech_xor2 i_3380744(.A(cacheQ[143]), .B(axi_AW[29]), .Z(n_911));
	notech_xor2 i_3480745(.A(n_8555), .B(axi_AW[30]), .Z(n_910));
	notech_xor2 i_3580746(.A(n_8556), .B(axi_AW[31]), .Z(n_909));
	notech_or4 i_4780756(.A(n_926), .B(n_925), .C(n_924), .D(n_923), .Z(n_900
		));
	notech_or4 i_4880757(.A(n_922), .B(n_921), .C(n_920), .D(n_919), .Z(n_899
		));
	notech_or4 i_4980758(.A(n_918), .B(n_917), .C(n_916), .D(n_915), .Z(n_898
		));
	notech_or4 i_5080759(.A(n_914), .B(n_913), .C(n_912), .D(n_911), .Z(n_897
		));
	notech_or4 i_5580762(.A(n_900), .B(n_899), .C(n_898), .D(n_897), .Z(n_894
		));
	notech_ao4 i_56354(.A(n_1061), .B(n_8393), .C(n_2010), .D(n_8431), .Z(n_989
		));
	notech_ao4 i_56348(.A(n_1061), .B(n_8392), .C(n_2010), .D(n_8430), .Z(n_992
		));
	notech_ao4 i_56342(.A(n_1061), .B(n_8391), .C(n_2010), .D(n_8429), .Z(n_995
		));
	notech_ao4 i_56336(.A(n_1061), .B(n_8390), .C(n_2010), .D(n_8428), .Z(n_998
		));
	notech_ao4 i_56330(.A(n_1061), .B(n_8389), .C(n_2010), .D(n_8427), .Z(n_1001
		));
	notech_ao4 i_56324(.A(n_1061), .B(n_8388), .C(n_2010), .D(n_8426), .Z(n_1004
		));
	notech_ao4 i_56318(.A(n_1061), .B(n_8387), .C(n_2010), .D(n_8425), .Z(n_1007
		));
	notech_ao4 i_56312(.A(n_1061), .B(n_8386), .C(n_2010), .D(n_8424), .Z(n_1010
		));
	notech_ao4 i_56306(.A(n_1061), .B(n_8385), .C(n_2010), .D(n_8423), .Z(n_1013
		));
	notech_ao4 i_56300(.A(n_1061), .B(n_8384), .C(n_2010), .D(n_8422), .Z(n_1016
		));
	notech_ao4 i_56294(.A(n_1061), .B(n_8383), .C(n_2010), .D(n_8421), .Z(n_1019
		));
	notech_ao4 i_56288(.A(n_62141), .B(n_8382), .C(n_2010), .D(n_8420), .Z(n_1022
		));
	notech_ao4 i_56282(.A(n_62141), .B(n_8381), .C(n_2010), .D(n_8419), .Z(n_1025
		));
	notech_ao4 i_56276(.A(n_62141), .B(n_8380), .C(n_2010), .D(n_8418), .Z(n_1028
		));
	notech_ao4 i_56270(.A(n_62141), .B(n_8379), .C(n_62161), .D(n_8417), .Z(n_1031
		));
	notech_ao4 i_56264(.A(n_62141), .B(n_8369), .C(n_62161), .D(n_8416), .Z(n_1034
		));
	notech_ao4 i_56258(.A(n_62141), .B(n_8370), .C(n_62161), .D(n_8415), .Z(n_1037
		));
	notech_ao4 i_56252(.A(n_62141), .B(n_8371), .C(n_62161), .D(n_8414), .Z(n_1040
		));
	notech_ao4 i_56246(.A(n_62141), .B(n_8372), .C(n_62161), .D(n_8413), .Z(n_1043
		));
	notech_ao4 i_56240(.A(n_62141), .B(n_8373), .C(n_62161), .D(n_8412), .Z(n_1046
		));
	notech_ao4 i_56234(.A(n_1061), .B(n_8374), .C(n_62161), .D(n_8411), .Z(n_1049
		));
	notech_ao4 i_56228(.A(n_62141), .B(n_8375), .C(n_62161), .D(n_8410), .Z(n_1052
		));
	notech_ao4 i_56222(.A(n_62141), .B(n_8376), .C(n_62161), .D(n_8409), .Z(n_1055
		));
	notech_ao4 i_56216(.A(n_62141), .B(n_8377), .C(n_62161), .D(n_8408), .Z(n_1058
		));
	notech_and3 i_32(.A(n_2019), .B(n_1215), .C(n_62793), .Z(n_1061));
	notech_ao4 i_56210(.A(n_62141), .B(n_8378), .C(n_62161), .D(n_8407), .Z(n_1062
		));
	notech_ao4 i_56204(.A(n_2020), .B(n_8368), .C(n_62161), .D(n_8406), .Z(n_1065
		));
	notech_nao3 i_242(.A(axi_AR[30]), .B(n_8559), .C(n_2019), .Z(n_1066));
	notech_and4 i_58465(.A(n_1215), .B(n_62161), .C(n_1066), .D(n_62793), .Z
		(n_1067));
	notech_ao4 i_56199(.A(n_2020), .B(n_8367), .C(n_62161), .D(n_8405), .Z(n_1070
		));
	notech_ao4 i_56523(.A(n_62825), .B(n_8434), .C(n_62739), .D(n_8396), .Z(n_1073
		));
	notech_ao4 i_56518(.A(n_62825), .B(n_8433), .C(n_62739), .D(n_8395), .Z(n_1076
		));
	notech_ao4 i_56513(.A(n_62825), .B(n_8432), .C(n_62739), .D(n_8394), .Z(n_1079
		));
	notech_ao4 i_56508(.A(n_62825), .B(n_8431), .C(n_62739), .D(n_8393), .Z(n_1082
		));
	notech_ao4 i_56503(.A(n_62825), .B(n_8430), .C(n_62739), .D(n_8392), .Z(n_1085
		));
	notech_ao4 i_56498(.A(n_62825), .B(n_8429), .C(n_62739), .D(n_8391), .Z(n_1088
		));
	notech_ao4 i_56493(.A(n_62825), .B(n_8428), .C(n_62739), .D(n_8390), .Z(n_1091
		));
	notech_ao4 i_56488(.A(n_62825), .B(n_8427), .C(n_62739), .D(n_8389), .Z(n_1094
		));
	notech_ao4 i_56483(.A(n_62825), .B(n_8426), .C(n_62739), .D(n_8388), .Z(n_1097
		));
	notech_ao4 i_56478(.A(n_62825), .B(n_8425), .C(n_62739), .D(n_8387), .Z(n_1100
		));
	notech_ao4 i_56473(.A(n_62825), .B(n_8424), .C(n_62739), .D(n_8386), .Z(n_1103
		));
	notech_ao4 i_56468(.A(n_62825), .B(n_8423), .C(n_62739), .D(n_8385), .Z(n_1106
		));
	notech_ao4 i_56463(.A(n_62825), .B(n_8422), .C(n_62739), .D(n_8384), .Z(n_1109
		));
	notech_ao4 i_56458(.A(n_62825), .B(n_8421), .C(n_62739), .D(n_8383), .Z(n_1112
		));
	notech_ao4 i_56453(.A(n_62825), .B(n_8420), .C(n_62739), .D(n_8382), .Z(n_1115
		));
	notech_ao4 i_56448(.A(n_62825), .B(n_8419), .C(n_62739), .D(n_8381), .Z(n_1118
		));
	notech_ao4 i_56443(.A(n_62826), .B(n_8418), .C(n_62739), .D(n_8380), .Z(n_1121
		));
	notech_ao4 i_56438(.A(n_62826), .B(n_8417), .C(n_62739), .D(n_8379), .Z(n_1124
		));
	notech_ao4 i_56433(.A(n_62826), .B(n_8416), .C(n_62739), .D(n_8369), .Z(n_1127
		));
	notech_ao4 i_56428(.A(n_62826), .B(n_8415), .C(n_62734), .D(n_8370), .Z(n_1130
		));
	notech_ao4 i_56423(.A(n_62826), .B(n_8414), .C(n_62734), .D(n_8371), .Z(n_1133
		));
	notech_ao4 i_56418(.A(n_62826), .B(n_8413), .C(n_62734), .D(n_8372), .Z(n_1136
		));
	notech_ao4 i_56413(.A(n_62826), .B(n_8412), .C(n_62734), .D(n_8373), .Z(n_1139
		));
	notech_ao4 i_56408(.A(n_62826), .B(n_8411), .C(n_62734), .D(n_8374), .Z(n_1142
		));
	notech_ao4 i_56403(.A(n_62826), .B(n_8410), .C(n_62734), .D(n_8375), .Z(n_1145
		));
	notech_ao4 i_56398(.A(n_62826), .B(n_8409), .C(n_62734), .D(n_8376), .Z(n_1148
		));
	notech_ao4 i_56393(.A(n_62826), .B(n_8408), .C(n_62734), .D(n_8377), .Z(n_1151
		));
	notech_ao4 i_56388(.A(n_62826), .B(n_8407), .C(n_62734), .D(n_8378), .Z(n_1154
		));
	notech_ao4 i_56383(.A(n_62826), .B(n_8406), .C(n_62734), .D(n_8368), .Z(n_1157
		));
	notech_ao4 i_56378(.A(n_62826), .B(n_8405), .C(n_62734), .D(n_8367), .Z(n_1160
		));
	notech_nao3 i_348(.A(n_2033), .B(n_2035), .C(n_2040), .Z(n_1167));
	notech_and3 i_126(.A(n_8323), .B(n_973), .C(n_1167), .Z(n_1170));
	notech_ao4 i_58840(.A(n_1170), .B(n_8561), .C(n_2024), .D(n_2030), .Z(n_1171
		));
	notech_ao4 i_56528(.A(n_2024), .B(burst_idx[0]), .C(n_2032), .D(n_2000),
		 .Z(n_1173));
	notech_nand2 i_354(.A(axi_AWREADY), .B(n_8229), .Z(n_1174));
	notech_and4 i_57260(.A(n_62826), .B(n_62793), .C(n_8323), .D(n_1174), .Z
		(n_1175));
	notech_nand2 i_105(.A(n_62826), .B(n_8323), .Z(n_1176));
	notech_ao4 i_56592(.A(n_62826), .B(n_8404), .C(n_62734), .D(n_8442), .Z(n_1179
		));
	notech_ao4 i_56587(.A(n_62826), .B(n_8403), .C(n_62734), .D(n_8441), .Z(n_1182
		));
	notech_ao4 i_56582(.A(n_62815), .B(n_8402), .C(n_62734), .D(n_8440), .Z(n_1185
		));
	notech_ao4 i_56577(.A(n_62815), .B(n_8401), .C(n_62734), .D(n_8439), .Z(n_1188
		));
	notech_ao4 i_56572(.A(n_62815), .B(n_8400), .C(n_62734), .D(n_8438), .Z(n_1191
		));
	notech_ao4 i_56567(.A(n_62815), .B(n_8399), .C(n_62734), .D(n_8437), .Z(n_1194
		));
	notech_ao4 i_56562(.A(n_62815), .B(n_8398), .C(n_62734), .D(n_8436), .Z(n_1197
		));
	notech_ao4 i_56557(.A(n_62815), .B(n_8397), .C(n_62734), .D(n_8435), .Z(n_1200
		));
	notech_and4 i_59007(.A(n_2046), .B(n_62793), .C(n_8323), .D(n_973), .Z(n_1203
		));
	notech_nand2 i_56691(.A(n_2045), .B(n_8265), .Z(n_1204));
	notech_or2 i_389(.A(n_1995), .B(n_2017), .Z(n_1205));
	notech_nao3 i_391(.A(read_req), .B(n_2052), .C(n_2045), .Z(n_1207));
	notech_and4 i_57897(.A(n_62782), .B(n_2051), .C(n_973), .D(n_1207), .Z(n_1208
		));
	notech_or2 i_396(.A(abort), .B(n_2045), .Z(n_1209));
	notech_nand3 i_56694(.A(n_2019), .B(n_1205), .C(n_1209), .Z(n_1210));
	notech_ao3 i_57851(.A(n_62782), .B(n_973), .C(n_2033), .Z(n_1211));
	notech_nand3 i_56706(.A(n_62161), .B(n_2058), .C(n_62815), .Z(n_1212));
	notech_and4 i_56704(.A(n_2061), .B(n_62815), .C(n_2024), .D(n_2056), .Z(n_1213
		));
	notech_nand2 i_56703(.A(n_1066), .B(n_2058), .Z(n_1214));
	notech_or4 i_60(.A(read_ack), .B(n_2003), .C(busy), .D(n_8565), .Z(n_1215
		));
	notech_nao3 i_56701(.A(n_1215), .B(n_2058), .C(n_1221), .Z(n_1216));
	notech_nand2 i_410(.A(axi_WREADY), .B(n_8229), .Z(n_1217));
	notech_and4 i_57881(.A(n_62815), .B(n_1217), .C(n_62793), .D(n_8323), .Z
		(n_1218));
	notech_ao3 i_61(.A(fsm[3]), .B(fsm[0]), .C(n_2000), .Z(n_1221));
	notech_and4 i_58067(.A(n_62782), .B(n_2064), .C(n_2066), .D(n_1217), .Z(n_1222
		));
	notech_and4 i_56699(.A(n_2024), .B(n_8323), .C(n_2057), .D(n_973), .Z(n_1223
		));
	notech_nand2 i_57175(.A(n_8212), .B(n_8221), .Z(n_1224));
	notech_ao4 i_57169(.A(n_8212), .B(n_8396), .C(n_8556), .D(n_8221), .Z(n_1227
		));
	notech_ao4 i_57166(.A(n_8212), .B(n_8395), .C(n_8555), .D(n_8221), .Z(n_1230
		));
	notech_ao4 i_57163(.A(n_8212), .B(n_8394), .C(n_8221), .D(n_8554), .Z(n_1233
		));
	notech_ao4 i_57160(.A(n_8212), .B(n_8393), .C(n_8221), .D(n_8553), .Z(n_1236
		));
	notech_ao4 i_57157(.A(n_8212), .B(n_8392), .C(n_8221), .D(n_8552), .Z(n_1239
		));
	notech_ao4 i_57154(.A(n_8212), .B(n_8391), .C(n_8221), .D(n_8551), .Z(n_1242
		));
	notech_ao4 i_57151(.A(n_8212), .B(n_8390), .C(n_8221), .D(n_8550), .Z(n_1245
		));
	notech_ao4 i_57148(.A(n_8212), .B(n_8389), .C(n_8221), .D(n_8549), .Z(n_1248
		));
	notech_ao4 i_57145(.A(n_8212), .B(n_8388), .C(n_8221), .D(n_8548), .Z(n_1251
		));
	notech_ao4 i_57142(.A(n_8212), .B(n_8387), .C(n_8221), .D(n_8547), .Z(n_1254
		));
	notech_ao4 i_57139(.A(n_8212), .B(n_8386), .C(n_8221), .D(n_8546), .Z(n_1257
		));
	notech_ao4 i_57136(.A(n_62123), .B(n_8385), .C(n_8221), .D(n_8545), .Z(n_1260
		));
	notech_ao4 i_57133(.A(n_62123), .B(n_8384), .C(n_8221), .D(n_8544), .Z(n_1263
		));
	notech_ao4 i_57130(.A(n_62123), .B(n_8383), .C(n_8221), .D(n_8543), .Z(n_1266
		));
	notech_ao4 i_57127(.A(n_62123), .B(n_8382), .C(n_8221), .D(n_8542), .Z(n_1269
		));
	notech_ao4 i_57124(.A(n_62123), .B(n_8381), .C(n_8221), .D(n_8541), .Z(n_1272
		));
	notech_ao4 i_57121(.A(n_62123), .B(n_8380), .C(n_8221), .D(n_8540), .Z(n_1275
		));
	notech_ao4 i_57679(.A(n_62123), .B(n_2071), .C(n_2070), .D(n_8561), .Z(n_1277
		));
	notech_ao4 i_57118(.A(n_62123), .B(n_8379), .C(n_8221), .D(n_8539), .Z(n_1280
		));
	notech_nand2 i_480(.A(cacheQ[127]), .B(n_1377), .Z(n_1281));
	notech_nand3 i_479(.A(n_60778), .B(axi_W[31]), .C(n_60760), .Z(n_1282)
		);
	notech_nand3 i_57115(.A(n_1282), .B(n_1579), .C(n_1281), .Z(n_1283));
	notech_nand2 i_484(.A(n_1377), .B(cacheQ[126]), .Z(n_1284));
	notech_nand3 i_483(.A(n_60778), .B(axi_W[30]), .C(n_60760), .Z(n_1285)
		);
	notech_nand3 i_57112(.A(n_1285), .B(n_1583), .C(n_1284), .Z(n_1286));
	notech_nand2 i_488(.A(n_1377), .B(cacheQ[125]), .Z(n_1287));
	notech_nand3 i_487(.A(n_60778), .B(axi_W[29]), .C(n_60756), .Z(n_1288)
		);
	notech_nand3 i_57109(.A(n_1288), .B(n_1587), .C(n_1287), .Z(n_1289));
	notech_nand2 i_492(.A(n_1377), .B(cacheQ[124]), .Z(n_1290));
	notech_nand3 i_491(.A(n_60778), .B(axi_W[28]), .C(n_60760), .Z(n_1291)
		);
	notech_nand3 i_57106(.A(n_1291), .B(n_1591), .C(n_1290), .Z(n_1292));
	notech_nand2 i_496(.A(n_1377), .B(cacheQ[123]), .Z(n_1293));
	notech_nand3 i_495(.A(n_60778), .B(axi_W[27]), .C(n_60760), .Z(n_1294)
		);
	notech_nand3 i_57103(.A(n_1294), .B(n_1595), .C(n_1293), .Z(n_1295));
	notech_nand2 i_500(.A(n_1377), .B(cacheQ[122]), .Z(n_1296));
	notech_nand3 i_499(.A(n_60779), .B(axi_W[26]), .C(n_60760), .Z(n_1297)
		);
	notech_nand3 i_57100(.A(n_1297), .B(n_1599), .C(n_1296), .Z(n_1298));
	notech_nand2 i_504(.A(n_1377), .B(cacheQ[121]), .Z(n_1299));
	notech_nand3 i_503(.A(n_60779), .B(axi_W[25]), .C(n_60760), .Z(n_1300)
		);
	notech_nand3 i_57097(.A(n_1300), .B(n_1603), .C(n_1299), .Z(n_1301));
	notech_nand2 i_508(.A(n_1377), .B(cacheQ[120]), .Z(n_1302));
	notech_nand3 i_507(.A(n_60778), .B(axi_W[24]), .C(n_60760), .Z(n_1303)
		);
	notech_nand3 i_57094(.A(n_1303), .B(n_1607), .C(n_1302), .Z(n_1304));
	notech_nand2 i_512(.A(n_1377), .B(cacheQ[119]), .Z(n_1305));
	notech_nand3 i_511(.A(n_60778), .B(axi_W[23]), .C(n_60760), .Z(n_1306)
		);
	notech_nand3 i_57091(.A(n_1306), .B(n_1611), .C(n_1305), .Z(n_1307));
	notech_nand2 i_516(.A(n_1377), .B(cacheQ[118]), .Z(n_1308));
	notech_nand3 i_515(.A(n_60778), .B(axi_W[22]), .C(n_60756), .Z(n_1309)
		);
	notech_nand3 i_57088(.A(n_1309), .B(n_1615), .C(n_1308), .Z(n_1310));
	notech_nand2 i_520(.A(n_1377), .B(cacheQ[117]), .Z(n_1311));
	notech_nand3 i_519(.A(n_60778), .B(axi_W[21]), .C(n_60756), .Z(n_1312)
		);
	notech_nand3 i_57085(.A(n_1312), .B(n_1619), .C(n_1311), .Z(n_1313));
	notech_nand2 i_524(.A(n_1377), .B(cacheQ[116]), .Z(n_1314));
	notech_nand3 i_523(.A(n_60778), .B(axi_W[20]), .C(n_60756), .Z(n_1315)
		);
	notech_nand3 i_57082(.A(n_1315), .B(n_1623), .C(n_1314), .Z(n_1316));
	notech_nand2 i_528(.A(n_1377), .B(cacheQ[115]), .Z(n_1317));
	notech_nand3 i_527(.A(n_60778), .B(axi_W[19]), .C(n_60756), .Z(n_1318)
		);
	notech_nand3 i_57079(.A(n_1318), .B(n_1627), .C(n_1317), .Z(n_1319));
	notech_nand2 i_532(.A(n_1377), .B(cacheQ[114]), .Z(n_1320));
	notech_nand3 i_531(.A(n_60778), .B(axi_W[18]), .C(n_60756), .Z(n_1321)
		);
	notech_nand3 i_57076(.A(n_1321), .B(n_1631), .C(n_1320), .Z(n_1322));
	notech_nand2 i_536(.A(n_1377), .B(cacheQ[113]), .Z(n_1323));
	notech_nand3 i_535(.A(n_60778), .B(axi_W[17]), .C(n_60756), .Z(n_1324)
		);
	notech_nand3 i_57073(.A(n_1324), .B(n_1635), .C(n_1323), .Z(n_1325));
	notech_nand2 i_540(.A(n_1377), .B(cacheQ[112]), .Z(n_1326));
	notech_nand3 i_539(.A(n_60778), .B(axi_W[16]), .C(n_60756), .Z(n_1327)
		);
	notech_nand3 i_57070(.A(n_1327), .B(n_1639), .C(n_1326), .Z(n_1328));
	notech_nand2 i_544(.A(n_60704), .B(cacheQ[111]), .Z(n_1329));
	notech_nand3 i_543(.A(n_60778), .B(axi_W[15]), .C(n_60756), .Z(n_1330)
		);
	notech_nand3 i_57067(.A(n_1330), .B(n_1643), .C(n_1329), .Z(n_1331));
	notech_nand2 i_548(.A(n_60704), .B(cacheQ[110]), .Z(n_1332));
	notech_nand3 i_547(.A(n_60778), .B(axi_W[14]), .C(n_60756), .Z(n_1333)
		);
	notech_nand3 i_57064(.A(n_1333), .B(n_1647), .C(n_1332), .Z(n_1334));
	notech_nand2 i_552(.A(n_60704), .B(cacheQ[109]), .Z(n_1335));
	notech_nand3 i_551(.A(n_60779), .B(axi_W[13]), .C(n_60756), .Z(n_1336)
		);
	notech_nand3 i_57061(.A(n_1336), .B(n_1651), .C(n_1335), .Z(n_1337));
	notech_nand2 i_556(.A(n_60704), .B(cacheQ[108]), .Z(n_1338));
	notech_nand3 i_555(.A(n_60779), .B(axi_W[12]), .C(n_60760), .Z(n_1339)
		);
	notech_nand3 i_57058(.A(n_1339), .B(n_1655), .C(n_1338), .Z(n_1340));
	notech_nand2 i_560(.A(n_60704), .B(cacheQ[107]), .Z(n_1341));
	notech_nand3 i_559(.A(n_60779), .B(axi_W[11]), .C(n_60762), .Z(n_1342)
		);
	notech_nand3 i_57055(.A(n_1342), .B(n_1659), .C(n_1341), .Z(n_1343));
	notech_nand2 i_564(.A(n_60704), .B(cacheQ[106]), .Z(n_1344));
	notech_nand3 i_563(.A(n_60779), .B(axi_W[10]), .C(n_60762), .Z(n_1345)
		);
	notech_nand3 i_57052(.A(n_1345), .B(n_1663), .C(n_1344), .Z(n_1346));
	notech_nand2 i_568(.A(n_60704), .B(cacheQ[105]), .Z(n_1347));
	notech_nand3 i_567(.A(n_60779), .B(axi_W[9]), .C(n_60762), .Z(n_1348));
	notech_nand3 i_57049(.A(n_1348), .B(n_1667), .C(n_1347), .Z(n_1349));
	notech_nand2 i_572(.A(n_60704), .B(cacheQ[104]), .Z(n_1350));
	notech_nand3 i_571(.A(n_60779), .B(axi_W[8]), .C(n_60762), .Z(n_1351));
	notech_nand3 i_57046(.A(n_1351), .B(n_1671), .C(n_1350), .Z(n_1352));
	notech_nand2 i_576(.A(n_60704), .B(cacheQ[103]), .Z(n_1353));
	notech_nand3 i_575(.A(n_60779), .B(axi_W[7]), .C(n_60762), .Z(n_1354));
	notech_nand3 i_57043(.A(n_1354), .B(n_1675), .C(n_1353), .Z(n_1355));
	notech_nand2 i_580(.A(n_60704), .B(cacheQ[102]), .Z(n_1356));
	notech_nand3 i_579(.A(n_60779), .B(axi_W[6]), .C(n_60762), .Z(n_1357));
	notech_nand3 i_57040(.A(n_1357), .B(n_1679), .C(n_1356), .Z(n_1358));
	notech_nand2 i_584(.A(n_60704), .B(cacheQ[101]), .Z(n_1359));
	notech_nand3 i_583(.A(n_60779), .B(axi_W[5]), .C(n_60762), .Z(n_1360));
	notech_nand3 i_57037(.A(n_1360), .B(n_1683), .C(n_1359), .Z(n_1361));
	notech_nand2 i_588(.A(n_60704), .B(cacheQ[100]), .Z(n_1362));
	notech_nand3 i_587(.A(n_60779), .B(axi_W[4]), .C(n_60762), .Z(n_1363));
	notech_nand3 i_57034(.A(n_1363), .B(n_1687), .C(n_1362), .Z(n_1364));
	notech_nand2 i_592(.A(n_60704), .B(cacheQ[99]), .Z(n_1365));
	notech_nand3 i_591(.A(n_60779), .B(axi_W[3]), .C(n_60762), .Z(n_1366));
	notech_nand3 i_57031(.A(n_1366), .B(n_1691), .C(n_1365), .Z(n_1367));
	notech_nand2 i_596(.A(n_60704), .B(cacheQ[98]), .Z(n_1368));
	notech_nand3 i_595(.A(n_60779), .B(axi_W[2]), .C(n_60762), .Z(n_1369));
	notech_nand3 i_57028(.A(n_1369), .B(n_1695), .C(n_1368), .Z(n_1370));
	notech_nand2 i_600(.A(n_60704), .B(cacheQ[97]), .Z(n_1371));
	notech_nand3 i_599(.A(n_60779), .B(axi_W[1]), .C(n_60760), .Z(n_1372));
	notech_nand3 i_57025(.A(n_1372), .B(n_1699), .C(n_1371), .Z(n_1373));
	notech_ao4 i_57678(.A(n_210856366), .B(n_2025), .C(n_2070), .D(n_8561), 
		.Z(n_1375));
	notech_nand2 i_606(.A(n_60704), .B(cacheQ[96]), .Z(n_1376));
	notech_nand2 i_19(.A(n_60743), .B(n_2073), .Z(n_1377));
	notech_nand3 i_605(.A(n_60779), .B(axi_W[0]), .C(n_60760), .Z(n_1378));
	notech_nand3 i_57022(.A(n_1378), .B(n_1706), .C(n_1376), .Z(n_1379));
	notech_nand2 i_610(.A(cacheQ[95]), .B(n_1476), .Z(n_1380));
	notech_nand3 i_609(.A(n_60779), .B(axi_W[31]), .C(n_60722), .Z(n_1381)
		);
	notech_nand3 i_57019(.A(n_1579), .B(n_1381), .C(n_1380), .Z(n_1382));
	notech_nand2 i_614(.A(n_1476), .B(cacheQ[94]), .Z(n_1383));
	notech_nand3 i_613(.A(n_60779), .B(axi_W[30]), .C(n_60725), .Z(n_1384)
		);
	notech_nand3 i_57016(.A(n_1583), .B(n_1384), .C(n_1383), .Z(n_1385));
	notech_nand2 i_618(.A(n_1476), .B(cacheQ[93]), .Z(n_1386));
	notech_nand3 i_617(.A(n_60779), .B(axi_W[29]), .C(n_60725), .Z(n_1387)
		);
	notech_nand3 i_57013(.A(n_1587), .B(n_1387), .C(n_1386), .Z(n_1388));
	notech_nand2 i_622(.A(n_1476), .B(cacheQ[92]), .Z(n_1389));
	notech_nand3 i_621(.A(n_60779), .B(axi_W[28]), .C(n_60722), .Z(n_1390)
		);
	notech_nand3 i_57010(.A(n_1591), .B(n_1390), .C(n_1389), .Z(n_1391));
	notech_nand2 i_626(.A(n_1476), .B(cacheQ[91]), .Z(n_1392));
	notech_nand3 i_625(.A(n_60778), .B(axi_W[27]), .C(n_60722), .Z(n_1393)
		);
	notech_nand3 i_57007(.A(n_1595), .B(n_1393), .C(n_1392), .Z(n_1394));
	notech_nand2 i_630(.A(n_1476), .B(cacheQ[90]), .Z(n_1395));
	notech_nand3 i_629(.A(n_60766), .B(axi_W[26]), .C(n_60722), .Z(n_1396)
		);
	notech_nand3 i_57004(.A(n_1599), .B(n_1396), .C(n_1395), .Z(n_1397));
	notech_nand2 i_634(.A(n_1476), .B(cacheQ[89]), .Z(n_1398));
	notech_nand3 i_633(.A(n_60766), .B(axi_W[25]), .C(n_60725), .Z(n_1399)
		);
	notech_nand3 i_57001(.A(n_1603), .B(n_1399), .C(n_1398), .Z(n_1400));
	notech_nand2 i_638(.A(n_1476), .B(cacheQ[88]), .Z(n_1401));
	notech_nand3 i_637(.A(n_60766), .B(axi_W[24]), .C(n_60725), .Z(n_1402)
		);
	notech_nand3 i_56998(.A(n_1607), .B(n_1402), .C(n_1401), .Z(n_1403));
	notech_nand2 i_642(.A(n_1476), .B(cacheQ[87]), .Z(n_1404));
	notech_nand3 i_641(.A(n_60766), .B(axi_W[23]), .C(n_60725), .Z(n_1405)
		);
	notech_nand3 i_56995(.A(n_1611), .B(n_1405), .C(n_1404), .Z(n_1406));
	notech_nand2 i_646(.A(n_1476), .B(cacheQ[86]), .Z(n_1407));
	notech_nand3 i_645(.A(n_60772), .B(axi_W[22]), .C(n_60725), .Z(n_1408)
		);
	notech_nand3 i_56992(.A(n_1615), .B(n_1408), .C(n_1407), .Z(n_1409));
	notech_nand2 i_650(.A(n_1476), .B(cacheQ[85]), .Z(n_1410));
	notech_nand3 i_649(.A(n_60772), .B(axi_W[21]), .C(n_60725), .Z(n_1411)
		);
	notech_nand3 i_56989(.A(n_1619), .B(n_1411), .C(n_1410), .Z(n_1412));
	notech_nand2 i_654(.A(n_1476), .B(cacheQ[84]), .Z(n_1413));
	notech_nand3 i_653(.A(n_60772), .B(axi_W[20]), .C(n_60725), .Z(n_1414)
		);
	notech_nand3 i_56986(.A(n_1623), .B(n_1414), .C(n_1413), .Z(n_1415));
	notech_nand2 i_658(.A(n_1476), .B(cacheQ[83]), .Z(n_1416));
	notech_nand3 i_657(.A(n_60772), .B(axi_W[19]), .C(n_60725), .Z(n_1417)
		);
	notech_nand3 i_56983(.A(n_1627), .B(n_1417), .C(n_1416), .Z(n_1418));
	notech_nand2 i_662(.A(n_1476), .B(cacheQ[82]), .Z(n_1419));
	notech_nand3 i_661(.A(n_60772), .B(axi_W[18]), .C(n_60722), .Z(n_1420)
		);
	notech_nand3 i_56980(.A(n_1631), .B(n_1420), .C(n_1419), .Z(n_1421));
	notech_nand2 i_666(.A(n_1476), .B(cacheQ[81]), .Z(n_1422));
	notech_nand3 i_665(.A(n_60766), .B(axi_W[17]), .C(n_60722), .Z(n_1423)
		);
	notech_nand3 i_56977(.A(n_1635), .B(n_1423), .C(n_1422), .Z(n_1424));
	notech_nand2 i_670(.A(n_1476), .B(cacheQ[80]), .Z(n_1425));
	notech_nand3 i_669(.A(n_60766), .B(axi_W[16]), .C(n_60722), .Z(n_1426)
		);
	notech_nand3 i_56974(.A(n_1639), .B(n_1426), .C(n_1425), .Z(n_1427));
	notech_nand2 i_674(.A(n_60682), .B(cacheQ[79]), .Z(n_1428));
	notech_nand3 i_673(.A(n_60766), .B(axi_W[15]), .C(n_60722), .Z(n_1429)
		);
	notech_nand3 i_56971(.A(n_1643), .B(n_1429), .C(n_1428), .Z(n_1430));
	notech_nand2 i_678(.A(n_60682), .B(cacheQ[78]), .Z(n_1431));
	notech_nand3 i_677(.A(n_60766), .B(axi_W[14]), .C(n_60722), .Z(n_1432)
		);
	notech_nand3 i_56968(.A(n_1647), .B(n_1432), .C(n_1431), .Z(n_1433));
	notech_nand2 i_682(.A(n_60682), .B(cacheQ[77]), .Z(n_1434));
	notech_nand3 i_681(.A(n_60766), .B(axi_W[13]), .C(n_60722), .Z(n_1435)
		);
	notech_nand3 i_56965(.A(n_1651), .B(n_1435), .C(n_1434), .Z(n_1436));
	notech_nand2 i_686(.A(n_60682), .B(cacheQ[76]), .Z(n_1437));
	notech_nand3 i_685(.A(n_60766), .B(axi_W[12]), .C(n_60722), .Z(n_1438)
		);
	notech_nand3 i_56962(.A(n_1655), .B(n_1438), .C(n_1437), .Z(n_1439));
	notech_nand2 i_690(.A(n_60682), .B(cacheQ[75]), .Z(n_1440));
	notech_nand3 i_689(.A(n_60766), .B(axi_W[11]), .C(n_60722), .Z(n_1441)
		);
	notech_nand3 i_56959(.A(n_1659), .B(n_1441), .C(n_1440), .Z(n_1442));
	notech_nand2 i_694(.A(n_60682), .B(cacheQ[74]), .Z(n_1443));
	notech_nand3 i_693(.A(n_60766), .B(axi_W[10]), .C(n_60722), .Z(n_1444)
		);
	notech_nand3 i_56956(.A(n_1663), .B(n_1444), .C(n_1443), .Z(n_1445));
	notech_nand2 i_698(.A(n_60682), .B(cacheQ[73]), .Z(n_1446));
	notech_nand3 i_697(.A(n_60766), .B(axi_W[9]), .C(n_60722), .Z(n_1447));
	notech_nand3 i_56953(.A(n_1667), .B(n_1447), .C(n_1446), .Z(n_1448));
	notech_nand2 i_702(.A(n_60682), .B(cacheQ[72]), .Z(n_1449));
	notech_nand3 i_701(.A(n_60772), .B(axi_W[8]), .C(n_60722), .Z(n_1450));
	notech_nand3 i_56950(.A(n_1671), .B(n_1450), .C(n_1449), .Z(n_1451));
	notech_nand2 i_706(.A(n_60682), .B(cacheQ[71]), .Z(n_1452));
	notech_nand3 i_705(.A(n_60772), .B(axi_W[7]), .C(n_60722), .Z(n_1453));
	notech_nand3 i_56947(.A(n_1675), .B(n_1453), .C(n_1452), .Z(n_1454));
	notech_nand2 i_710(.A(n_60682), .B(cacheQ[70]), .Z(n_1455));
	notech_nand3 i_709(.A(n_60772), .B(axi_W[6]), .C(n_60722), .Z(n_1456));
	notech_nand3 i_56944(.A(n_1679), .B(n_1456), .C(n_1455), .Z(n_1457));
	notech_nand2 i_714(.A(n_60682), .B(cacheQ[69]), .Z(n_1458));
	notech_nand3 i_713(.A(n_60772), .B(axi_W[5]), .C(n_60725), .Z(n_1459));
	notech_nand3 i_56941(.A(n_1683), .B(n_1459), .C(n_1458), .Z(n_1460));
	notech_nand2 i_718(.A(n_60682), .B(cacheQ[68]), .Z(n_1461));
	notech_nand3 i_717(.A(n_60772), .B(axi_W[4]), .C(n_60727), .Z(n_1462));
	notech_nand3 i_56938(.A(n_1687), .B(n_1462), .C(n_1461), .Z(n_1463));
	notech_nand2 i_722(.A(n_60682), .B(cacheQ[67]), .Z(n_1464));
	notech_nand3 i_721(.A(n_60778), .B(axi_W[3]), .C(n_60727), .Z(n_1465));
	notech_nand3 i_56935(.A(n_1691), .B(n_1465), .C(n_1464), .Z(n_1466));
	notech_nand2 i_726(.A(n_60682), .B(cacheQ[66]), .Z(n_1467));
	notech_nand3 i_725(.A(n_60778), .B(axi_W[2]), .C(n_60727), .Z(n_1468));
	notech_nand3 i_56932(.A(n_1695), .B(n_1468), .C(n_1467), .Z(n_1469));
	notech_nand2 i_730(.A(n_60682), .B(cacheQ[65]), .Z(n_1470));
	notech_nand3 i_729(.A(n_60772), .B(axi_W[1]), .C(n_60727), .Z(n_1471));
	notech_nand3 i_56929(.A(n_1699), .B(n_1471), .C(n_1470), .Z(n_1472));
	notech_ao4 i_57677(.A(n_210856366), .B(n_8223), .C(n_2070), .D(n_8561), 
		.Z(n_1474));
	notech_nand2 i_736(.A(n_60682), .B(cacheQ[64]), .Z(n_1475));
	notech_nand2 i_18(.A(n_60743), .B(n_2075), .Z(n_1476));
	notech_nand3 i_735(.A(n_60778), .B(axi_W[0]), .C(n_60727), .Z(n_1477));
	notech_nand3 i_56926(.A(n_1706), .B(n_1477), .C(n_1475), .Z(n_1478));
	notech_nand2 i_740(.A(cacheQ[63]), .B(n_1575), .Z(n_1479));
	notech_nao3 i_739(.A(axi_W[31]), .B(n_60760), .C(n_60743), .Z(n_1480));
	notech_nand3 i_56923(.A(n_1579), .B(n_1480), .C(n_1479), .Z(n_1481));
	notech_nand2 i_744(.A(n_1575), .B(cacheQ[62]), .Z(n_1482));
	notech_nao3 i_743(.A(axi_W[30]), .B(n_60760), .C(n_60743), .Z(n_1483));
	notech_nand3 i_56920(.A(n_1583), .B(n_1483), .C(n_1482), .Z(n_1484));
	notech_nand2 i_748(.A(n_1575), .B(cacheQ[61]), .Z(n_1485));
	notech_nao3 i_747(.A(axi_W[29]), .B(n_60760), .C(n_60743), .Z(n_1486));
	notech_nand3 i_56917(.A(n_1587), .B(n_1486), .C(n_1485), .Z(n_1487));
	notech_nand2 i_752(.A(n_1575), .B(cacheQ[60]), .Z(n_1488));
	notech_nao3 i_751(.A(axi_W[28]), .B(n_60762), .C(n_60743), .Z(n_1489));
	notech_nand3 i_56914(.A(n_1591), .B(n_1489), .C(n_1488), .Z(n_1490));
	notech_nand2 i_756(.A(n_1575), .B(cacheQ[59]), .Z(n_1491));
	notech_nao3 i_755(.A(axi_W[27]), .B(n_60762), .C(n_60744), .Z(n_1492));
	notech_nand3 i_56911(.A(n_1595), .B(n_1492), .C(n_1491), .Z(n_1493));
	notech_nand2 i_760(.A(n_1575), .B(cacheQ[58]), .Z(n_1494));
	notech_nao3 i_759(.A(axi_W[26]), .B(n_60762), .C(n_60743), .Z(n_1495));
	notech_nand3 i_56908(.A(n_1599), .B(n_1495), .C(n_1494), .Z(n_1496));
	notech_nand2 i_764(.A(n_1575), .B(cacheQ[57]), .Z(n_1497));
	notech_nao3 i_763(.A(axi_W[25]), .B(n_60762), .C(n_60743), .Z(n_1498));
	notech_nand3 i_56905(.A(n_1603), .B(n_1498), .C(n_1497), .Z(n_1499));
	notech_nand2 i_768(.A(n_1575), .B(cacheQ[56]), .Z(n_1500));
	notech_nao3 i_767(.A(axi_W[24]), .B(n_60762), .C(n_60743), .Z(n_1501));
	notech_nand3 i_56902(.A(n_1607), .B(n_1501), .C(n_1500), .Z(n_1502));
	notech_nand2 i_772(.A(n_1575), .B(cacheQ[55]), .Z(n_1503));
	notech_nao3 i_771(.A(axi_W[23]), .B(n_60762), .C(n_60743), .Z(n_1504));
	notech_nand3 i_56899(.A(n_1611), .B(n_1504), .C(n_1503), .Z(n_1505));
	notech_nand2 i_776(.A(n_1575), .B(cacheQ[54]), .Z(n_1506));
	notech_nao3 i_775(.A(axi_W[22]), .B(n_60755), .C(n_60743), .Z(n_1507));
	notech_nand3 i_56896(.A(n_1615), .B(n_1507), .C(n_1506), .Z(n_1508));
	notech_nand2 i_780(.A(n_1575), .B(cacheQ[53]), .Z(n_1509));
	notech_nao3 i_779(.A(axi_W[21]), .B(n_60755), .C(n_60743), .Z(n_1510));
	notech_nand3 i_56893(.A(n_1619), .B(n_1510), .C(n_1509), .Z(n_1511));
	notech_nand2 i_784(.A(n_1575), .B(cacheQ[52]), .Z(n_1512));
	notech_nao3 i_783(.A(axi_W[20]), .B(n_60762), .C(n_60743), .Z(n_1513));
	notech_nand3 i_56890(.A(n_1623), .B(n_1513), .C(n_1512), .Z(n_1514));
	notech_nand2 i_788(.A(n_1575), .B(cacheQ[51]), .Z(n_1515));
	notech_nao3 i_787(.A(axi_W[19]), .B(n_60762), .C(n_60743), .Z(n_1516));
	notech_nand3 i_56887(.A(n_1627), .B(n_1516), .C(n_1515), .Z(n_1517));
	notech_nand2 i_792(.A(n_1575), .B(cacheQ[50]), .Z(n_1518));
	notech_nao3 i_791(.A(axi_W[18]), .B(n_60760), .C(n_60743), .Z(n_1519));
	notech_nand3 i_56884(.A(n_1631), .B(n_1519), .C(n_1518), .Z(n_1520));
	notech_nand2 i_796(.A(n_1575), .B(cacheQ[49]), .Z(n_1521));
	notech_nao3 i_795(.A(axi_W[17]), .B(n_60762), .C(n_60743), .Z(n_1522));
	notech_nand3 i_56881(.A(n_1635), .B(n_1522), .C(n_1521), .Z(n_1523));
	notech_nand2 i_800(.A(n_1575), .B(cacheQ[48]), .Z(n_1524));
	notech_nao3 i_799(.A(axi_W[16]), .B(n_60762), .C(n_60743), .Z(n_1525));
	notech_nand3 i_56878(.A(n_1639), .B(n_1525), .C(n_1524), .Z(n_1526));
	notech_nand2 i_804(.A(n_60660), .B(cacheQ[47]), .Z(n_1527));
	notech_nao3 i_803(.A(axi_W[15]), .B(n_60755), .C(n_60744), .Z(n_1528));
	notech_nand3 i_56875(.A(n_1643), .B(n_1528), .C(n_1527), .Z(n_1529));
	notech_nand2 i_808(.A(n_60660), .B(cacheQ[46]), .Z(n_1530));
	notech_nao3 i_807(.A(axi_W[14]), .B(n_60750), .C(n_60744), .Z(n_1531));
	notech_nand3 i_56872(.A(n_1647), .B(n_1531), .C(n_1530), .Z(n_1532));
	notech_nand2 i_812(.A(n_60660), .B(cacheQ[45]), .Z(n_1533));
	notech_nao3 i_811(.A(axi_W[13]), .B(n_60750), .C(n_60744), .Z(n_1534));
	notech_nand3 i_56869(.A(n_1651), .B(n_1534), .C(n_1533), .Z(n_1535));
	notech_nand2 i_816(.A(n_60660), .B(cacheQ[44]), .Z(n_1536));
	notech_nao3 i_815(.A(axi_W[12]), .B(n_60750), .C(n_60744), .Z(n_1537));
	notech_nand3 i_56866(.A(n_1655), .B(n_1537), .C(n_1536), .Z(n_1538));
	notech_nand2 i_820(.A(n_60660), .B(cacheQ[43]), .Z(n_1539));
	notech_nao3 i_819(.A(axi_W[11]), .B(n_60750), .C(n_60744), .Z(n_1540));
	notech_nand3 i_56863(.A(n_1659), .B(n_1540), .C(n_1539), .Z(n_1541));
	notech_nand2 i_824(.A(n_60660), .B(cacheQ[42]), .Z(n_1542));
	notech_nao3 i_823(.A(axi_W[10]), .B(n_60750), .C(n_60744), .Z(n_1543));
	notech_nand3 i_56860(.A(n_1663), .B(n_1543), .C(n_1542), .Z(n_1544));
	notech_nand2 i_828(.A(n_60660), .B(cacheQ[41]), .Z(n_1545));
	notech_nao3 i_827(.A(axi_W[9]), .B(n_60755), .C(n_60744), .Z(n_1546));
	notech_nand3 i_56857(.A(n_1667), .B(n_1546), .C(n_1545), .Z(n_1547));
	notech_nand2 i_832(.A(n_60660), .B(cacheQ[40]), .Z(n_1548));
	notech_nao3 i_831(.A(axi_W[8]), .B(n_60755), .C(n_60744), .Z(n_1549));
	notech_nand3 i_56854(.A(n_1671), .B(n_1549), .C(n_1548), .Z(n_1550));
	notech_nand2 i_836(.A(n_60660), .B(cacheQ[39]), .Z(n_1551));
	notech_nao3 i_835(.A(axi_W[7]), .B(n_60750), .C(n_60744), .Z(n_1552));
	notech_nand3 i_56851(.A(n_1675), .B(n_1552), .C(n_1551), .Z(n_1553));
	notech_nand2 i_840(.A(n_60660), .B(cacheQ[38]), .Z(n_1554));
	notech_nao3 i_839(.A(axi_W[6]), .B(n_60755), .C(n_60744), .Z(n_1555));
	notech_nand3 i_56848(.A(n_1679), .B(n_1555), .C(n_1554), .Z(n_1556));
	notech_nand2 i_844(.A(n_60660), .B(cacheQ[37]), .Z(n_1557));
	notech_nao3 i_843(.A(axi_W[5]), .B(n_60760), .C(n_60744), .Z(n_1558));
	notech_nand3 i_56845(.A(n_1683), .B(n_1558), .C(n_1557), .Z(n_1559));
	notech_nand2 i_848(.A(n_60660), .B(cacheQ[36]), .Z(n_1560));
	notech_nao3 i_847(.A(axi_W[4]), .B(n_60756), .C(n_60744), .Z(n_1561));
	notech_nand3 i_56842(.A(n_1687), .B(n_1561), .C(n_1560), .Z(n_1562));
	notech_nand2 i_852(.A(n_60660), .B(cacheQ[35]), .Z(n_1563));
	notech_nao3 i_851(.A(axi_W[3]), .B(n_60756), .C(n_60744), .Z(n_1564));
	notech_nand3 i_56839(.A(n_1691), .B(n_1564), .C(n_1563), .Z(n_1565));
	notech_nand2 i_856(.A(n_60660), .B(cacheQ[34]), .Z(n_1566));
	notech_nao3 i_855(.A(axi_W[2]), .B(n_60756), .C(n_60744), .Z(n_1567));
	notech_nand3 i_56836(.A(n_1695), .B(n_1567), .C(n_1566), .Z(n_1568));
	notech_nand2 i_860(.A(n_60660), .B(cacheQ[33]), .Z(n_1569));
	notech_nao3 i_859(.A(axi_W[1]), .B(n_60756), .C(n_60744), .Z(n_1570));
	notech_nand3 i_56833(.A(n_1699), .B(n_1570), .C(n_1569), .Z(n_1571));
	notech_ao4 i_57676(.A(n_210856366), .B(n_8222), .C(n_2070), .D(n_8561), 
		.Z(n_1573));
	notech_nand2 i_866(.A(n_60660), .B(cacheQ[32]), .Z(n_1574));
	notech_or2 i_17(.A(n_60772), .B(n_214256400), .Z(n_1575));
	notech_nao3 i_865(.A(axi_W[0]), .B(n_60756), .C(n_60744), .Z(n_1576));
	notech_nand3 i_56830(.A(n_1706), .B(n_1576), .C(n_1574), .Z(n_1577));
	notech_nand2 i_870(.A(cacheQ[31]), .B(n_1705), .Z(n_1578));
	notech_nand2 i_104(.A(axi_R[31]), .B(n_2023), .Z(n_1579));
	notech_nao3 i_869(.A(axi_W[31]), .B(n_60727), .C(n_60744), .Z(n_1580));
	notech_nand3 i_56827(.A(n_1579), .B(n_1580), .C(n_1578), .Z(n_1581));
	notech_nand2 i_874(.A(n_1705), .B(cacheQ[30]), .Z(n_1582));
	notech_nand2 i_102(.A(axi_R[30]), .B(n_2023), .Z(n_1583));
	notech_nao3 i_873(.A(axi_W[30]), .B(n_60727), .C(n_60744), .Z(n_1584));
	notech_nand3 i_56824(.A(n_1583), .B(n_1584), .C(n_1582), .Z(n_1585));
	notech_nand2 i_878(.A(n_1705), .B(cacheQ[29]), .Z(n_1586));
	notech_nand2 i_101(.A(axi_R[29]), .B(n_2023), .Z(n_1587));
	notech_nao3 i_877(.A(axi_W[29]), .B(n_60727), .C(n_60744), .Z(n_1588));
	notech_nand3 i_56821(.A(n_1587), .B(n_1588), .C(n_1586), .Z(n_1589));
	notech_nand2 i_882(.A(n_1705), .B(cacheQ[28]), .Z(n_1590));
	notech_nand2 i_106(.A(axi_R[28]), .B(n_2023), .Z(n_1591));
	notech_nao3 i_881(.A(axi_W[28]), .B(n_60727), .C(n_60731), .Z(n_1592));
	notech_nand3 i_56818(.A(n_1591), .B(n_1592), .C(n_1590), .Z(n_1593));
	notech_nand2 i_886(.A(n_1705), .B(cacheQ[27]), .Z(n_1594));
	notech_nand2 i_99(.A(axi_R[27]), .B(n_2023), .Z(n_1595));
	notech_nao3 i_885(.A(axi_W[27]), .B(n_60727), .C(n_60731), .Z(n_1596));
	notech_nand3 i_56815(.A(n_1595), .B(n_1596), .C(n_1594), .Z(n_1597));
	notech_nand2 i_890(.A(n_1705), .B(cacheQ[26]), .Z(n_1598));
	notech_nand2 i_97(.A(axi_R[26]), .B(n_2023), .Z(n_1599));
	notech_nao3 i_889(.A(axi_W[26]), .B(n_60727), .C(n_60731), .Z(n_1600));
	notech_nand3 i_56812(.A(n_1599), .B(n_1600), .C(n_1598), .Z(n_1601));
	notech_nand2 i_901(.A(n_1705), .B(cacheQ[25]), .Z(n_1602));
	notech_nand2 i_76(.A(axi_R[25]), .B(n_2023), .Z(n_1603));
	notech_nao3 i_897(.A(axi_W[25]), .B(n_60727), .C(n_60731), .Z(n_1604));
	notech_nand3 i_56809(.A(n_1603), .B(n_1604), .C(n_1602), .Z(n_1605));
	notech_nand2 i_905(.A(n_1705), .B(cacheQ[24]), .Z(n_1606));
	notech_nand2 i_108(.A(axi_R[24]), .B(n_2023), .Z(n_1607));
	notech_nao3 i_904(.A(axi_W[24]), .B(n_60727), .C(n_60731), .Z(n_1608));
	notech_nand3 i_56806(.A(n_1607), .B(n_1608), .C(n_1606), .Z(n_1609));
	notech_nand2 i_909(.A(n_1705), .B(cacheQ[23]), .Z(n_1610));
	notech_nand2 i_96(.A(axi_R[23]), .B(n_2023), .Z(n_1611));
	notech_nao3 i_908(.A(axi_W[23]), .B(n_60725), .C(n_60737), .Z(n_1612));
	notech_nand3 i_56803(.A(n_1611), .B(n_1612), .C(n_1610), .Z(n_1613));
	notech_nand2 i_913(.A(n_1705), .B(cacheQ[22]), .Z(n_1614));
	notech_nand2 i_95(.A(axi_R[22]), .B(n_2023), .Z(n_1615));
	notech_nao3 i_912(.A(axi_W[22]), .B(n_60725), .C(n_60737), .Z(n_1616));
	notech_nand3 i_56800(.A(n_1615), .B(n_1616), .C(n_1614), .Z(n_1617));
	notech_nand2 i_917(.A(n_1705), .B(cacheQ[21]), .Z(n_1618));
	notech_nand2 i_94(.A(axi_R[21]), .B(n_2023), .Z(n_1619));
	notech_nao3 i_916(.A(axi_W[21]), .B(n_60725), .C(n_60737), .Z(n_1620));
	notech_nand3 i_56797(.A(n_1619), .B(n_1620), .C(n_1618), .Z(n_1621));
	notech_nand2 i_924(.A(n_1705), .B(cacheQ[20]), .Z(n_1622));
	notech_nand2 i_86(.A(axi_R[20]), .B(n_2023), .Z(n_1623));
	notech_nao3 i_923(.A(axi_W[20]), .B(n_60725), .C(n_60737), .Z(n_1624));
	notech_nand3 i_56794(.A(n_1623), .B(n_1624), .C(n_1622), .Z(n_1625));
	notech_nand2 i_928(.A(n_1705), .B(cacheQ[19]), .Z(n_1626));
	notech_nand2 i_88(.A(axi_R[19]), .B(n_2023), .Z(n_1627));
	notech_nao3 i_927(.A(axi_W[19]), .B(n_60725), .C(n_60731), .Z(n_1628));
	notech_nand3 i_56791(.A(n_1627), .B(n_1628), .C(n_1626), .Z(n_1629));
	notech_nand2 i_932(.A(n_1705), .B(cacheQ[18]), .Z(n_1630));
	notech_nand2 i_89(.A(axi_R[18]), .B(n_2023), .Z(n_1631));
	notech_nao3 i_931(.A(axi_W[18]), .B(n_60725), .C(n_60731), .Z(n_1632));
	notech_nand3 i_56788(.A(n_1631), .B(n_1632), .C(n_1630), .Z(n_1633));
	notech_nand2 i_936(.A(n_1705), .B(cacheQ[17]), .Z(n_1634));
	notech_nand2 i_90(.A(axi_R[17]), .B(n_2023), .Z(n_1635));
	notech_nao3 i_935(.A(axi_W[17]), .B(n_60725), .C(n_60731), .Z(n_1636));
	notech_nand3 i_56785(.A(n_1635), .B(n_1636), .C(n_1634), .Z(n_1637));
	notech_nand2 i_940(.A(n_1705), .B(cacheQ[16]), .Z(n_1638));
	notech_nand2 i_91(.A(axi_R[16]), .B(n_2023), .Z(n_1639));
	notech_nao3 i_939(.A(axi_W[16]), .B(n_60727), .C(n_60731), .Z(n_1640));
	notech_nand3 i_56782(.A(n_1639), .B(n_1640), .C(n_1638), .Z(n_1641));
	notech_nand2 i_944(.A(n_60638), .B(cacheQ[15]), .Z(n_1642));
	notech_nand2 i_92(.A(axi_R[15]), .B(n_2023), .Z(n_1643));
	notech_nao3 i_943(.A(axi_W[15]), .B(n_60727), .C(n_60731), .Z(n_1644));
	notech_nand3 i_56779(.A(n_1643), .B(n_1644), .C(n_1642), .Z(n_1645));
	notech_nand2 i_948(.A(n_60638), .B(cacheQ[14]), .Z(n_1646));
	notech_nand2 i_93(.A(axi_R[14]), .B(n_2023), .Z(n_1647));
	notech_nao3 i_947(.A(axi_W[14]), .B(n_60727), .C(n_60731), .Z(n_1648));
	notech_nand3 i_56776(.A(n_1647), .B(n_1648), .C(n_1646), .Z(n_1649));
	notech_nand2 i_952(.A(n_60638), .B(cacheQ[13]), .Z(n_1650));
	notech_nand2 i_87(.A(axi_R[13]), .B(n_62132), .Z(n_1651));
	notech_nao3 i_951(.A(axi_W[13]), .B(n_60725), .C(n_60731), .Z(n_1652));
	notech_nand3 i_56773(.A(n_1651), .B(n_1652), .C(n_1650), .Z(n_1653));
	notech_nand2 i_956(.A(n_60638), .B(cacheQ[12]), .Z(n_1654));
	notech_nand2 i_103(.A(axi_R[12]), .B(n_62132), .Z(n_1655));
	notech_nao3 i_955(.A(axi_W[12]), .B(n_60727), .C(n_60731), .Z(n_1656));
	notech_nand3 i_56770(.A(n_1655), .B(n_1656), .C(n_1654), .Z(n_1657));
	notech_nand2 i_960(.A(n_60638), .B(cacheQ[11]), .Z(n_1658));
	notech_nand2 i_85(.A(axi_R[11]), .B(n_62132), .Z(n_1659));
	notech_nao3 i_959(.A(axi_W[11]), .B(n_60727), .C(n_60731), .Z(n_1660));
	notech_nand3 i_56767(.A(n_1659), .B(n_1660), .C(n_1658), .Z(n_1661));
	notech_nand2 i_964(.A(n_60638), .B(cacheQ[10]), .Z(n_1662));
	notech_nand2 i_84(.A(axi_R[10]), .B(n_62132), .Z(n_1663));
	notech_nao3 i_963(.A(axi_W[10]), .B(n_60722), .C(n_60737), .Z(n_1664));
	notech_nand3 i_56764(.A(n_1663), .B(n_1664), .C(n_1662), .Z(n_1665));
	notech_nand2 i_968(.A(n_60638), .B(cacheQ[9]), .Z(n_1666));
	notech_nand2 i_83(.A(axi_R[9]), .B(n_62132), .Z(n_1667));
	notech_nao3 i_967(.A(axi_W[9]), .B(n_60715), .C(n_60737), .Z(n_1668));
	notech_nand3 i_56761(.A(n_1667), .B(n_1668), .C(n_1666), .Z(n_1669));
	notech_nand2 i_972(.A(n_60638), .B(cacheQ[8]), .Z(n_1670));
	notech_nand2 i_82(.A(axi_R[8]), .B(n_62132), .Z(n_1671));
	notech_nao3 i_971(.A(axi_W[8]), .B(n_60717), .C(n_60737), .Z(n_1672));
	notech_nand3 i_56758(.A(n_1671), .B(n_1672), .C(n_1670), .Z(n_1673));
	notech_nand2 i_976(.A(n_60638), .B(cacheQ[7]), .Z(n_1674));
	notech_nand2 i_81(.A(axi_R[7]), .B(n_62132), .Z(n_1675));
	notech_nao3 i_975(.A(axi_W[7]), .B(n_60717), .C(n_60737), .Z(n_1676));
	notech_nand3 i_56755(.A(n_1675), .B(n_1676), .C(n_1674), .Z(n_1677));
	notech_nand2 i_980(.A(n_60638), .B(cacheQ[6]), .Z(n_1678));
	notech_nand2 i_80(.A(axi_R[6]), .B(n_62132), .Z(n_1679));
	notech_nao3 i_979(.A(axi_W[6]), .B(n_60715), .C(n_60737), .Z(n_1680));
	notech_nand3 i_56752(.A(n_1679), .B(n_1680), .C(n_1678), .Z(n_1681));
	notech_nand2 i_984(.A(n_60638), .B(cacheQ[5]), .Z(n_1682));
	notech_nand2 i_79(.A(axi_R[5]), .B(n_62132), .Z(n_1683));
	notech_nao3 i_983(.A(axi_W[5]), .B(n_60715), .C(n_60737), .Z(n_1684));
	notech_nand3 i_56749(.A(n_1683), .B(n_1684), .C(n_1682), .Z(n_1685));
	notech_nand2 i_988(.A(n_60638), .B(cacheQ[4]), .Z(n_1686));
	notech_nand2 i_107(.A(axi_R[4]), .B(n_62132), .Z(n_1687));
	notech_nao3 i_987(.A(axi_W[4]), .B(n_60715), .C(n_60743), .Z(n_1688));
	notech_nand3 i_56746(.A(n_1687), .B(n_1688), .C(n_1686), .Z(n_1689));
	notech_nand2 i_992(.A(n_60638), .B(cacheQ[3]), .Z(n_1690));
	notech_nand2 i_100(.A(axi_R[3]), .B(n_62132), .Z(n_1691));
	notech_nao3 i_991(.A(axi_W[3]), .B(n_60717), .C(n_60743), .Z(n_1692));
	notech_nand3 i_56743(.A(n_1691), .B(n_1692), .C(n_1690), .Z(n_1693));
	notech_nand2 i_996(.A(n_60638), .B(cacheQ[2]), .Z(n_1694));
	notech_nand2 i_77(.A(axi_R[2]), .B(n_62132), .Z(n_1695));
	notech_nao3 i_995(.A(axi_W[2]), .B(n_60717), .C(n_60737), .Z(n_1696));
	notech_nand3 i_56740(.A(n_1695), .B(n_1696), .C(n_1694), .Z(n_1697));
	notech_nand2 i_1000(.A(n_60638), .B(cacheQ[1]), .Z(n_1698));
	notech_nand2 i_74(.A(axi_R[1]), .B(n_62132), .Z(n_1699));
	notech_nao3 i_999(.A(axi_W[1]), .B(n_60717), .C(n_60743), .Z(n_1700));
	notech_nand3 i_56737(.A(n_1699), .B(n_1700), .C(n_1698), .Z(n_1701));
	notech_ao4 i_57675(.A(n_210856366), .B(n_2036), .C(n_2070), .D(n_8561), 
		.Z(n_1703));
	notech_nand2 i_1006(.A(n_60638), .B(cacheQ[0]), .Z(n_1704));
	notech_or2 i_16(.A(n_60772), .B(n_214356401), .Z(n_1705));
	notech_nand2 i_98(.A(axi_R[0]), .B(n_62132), .Z(n_1706));
	notech_nao3 i_1005(.A(axi_W[0]), .B(n_60717), .C(n_60737), .Z(n_1707));
	notech_nand3 i_56734(.A(n_1706), .B(n_1707), .C(n_1704), .Z(n_1708));
	notech_ao4 i_56147(.A(n_8323), .B(n_8558), .C(n_2002), .D(n_2007), .Z(n_1710
		));
	notech_nand2 i_1011(.A(n_2033), .B(n_21466), .Z(n_1711));
	notech_nand3 i_1014(.A(n_60772), .B(axi_WSTRB[3]), .C(n_60756), .Z(n_1712
		));
	notech_nand3 i_57211(.A(n_62815), .B(n_220956467), .C(n_1712), .Z(n_1713
		));
	notech_nand3 i_1016(.A(n_60772), .B(axi_WSTRB[2]), .C(n_60756), .Z(n_1714
		));
	notech_nand3 i_57209(.A(n_62815), .B(n_220956467), .C(n_1714), .Z(n_1715
		));
	notech_nand3 i_1018(.A(n_60772), .B(axi_WSTRB[1]), .C(n_60756), .Z(n_1716
		));
	notech_nand3 i_57207(.A(n_62815), .B(n_220956467), .C(n_1716), .Z(n_1717
		));
	notech_and4 i_1020(.A(A4[1]), .B(n_60756), .C(axi_WSTRB[0]), .D(n_2069),
		 .Z(n_1718));
	notech_nao3 i_57205(.A(n_62815), .B(n_220956467), .C(n_1718), .Z(n_1719)
		);
	notech_nand3 i_1022(.A(n_60772), .B(axi_WSTRB[3]), .C(n_60717), .Z(n_1720
		));
	notech_nand3 i_57203(.A(n_62815), .B(n_220956467), .C(n_1720), .Z(n_1721
		));
	notech_nand3 i_1024(.A(n_60772), .B(axi_WSTRB[2]), .C(n_60717), .Z(n_1722
		));
	notech_nand3 i_57201(.A(n_62815), .B(n_220956467), .C(n_1722), .Z(n_1723
		));
	notech_nand3 i_1026(.A(n_60772), .B(axi_WSTRB[1]), .C(n_60717), .Z(n_1724
		));
	notech_nand3 i_57199(.A(n_62815), .B(n_220956467), .C(n_1724), .Z(n_1725
		));
	notech_nand3 i_1028(.A(axi_WSTRB[0]), .B(n_60715), .C(n_60772), .Z(n_1726
		));
	notech_nand3 i_57197(.A(n_62815), .B(n_220956467), .C(n_1726), .Z(n_1727
		));
	notech_nao3 i_1030(.A(axi_WSTRB[3]), .B(n_60755), .C(n_60737), .Z(n_1728
		));
	notech_nand3 i_57195(.A(n_62815), .B(n_220956467), .C(n_1728), .Z(n_1729
		));
	notech_nao3 i_1032(.A(axi_WSTRB[2]), .B(n_60760), .C(n_60737), .Z(n_1730
		));
	notech_nand3 i_57193(.A(n_62820), .B(n_220956467), .C(n_1730), .Z(n_1731
		));
	notech_nao3 i_1034(.A(axi_WSTRB[1]), .B(n_60760), .C(n_60737), .Z(n_1732
		));
	notech_nand3 i_57191(.A(n_62820), .B(n_220956467), .C(n_1732), .Z(n_1733
		));
	notech_nao3 i_1036(.A(axi_WSTRB[0]), .B(n_60760), .C(n_60737), .Z(n_1734
		));
	notech_nand3 i_57189(.A(n_62820), .B(n_220956467), .C(n_1734), .Z(n_1735
		));
	notech_nao3 i_1038(.A(axi_WSTRB[3]), .B(n_60715), .C(n_60737), .Z(n_1736
		));
	notech_nand3 i_57187(.A(n_62820), .B(n_220956467), .C(n_1736), .Z(n_1737
		));
	notech_nao3 i_1040(.A(axi_WSTRB[2]), .B(n_60715), .C(n_60737), .Z(n_1738
		));
	notech_nand3 i_57185(.A(n_62820), .B(n_220956467), .C(n_1738), .Z(n_1739
		));
	notech_nao3 i_1042(.A(axi_WSTRB[1]), .B(n_60715), .C(n_60737), .Z(n_1740
		));
	notech_nand3 i_57183(.A(n_62820), .B(n_220956467), .C(n_1740), .Z(n_1741
		));
	notech_ao3 i_123(.A(fsm[4]), .B(fsm[2]), .C(n_1998), .Z(n_1742));
	notech_nand2 i_1044(.A(n_2049), .B(n_2050), .Z(n_1743));
	notech_ao3 i_58707(.A(n_2070), .B(n_1743), .C(n_1742), .Z(n_1744));
	notech_nao3 i_1047(.A(axi_WSTRB[0]), .B(n_60715), .C(n_60737), .Z(n_1745
		));
	notech_nand3 i_57181(.A(n_62820), .B(n_220956467), .C(n_1745), .Z(n_1746
		));
	notech_nand3 i_1050(.A(axi_RVALID), .B(axi_RLAST), .C(n_62132), .Z(n_1747
		));
	notech_and4 i_1051(.A(axi_AWREADY), .B(axi_AWVALID), .C(n_2037), .D(n_25047
		), .Z(n_1748));
	notech_ao3 i_57840(.A(n_62793), .B(n_1747), .C(n_221656474), .Z(n_1749)
		);
	notech_and2 i_1061(.A(n_2041), .B(n_2033), .Z(n_1750));
	notech_or4 i_57216(.A(n_1221), .B(n_974), .C(n_1750), .D(n_8224), .Z(n_1751
		));
	notech_nand2 i_1066(.A(axi_ARREADY), .B(n_8215), .Z(n_1754));
	notech_and4 i_59029(.A(n_2064), .B(n_62793), .C(n_973), .D(n_1754), .Z(n_1755
		));
	notech_nand2 i_57221(.A(n_62161), .B(n_221956477), .Z(n_1756));
	notech_nand2 i_1072(.A(axi_ARREADY), .B(n_1758), .Z(n_1757));
	notech_nand3 i_128(.A(n_2045), .B(n_8265), .C(n_62123), .Z(n_1758));
	notech_and4 i_58995(.A(n_62161), .B(n_1743), .C(n_2022), .D(n_1757), .Z(n_1759
		));
	notech_nand2 i_56157(.A(n_62161), .B(n_2019), .Z(n_1760));
	notech_ao4 i_69(.A(n_222656484), .B(n_222556483), .C(n_222456482), .D(n_8333
		), .Z(n_1763));
	notech_ao4 i_57618(.A(n_223056488), .B(n_223356491), .C(n_222756485), .D
		(n_8330), .Z(n_1765));
	notech_ao4 i_57860(.A(n_8219), .B(n_8218), .C(n_222756485), .D(n_8330), 
		.Z(n_1766));
	notech_ao4 i_58525(.A(readio_ack), .B(n_8560), .C(n_222656484), .D(n_222556483
		), .Z(n_1769));
	notech_ao4 i_58980(.A(n_223056488), .B(n_223156489), .C(n_8333), .D(n_222456482
		), .Z(n_1770));
	notech_mux2 i_1(.S(n_2033), .A(Daddr[4]), .B(axi_AW[4]), .Z(cacheA[0])
		);
	notech_mux2 i_211482(.S(n_2033), .A(Daddr[5]), .B(axi_AW[5]), .Z(cacheA[
		1]));
	notech_mux2 i_3(.S(n_2033), .A(Daddr[6]), .B(axi_AW[6]), .Z(cacheA[2])
		);
	notech_mux2 i_4(.S(n_2033), .A(Daddr[7]), .B(axi_AW[7]), .Z(cacheA[3])
		);
	notech_mux2 i_5(.S(n_2033), .A(Daddr[8]), .B(axi_AW[8]), .Z(cacheA[4])
		);
	notech_mux2 i_6(.S(n_2033), .A(Daddr[9]), .B(axi_AW[9]), .Z(cacheA[5])
		);
	notech_mux2 i_7(.S(n_2033), .A(Daddr[10]), .B(axi_AW[10]), .Z(cacheA[6])
		);
	notech_mux2 i_8(.S(n_62170), .A(Daddr[11]), .B(axi_AW[11]), .Z(cacheA[7]
		));
	notech_mux2 i_9(.S(n_62170), .A(Daddr[12]), .B(axi_AW[12]), .Z(cacheA[8]
		));
	notech_mux2 i_10(.S(n_62170), .A(Daddr[13]), .B(axi_AW[13]), .Z(cacheA[9
		]));
	notech_and4 i_1161(.A(n_60789), .B(n_62809), .C(cacheQ[64]), .D(n_60715)
		, .Z(n_1805));
	notech_nao3 i_122015(.A(n_2245), .B(n_2240), .C(n_1805), .Z(read_data[0]
		));
	notech_reg code_wack_reg(.CP(n_63282), .D(n_4740), .CD(n_62726), .Q(code_wack
		));
	notech_mux2 i_2330(.S(n_975), .A(n_25047), .B(code_wack), .Z(n_4740));
	notech_and4 i_1170(.A(A4[1]), .B(n_62809), .C(cacheQ[65]), .D(n_60715), 
		.Z(n_1811));
	notech_reg code_ack_slow_reg(.CP(n_63282), .D(n_4746), .CD(n_62726), .Q(code_ack
		));
	notech_mux2 i_2338(.S(n_977), .A(n_22714), .B(code_ack), .Z(n_4746));
	notech_nao3 i_222016(.A(n_2248), .B(n_2247), .C(n_1811), .Z(read_data[1]
		));
	notech_reg axi_AR_reg_0(.CP(n_63282), .D(n_4755), .CD(n_62726), .Q(axi_AR
		[0]));
	notech_and4 i_2348(.A(n_1066), .B(n_973), .C(axi_AR[0]), .D(n_62793), .Z
		(n_4755));
	notech_reg axi_AR_reg_1(.CP(n_63282), .D(n_4761), .CD(n_62726), .Q(axi_AR
		[1]));
	notech_and4 i_2356(.A(n_62793), .B(n_1066), .C(n_973), .D(axi_AR[1]), .Z
		(n_4761));
	notech_reg axi_AR_reg_2(.CP(n_63282), .D(n_4764), .CD(n_62726), .Q(axi_AR
		[2]));
	notech_mux2 i_2362(.S(n_1067), .A(n_8258), .B(axi_AR[2]), .Z(n_4764));
	notech_reg axi_AR_reg_3(.CP(n_63282), .D(n_4770), .CD(n_62726), .Q(axi_AR
		[3]));
	notech_mux2 i_2370(.S(n_1067), .A(n_8257), .B(axi_AR[3]), .Z(n_4770));
	notech_reg axi_AR_reg_4(.CP(n_63282), .D(n_4776), .CD(n_62726), .Q(axi_AR
		[4]));
	notech_mux2 i_2378(.S(n_1067), .A(n_8256), .B(axi_AR[4]), .Z(n_4776));
	notech_and4 i_1179(.A(A4[1]), .B(n_62809), .C(cacheQ[66]), .D(n_60715), 
		.Z(n_1817));
	notech_reg axi_AR_reg_5(.CP(n_63282), .D(n_4782), .CD(n_62726), .Q(axi_AR
		[5]));
	notech_mux2 i_2386(.S(n_1067), .A(n_8255), .B(axi_AR[5]), .Z(n_4782));
	notech_nao3 i_322017(.A(n_2251), .B(n_2250), .C(n_1817), .Z(read_data[2]
		));
	notech_reg axi_AR_reg_6(.CP(n_63282), .D(n_4788), .CD(n_62724), .Q(axi_AR
		[6]));
	notech_mux2 i_2394(.S(n_1067), .A(n_8254), .B(axi_AR[6]), .Z(n_4788));
	notech_reg axi_AR_reg_7(.CP(n_63282), .D(n_4794), .CD(n_62724), .Q(axi_AR
		[7]));
	notech_mux2 i_2402(.S(n_1067), .A(n_8253), .B(axi_AR[7]), .Z(n_4794));
	notech_reg axi_AR_reg_8(.CP(n_63282), .D(n_4800), .CD(n_62724), .Q(axi_AR
		[8]));
	notech_mux2 i_2410(.S(n_1067), .A(n_8252), .B(axi_AR[8]), .Z(n_4800));
	notech_reg axi_AR_reg_9(.CP(n_63282), .D(n_4806), .CD(n_62724), .Q(axi_AR
		[9]));
	notech_mux2 i_2418(.S(n_1067), .A(n_8251), .B(axi_AR[9]), .Z(n_4806));
	notech_reg axi_AR_reg_10(.CP(n_63282), .D(n_4812), .CD(n_62724), .Q(axi_AR
		[10]));
	notech_mux2 i_2426(.S(n_1067), .A(n_8250), .B(axi_AR[10]), .Z(n_4812));
	notech_and4 i_1188(.A(A4[1]), .B(n_62809), .C(cacheQ[67]), .D(n_60715), 
		.Z(n_1823));
	notech_reg axi_AR_reg_11(.CP(n_63282), .D(n_4818), .CD(n_62724), .Q(axi_AR
		[11]));
	notech_mux2 i_2434(.S(n_1067), .A(n_8249), .B(axi_AR[11]), .Z(n_4818));
	notech_nao3 i_422018(.A(n_2254), .B(n_2253), .C(n_1823), .Z(read_data[3]
		));
	notech_reg axi_AR_reg_12(.CP(n_63282), .D(n_4824), .CD(n_62724), .Q(axi_AR
		[12]));
	notech_mux2 i_2442(.S(n_1067), .A(n_8248), .B(axi_AR[12]), .Z(n_4824));
	notech_reg axi_AR_reg_13(.CP(n_63282), .D(n_4830), .CD(n_62724), .Q(axi_AR
		[13]));
	notech_mux2 i_2450(.S(n_1067), .A(n_8247), .B(axi_AR[13]), .Z(n_4830));
	notech_reg axi_AR_reg_14(.CP(n_63282), .D(n_4836), .CD(n_62726), .Q(axi_AR
		[14]));
	notech_mux2 i_2458(.S(n_1067), .A(n_8246), .B(axi_AR[14]), .Z(n_4836));
	notech_reg axi_AR_reg_15(.CP(n_63282), .D(n_4842), .CD(n_62727), .Q(axi_AR
		[15]));
	notech_mux2 i_2466(.S(n_1067), .A(n_8245), .B(axi_AR[15]), .Z(n_4842));
	notech_reg axi_AR_reg_16(.CP(n_63282), .D(n_4848), .CD(n_62727), .Q(axi_AR
		[16]));
	notech_mux2 i_2474(.S(n_1067), .A(n_8244), .B(axi_AR[16]), .Z(n_4848));
	notech_and4 i_1197(.A(n_60789), .B(n_62809), .C(cacheQ[68]), .D(n_60715)
		, .Z(n_1829));
	notech_reg axi_AR_reg_17(.CP(n_63298), .D(n_4854), .CD(n_62727), .Q(axi_AR
		[17]));
	notech_mux2 i_2482(.S(n_1067), .A(n_8243), .B(axi_AR[17]), .Z(n_4854));
	notech_nao3 i_522019(.A(n_2257), .B(n_2256), .C(n_1829), .Z(read_data[4]
		));
	notech_reg axi_AR_reg_18(.CP(n_63298), .D(n_4860), .CD(n_62727), .Q(axi_AR
		[18]));
	notech_mux2 i_2490(.S(n_62150), .A(n_8242), .B(axi_AR[18]), .Z(n_4860)
		);
	notech_reg axi_AR_reg_19(.CP(n_63298), .D(n_4866), .CD(n_62727), .Q(axi_AR
		[19]));
	notech_mux2 i_2498(.S(n_62150), .A(n_8241), .B(axi_AR[19]), .Z(n_4866)
		);
	notech_reg axi_AR_reg_20(.CP(n_63298), .D(n_4872), .CD(n_62727), .Q(axi_AR
		[20]));
	notech_mux2 i_2506(.S(n_62150), .A(n_8240), .B(axi_AR[20]), .Z(n_4872)
		);
	notech_reg axi_AR_reg_21(.CP(n_63298), .D(n_4878), .CD(n_62727), .Q(axi_AR
		[21]));
	notech_mux2 i_2514(.S(n_62150), .A(n_8239), .B(axi_AR[21]), .Z(n_4878)
		);
	notech_reg axi_AR_reg_22(.CP(n_63298), .D(n_4884), .CD(n_62727), .Q(axi_AR
		[22]));
	notech_mux2 i_2522(.S(n_62150), .A(n_8238), .B(axi_AR[22]), .Z(n_4884)
		);
	notech_and4 i_1206(.A(n_60789), .B(n_62809), .C(cacheQ[69]), .D(n_60715)
		, .Z(n_1835));
	notech_reg axi_AR_reg_23(.CP(n_63298), .D(n_4890), .CD(n_62726), .Q(axi_AR
		[23]));
	notech_mux2 i_2530(.S(n_62150), .A(n_8237), .B(axi_AR[23]), .Z(n_4890)
		);
	notech_nao3 i_622020(.A(n_2260), .B(n_2259), .C(n_1835), .Z(read_data[5]
		));
	notech_reg axi_AR_reg_24(.CP(n_63298), .D(n_4896), .CD(n_62726), .Q(axi_AR
		[24]));
	notech_mux2 i_2538(.S(n_62150), .A(n_8236), .B(axi_AR[24]), .Z(n_4896)
		);
	notech_reg axi_AR_reg_25(.CP(n_63298), .D(n_4902), .CD(n_62726), .Q(axi_AR
		[25]));
	notech_mux2 i_2546(.S(n_62150), .A(n_8235), .B(axi_AR[25]), .Z(n_4902)
		);
	notech_reg axi_AR_reg_26(.CP(n_63298), .D(n_4908), .CD(n_62726), .Q(axi_AR
		[26]));
	notech_mux2 i_2554(.S(n_62150), .A(n_8234), .B(axi_AR[26]), .Z(n_4908)
		);
	notech_reg axi_AR_reg_27(.CP(n_63298), .D(n_4914), .CD(n_62727), .Q(axi_AR
		[27]));
	notech_mux2 i_2562(.S(n_62150), .A(n_8232), .B(axi_AR[27]), .Z(n_4914)
		);
	notech_reg axi_AR_reg_28(.CP(n_63298), .D(n_4920), .CD(n_62727), .Q(axi_AR
		[28]));
	notech_mux2 i_2570(.S(n_62150), .A(n_8231), .B(axi_AR[28]), .Z(n_4920)
		);
	notech_and4 i_1215(.A(n_60789), .B(n_62809), .C(cacheQ[70]), .D(n_60715)
		, .Z(n_1841));
	notech_reg axi_AR_reg_29(.CP(n_63298), .D(n_4926), .CD(n_62726), .Q(axi_AR
		[29]));
	notech_mux2 i_2578(.S(n_62150), .A(n_8230), .B(axi_AR[29]), .Z(n_4926)
		);
	notech_nao3 i_722021(.A(n_2263), .B(n_2262), .C(n_1841), .Z(read_data[6]
		));
	notech_reg axi_AR_reg_30(.CP(n_63298), .D(n_4932), .CD(n_62726), .Q(axi_AR
		[30]));
	notech_mux2 i_2586(.S(n_62150), .A(n_8228), .B(axi_AR[30]), .Z(n_4932)
		);
	notech_reg axi_AR_reg_31(.CP(n_63298), .D(n_4938), .CD(n_62724), .Q(axi_AR
		[31]));
	notech_mux2 i_2594(.S(n_62150), .A(n_8227), .B(axi_AR[31]), .Z(n_4938)
		);
	notech_reg axi_AW_reg_0(.CP(n_63298), .D(n_4947), .CD(n_62722), .Q(axi_AW
		[0]));
	notech_and4 i_2604(.A(n_62793), .B(n_8323), .C(n_62820), .D(axi_AW[0]), 
		.Z(n_4947));
	notech_reg axi_AW_reg_1(.CP(n_63298), .D(n_4953), .CD(n_62722), .Q(axi_AW
		[1]));
	notech_and4 i_2612(.A(n_62793), .B(n_8323), .C(n_62820), .D(axi_AW[1]), 
		.Z(n_4953));
	notech_reg axi_AW_reg_2(.CP(n_63298), .D(n_4956), .CD(n_62722), .Q(axi_AW
		[2]));
	notech_mux2 i_2618(.S(n_62782), .A(n_8289), .B(axi_AW[2]), .Z(n_4956));
	notech_and4 i_1224(.A(n_60789), .B(n_62809), .C(cacheQ[71]), .D(n_60715)
		, .Z(n_1847));
	notech_reg axi_AW_reg_3(.CP(n_63298), .D(n_4962), .CD(n_62722), .Q(axi_AW
		[3]));
	notech_mux2 i_2626(.S(n_62782), .A(n_8288), .B(axi_AW[3]), .Z(n_4962));
	notech_nao3 i_822022(.A(n_2266), .B(n_2265), .C(n_1847), .Z(read_data[7]
		));
	notech_reg axi_AW_reg_4(.CP(n_63344), .D(n_4968), .CD(n_62723), .Q(axi_AW
		[4]));
	notech_mux2 i_2634(.S(n_62782), .A(n_8287), .B(axi_AW[4]), .Z(n_4968));
	notech_reg axi_AW_reg_5(.CP(n_63296), .D(n_4974), .CD(n_62723), .Q(axi_AW
		[5]));
	notech_mux2 i_2642(.S(n_62782), .A(n_8286), .B(axi_AW[5]), .Z(n_4974));
	notech_reg axi_AW_reg_6(.CP(n_63344), .D(n_4980), .CD(n_62723), .Q(axi_AW
		[6]));
	notech_mux2 i_2650(.S(n_62782), .A(n_8285), .B(axi_AW[6]), .Z(n_4980));
	notech_reg axi_AW_reg_7(.CP(n_63344), .D(n_4986), .CD(n_62723), .Q(axi_AW
		[7]));
	notech_mux2 i_2658(.S(n_62782), .A(n_8284), .B(axi_AW[7]), .Z(n_4986));
	notech_reg axi_AW_reg_8(.CP(n_63344), .D(n_4992), .CD(n_62722), .Q(axi_AW
		[8]));
	notech_mux2 i_2666(.S(n_62782), .A(n_8283), .B(axi_AW[8]), .Z(n_4992));
	notech_and4 i_1233(.A(n_60789), .B(n_62809), .C(cacheQ[72]), .D(n_60717)
		, .Z(n_1853));
	notech_reg axi_AW_reg_9(.CP(n_63344), .D(n_4998), .CD(n_62722), .Q(axi_AW
		[9]));
	notech_mux2 i_2674(.S(n_62782), .A(n_8282), .B(axi_AW[9]), .Z(n_4998));
	notech_nao3 i_922023(.A(n_2269), .B(n_2268), .C(n_1853), .Z(read_data[8]
		));
	notech_reg axi_AW_reg_10(.CP(n_63344), .D(n_5004), .CD(n_62722), .Q(axi_AW
		[10]));
	notech_mux2 i_2682(.S(n_62782), .A(n_8281), .B(axi_AW[10]), .Z(n_5004)
		);
	notech_reg axi_AW_reg_11(.CP(n_63344), .D(n_5010), .CD(n_62722), .Q(axi_AW
		[11]));
	notech_mux2 i_2690(.S(n_62782), .A(n_8280), .B(axi_AW[11]), .Z(n_5010)
		);
	notech_reg axi_AW_reg_12(.CP(n_63344), .D(n_5016), .CD(n_62722), .Q(axi_AW
		[12]));
	notech_mux2 i_2698(.S(n_62782), .A(n_8279), .B(axi_AW[12]), .Z(n_5016)
		);
	notech_reg axi_AW_reg_13(.CP(n_63344), .D(n_5022), .CD(n_62722), .Q(axi_AW
		[13]));
	notech_mux2 i_2706(.S(n_62782), .A(n_8278), .B(axi_AW[13]), .Z(n_5022)
		);
	notech_reg axi_AW_reg_14(.CP(n_63344), .D(n_5028), .CD(n_62722), .Q(axi_AW
		[14]));
	notech_mux2 i_2714(.S(n_62782), .A(n_8277), .B(axi_AW[14]), .Z(n_5028)
		);
	notech_and4 i_1242(.A(A4[1]), .B(n_62809), .C(cacheQ[73]), .D(n_60720), 
		.Z(n_1859));
	notech_reg axi_AW_reg_15(.CP(n_63344), .D(n_5034), .CD(n_62722), .Q(axi_AW
		[15]));
	notech_mux2 i_2722(.S(n_62783), .A(n_8276), .B(axi_AW[15]), .Z(n_5034)
		);
	notech_nao3 i_1022024(.A(n_2272), .B(n_2271), .C(n_1859), .Z(read_data[9
		]));
	notech_reg axi_AW_reg_16(.CP(n_63344), .D(n_5040), .CD(n_62723), .Q(axi_AW
		[16]));
	notech_mux2 i_2730(.S(n_62783), .A(n_8275), .B(axi_AW[16]), .Z(n_5040)
		);
	notech_reg axi_AW_reg_17(.CP(n_63344), .D(n_5046), .CD(n_62724), .Q(axi_AW
		[17]));
	notech_mux2 i_2738(.S(n_62783), .A(n_8274), .B(axi_AW[17]), .Z(n_5046)
		);
	notech_reg axi_AW_reg_18(.CP(n_63344), .D(n_5052), .CD(n_62724), .Q(axi_AW
		[18]));
	notech_mux2 i_2746(.S(n_62783), .A(n_8273), .B(axi_AW[18]), .Z(n_5052)
		);
	notech_reg axi_AW_reg_19(.CP(n_63344), .D(n_5058), .CD(n_62723), .Q(axi_AW
		[19]));
	notech_mux2 i_2754(.S(n_62783), .A(n_8272), .B(axi_AW[19]), .Z(n_5058)
		);
	notech_reg axi_AW_reg_20(.CP(n_63344), .D(n_5064), .CD(n_62723), .Q(axi_AW
		[20]));
	notech_mux2 i_2762(.S(n_62783), .A(n_8271), .B(axi_AW[20]), .Z(n_5064)
		);
	notech_and4 i_1251(.A(A4[1]), .B(n_62809), .C(cacheQ[74]), .D(n_60720), 
		.Z(n_1865));
	notech_reg axi_AW_reg_21(.CP(n_63344), .D(n_5070), .CD(n_62724), .Q(axi_AW
		[21]));
	notech_mux2 i_2770(.S(n_62783), .A(n_8270), .B(axi_AW[21]), .Z(n_5070)
		);
	notech_nao3 i_1122025(.A(n_2275), .B(n_2274), .C(n_1865), .Z(read_data[
		10]));
	notech_reg axi_AW_reg_22(.CP(n_63344), .D(n_5076), .CD(n_62724), .Q(axi_AW
		[22]));
	notech_mux2 i_2778(.S(n_62783), .A(n_8269), .B(axi_AW[22]), .Z(n_5076)
		);
	notech_reg axi_AW_reg_23(.CP(n_63322), .D(n_5082), .CD(n_62724), .Q(axi_AW
		[23]));
	notech_mux2 i_2786(.S(n_62783), .A(n_8268), .B(axi_AW[23]), .Z(n_5082)
		);
	notech_reg axi_AW_reg_24(.CP(n_63296), .D(n_5088), .CD(n_62724), .Q(axi_AW
		[24]));
	notech_mux2 i_2794(.S(n_62783), .A(n_8267), .B(axi_AW[24]), .Z(n_5088)
		);
	notech_reg axi_AW_reg_25(.CP(n_63296), .D(n_5094), .CD(n_62723), .Q(axi_AW
		[25]));
	notech_mux2 i_2802(.S(n_62783), .A(n_8266), .B(axi_AW[25]), .Z(n_5094)
		);
	notech_reg axi_AW_reg_26(.CP(n_63296), .D(n_5100), .CD(n_62723), .Q(axi_AW
		[26]));
	notech_mux2 i_2810(.S(n_62783), .A(n_8264), .B(axi_AW[26]), .Z(n_5100)
		);
	notech_and4 i_1260(.A(A4[1]), .B(n_62809), .C(cacheQ[75]), .D(n_60720), 
		.Z(n_1871));
	notech_reg axi_AW_reg_27(.CP(n_63296), .D(n_5106), .CD(n_62723), .Q(axi_AW
		[27]));
	notech_mux2 i_2818(.S(n_62783), .A(n_8263), .B(axi_AW[27]), .Z(n_5106)
		);
	notech_nao3 i_1222026(.A(n_2278), .B(n_2277), .C(n_1871), .Z(read_data[
		11]));
	notech_reg axi_AW_reg_28(.CP(n_63296), .D(n_5112), .CD(n_62723), .Q(axi_AW
		[28]));
	notech_mux2 i_2826(.S(n_62783), .A(n_8262), .B(axi_AW[28]), .Z(n_5112)
		);
	notech_reg axi_AW_reg_29(.CP(n_63296), .D(n_5118), .CD(n_62723), .Q(axi_AW
		[29]));
	notech_mux2 i_2834(.S(n_62783), .A(n_8261), .B(axi_AW[29]), .Z(n_5118)
		);
	notech_reg axi_AW_reg_30(.CP(n_63296), .D(n_5124), .CD(n_62723), .Q(axi_AW
		[30]));
	notech_mux2 i_2842(.S(n_62783), .A(n_8260), .B(axi_AW[30]), .Z(n_5124)
		);
	notech_reg axi_AW_reg_31(.CP(n_63296), .D(n_5130), .CD(n_62723), .Q(axi_AW
		[31]));
	notech_mux2 i_2850(.S(n_62783), .A(n_8259), .B(axi_AW[31]), .Z(n_5130)
		);
	notech_reg_set burst_idx_reg_0(.CP(n_63296), .D(n_5136), .SD(1'b1), .Q(burst_idx
		[0]));
	notech_mux2 i_2858(.S(n_1171), .A(n_8290), .B(burst_idx[0]), .Z(n_5136)
		);
	notech_and4 i_1269(.A(A4[1]), .B(n_62809), .C(cacheQ[76]), .D(n_60720), 
		.Z(n_1877));
	notech_reg_set burst_idx_reg_1(.CP(n_63296), .D(n_5142), .SD(1'b1), .Q(burst_idx
		[1]));
	notech_mux2 i_2866(.S(n_1171), .A(n_25495), .B(burst_idx[1]), .Z(n_5142)
		);
	notech_nao3 i_1322027(.A(n_2281), .B(n_2280), .C(n_1877), .Z(read_data[
		12]));
	notech_reg_set burst_idx_reg_2(.CP(n_63296), .D(n_5148), .SD(1'b1), .Q(burst_idx
		[2]));
	notech_mux2 i_2874(.S(n_1171), .A(n_25500), .B(burst_idx[2]), .Z(n_5148)
		);
	notech_reg_set burst_idx_reg_3(.CP(n_63296), .D(n_5154), .SD(1'b1), .Q(burst_idx
		[3]));
	notech_mux2 i_2882(.S(n_1171), .A(n_25505), .B(burst_idx[3]), .Z(n_5154)
		);
	notech_reg_set burst_idx_reg_4(.CP(n_63296), .D(n_5160), .SD(1'b1), .Q(burst_idx
		[4]));
	notech_mux2 i_2890(.S(n_1171), .A(n_25510), .B(burst_idx[4]), .Z(n_5160)
		);
	notech_reg axi_AWVALID_reg(.CP(n_63296), .D(n_5166), .CD(n_62723), .Q(axi_AWVALID
		));
	notech_mux2 i_2898(.S(n_1175), .A(n_1176), .B(axi_AWVALID), .Z(n_5166)
		);
	notech_reg_set A4_reg_0(.CP(n_63296), .D(n_5172), .SD(1'b1), .Q(A4[0])
		);
	notech_mux2 i_2906(.S(\nbus_11672[0] ), .A(n_60760), .B(Daddr[2]), .Z(n_5172
		));
	notech_and4 i_1278(.A(A4[1]), .B(n_62809), .C(cacheQ[77]), .D(n_60720), 
		.Z(n_1883));
	notech_reg_set A4_reg_1(.CP(n_63296), .D(n_5178), .SD(1'b1), .Q(A4[1])
		);
	notech_mux2 i_2914(.S(\nbus_11672[0] ), .A(A4[1]), .B(Daddr[3]), .Z(n_5178
		));
	notech_nao3 i_1422028(.A(n_2284), .B(n_2283), .C(n_1883), .Z(read_data[
		13]));
	notech_reg axi_W_reg_0(.CP(n_63296), .D(n_5184), .CD(n_62730), .Q(axi_W[
		0]));
	notech_mux2 i_2922(.S(n_62783), .A(n_8298), .B(axi_W[0]), .Z(n_5184));
	notech_reg axi_W_reg_1(.CP(n_63296), .D(n_5190), .CD(n_62730), .Q(axi_W[
		1]));
	notech_mux2 i_2930(.S(n_62782), .A(n_8297), .B(axi_W[1]), .Z(n_5190));
	notech_reg axi_W_reg_2(.CP(n_63344), .D(n_5196), .CD(n_62730), .Q(axi_W[
		2]));
	notech_mux2 i_2938(.S(n_62772), .A(n_8296), .B(axi_W[2]), .Z(n_5196));
	notech_reg axi_W_reg_3(.CP(n_63318), .D(n_5202), .CD(n_62730), .Q(axi_W[
		3]));
	notech_mux2 i_2946(.S(n_62772), .A(n_8295), .B(axi_W[3]), .Z(n_5202));
	notech_reg axi_W_reg_4(.CP(n_63294), .D(n_5208), .CD(n_62730), .Q(axi_W[
		4]));
	notech_mux2 i_2954(.S(n_62772), .A(n_8294), .B(axi_W[4]), .Z(n_5208));
	notech_and4 i_1287(.A(A4[1]), .B(n_62809), .C(cacheQ[78]), .D(n_60720), 
		.Z(n_1889));
	notech_reg axi_W_reg_5(.CP(n_63318), .D(n_5214), .CD(n_62730), .Q(axi_W[
		5]));
	notech_mux2 i_2962(.S(n_62772), .A(n_8293), .B(axi_W[5]), .Z(n_5214));
	notech_nao3 i_1522029(.A(n_2287), .B(n_2286), .C(n_1889), .Z(read_data[
		14]));
	notech_reg axi_W_reg_6(.CP(n_63318), .D(n_5220), .CD(n_62730), .Q(axi_W[
		6]));
	notech_mux2 i_2970(.S(n_62772), .A(n_8292), .B(axi_W[6]), .Z(n_5220));
	notech_reg axi_W_reg_7(.CP(n_63318), .D(n_5226), .CD(n_62730), .Q(axi_W[
		7]));
	notech_mux2 i_2978(.S(n_62772), .A(n_8291), .B(axi_W[7]), .Z(n_5226));
	notech_reg axi_W_reg_8(.CP(n_63318), .D(n_5232), .CD(n_62730), .Q(axi_W[
		8]));
	notech_mux2 i_2986(.S(n_62772), .A(n_24828), .B(axi_W[8]), .Z(n_5232));
	notech_reg axi_W_reg_9(.CP(n_63318), .D(n_5238), .CD(n_62730), .Q(axi_W[
		9]));
	notech_mux2 i_2994(.S(n_62772), .A(n_24834), .B(axi_W[9]), .Z(n_5238));
	notech_reg axi_W_reg_10(.CP(n_63318), .D(n_5244), .CD(n_62729), .Q(axi_W
		[10]));
	notech_mux2 i_3002(.S(n_62772), .A(n_24840), .B(axi_W[10]), .Z(n_5244)
		);
	notech_and4 i_1296(.A(A4[1]), .B(n_62809), .C(cacheQ[79]), .D(n_60720), 
		.Z(n_1895));
	notech_reg axi_W_reg_11(.CP(n_63318), .D(n_5250), .CD(n_62730), .Q(axi_W
		[11]));
	notech_mux2 i_3010(.S(n_62772), .A(n_24846), .B(axi_W[11]), .Z(n_5250)
		);
	notech_nao3 i_1622030(.A(n_2290), .B(n_2289), .C(n_1895), .Z(read_data[
		15]));
	notech_reg axi_W_reg_12(.CP(n_63318), .D(n_5256), .CD(n_62730), .Q(axi_W
		[12]));
	notech_mux2 i_3018(.S(n_62772), .A(n_24852), .B(axi_W[12]), .Z(n_5256)
		);
	notech_reg axi_W_reg_13(.CP(n_63318), .D(n_5262), .CD(n_62730), .Q(axi_W
		[13]));
	notech_mux2 i_3026(.S(n_62772), .A(n_24858), .B(axi_W[13]), .Z(n_5262)
		);
	notech_reg axi_W_reg_14(.CP(n_63318), .D(n_5268), .CD(n_62730), .Q(axi_W
		[14]));
	notech_mux2 i_3034(.S(n_62772), .A(n_24864), .B(axi_W[14]), .Z(n_5268)
		);
	notech_reg axi_W_reg_15(.CP(n_63318), .D(n_5274), .CD(n_62730), .Q(axi_W
		[15]));
	notech_mux2 i_3042(.S(n_62772), .A(n_24870), .B(axi_W[15]), .Z(n_5274)
		);
	notech_reg axi_W_reg_16(.CP(n_63318), .D(n_5280), .CD(n_62730), .Q(axi_W
		[16]));
	notech_mux2 i_3050(.S(n_62772), .A(n_24876), .B(axi_W[16]), .Z(n_5280)
		);
	notech_and4 i_1305(.A(A4[1]), .B(n_62810), .C(cacheQ[80]), .D(n_60720), 
		.Z(n_1901));
	notech_reg axi_W_reg_17(.CP(n_63318), .D(n_5286), .CD(n_62731), .Q(axi_W
		[17]));
	notech_mux2 i_3058(.S(n_62772), .A(n_24882), .B(axi_W[17]), .Z(n_5286)
		);
	notech_nao3 i_1722031(.A(n_2293), .B(n_2292), .C(n_1901), .Z(read_data[
		16]));
	notech_reg axi_W_reg_18(.CP(n_63318), .D(n_5292), .CD(n_62731), .Q(axi_W
		[18]));
	notech_mux2 i_3066(.S(n_62772), .A(n_24888), .B(axi_W[18]), .Z(n_5292)
		);
	notech_reg axi_W_reg_19(.CP(n_63318), .D(n_5298), .CD(n_62731), .Q(axi_W
		[19]));
	notech_mux2 i_3074(.S(n_62777), .A(n_24894), .B(axi_W[19]), .Z(n_5298)
		);
	notech_reg axi_W_reg_20(.CP(n_63318), .D(n_5304), .CD(n_62731), .Q(axi_W
		[20]));
	notech_mux2 i_3082(.S(n_62777), .A(n_24900), .B(axi_W[20]), .Z(n_5304)
		);
	notech_reg axi_W_reg_21(.CP(n_63318), .D(n_5310), .CD(n_62731), .Q(axi_W
		[21]));
	notech_mux2 i_3090(.S(n_62777), .A(n_24906), .B(axi_W[21]), .Z(n_5310)
		);
	notech_reg axi_W_reg_22(.CP(n_63354), .D(n_5316), .CD(n_62731), .Q(axi_W
		[22]));
	notech_mux2 i_3098(.S(n_62777), .A(n_24912), .B(axi_W[22]), .Z(n_5316)
		);
	notech_and4 i_1314(.A(A4[1]), .B(n_62810), .C(cacheQ[81]), .D(n_60720), 
		.Z(n_1907));
	notech_reg axi_W_reg_23(.CP(n_63340), .D(n_5322), .CD(n_62731), .Q(axi_W
		[23]));
	notech_mux2 i_3106(.S(n_62777), .A(n_24918), .B(axi_W[23]), .Z(n_5322)
		);
	notech_nao3 i_1822032(.A(n_2296), .B(n_2295), .C(n_1907), .Z(read_data[
		17]));
	notech_reg axi_W_reg_24(.CP(n_63354), .D(n_5328), .CD(n_62731), .Q(axi_W
		[24]));
	notech_mux2 i_3114(.S(n_62777), .A(n_24924), .B(axi_W[24]), .Z(n_5328)
		);
	notech_reg axi_W_reg_25(.CP(n_63354), .D(n_5334), .CD(n_62731), .Q(axi_W
		[25]));
	notech_mux2 i_3122(.S(n_62777), .A(n_24930), .B(axi_W[25]), .Z(n_5334)
		);
	notech_reg axi_W_reg_26(.CP(n_63354), .D(n_5340), .CD(n_62731), .Q(axi_W
		[26]));
	notech_mux2 i_3130(.S(n_62777), .A(n_24936), .B(axi_W[26]), .Z(n_5340)
		);
	notech_reg axi_W_reg_27(.CP(n_63354), .D(n_5346), .CD(n_62731), .Q(axi_W
		[27]));
	notech_mux2 i_3138(.S(n_62777), .A(n_24942), .B(axi_W[27]), .Z(n_5346)
		);
	notech_reg axi_W_reg_28(.CP(n_63354), .D(n_5352), .CD(n_62731), .Q(axi_W
		[28]));
	notech_mux2 i_3146(.S(n_62777), .A(n_24948), .B(axi_W[28]), .Z(n_5352)
		);
	notech_and4 i_1323(.A(A4[1]), .B(n_62810), .C(cacheQ[82]), .D(n_60720), 
		.Z(n_1913));
	notech_reg axi_W_reg_29(.CP(n_63354), .D(n_5358), .CD(n_62731), .Q(axi_W
		[29]));
	notech_mux2 i_3154(.S(n_62777), .A(n_24954), .B(axi_W[29]), .Z(n_5358)
		);
	notech_nao3 i_1922033(.A(n_2299), .B(n_2298), .C(n_1913), .Z(read_data[
		18]));
	notech_reg axi_W_reg_30(.CP(n_63354), .D(n_5364), .CD(n_62731), .Q(axi_W
		[30]));
	notech_mux2 i_3162(.S(n_62777), .A(n_24960), .B(axi_W[30]), .Z(n_5364)
		);
	notech_reg axi_W_reg_31(.CP(n_63354), .D(n_5370), .CD(n_62731), .Q(axi_W
		[31]));
	notech_mux2 i_3170(.S(n_62777), .A(n_24966), .B(axi_W[31]), .Z(n_5370)
		);
	notech_reg abort_reg(.CP(n_63354), .D(n_5376), .CD(n_62731), .Q(abort)
		);
	notech_mux2 i_3178(.S(n_1203), .A(n_1204), .B(abort), .Z(n_5376));
	notech_reg read_ack_slow_reg(.CP(n_63354), .D(n_5382), .CD(n_62729), .Q(read_ack
		));
	notech_mux2 i_3186(.S(n_1208), .A(n_1210), .B(read_ack), .Z(n_5382));
	notech_reg wrint_ack_reg(.CP(n_63354), .D(n_5388), .CD(n_62728), .Q(write_ack
		));
	notech_mux2 i_3194(.S(n_1211), .A(n_23557), .B(write_ack), .Z(n_5388));
	notech_and4 i_1332(.A(n_60789), .B(n_62810), .C(cacheQ[83]), .D(n_60720)
		, .Z(n_1919));
	notech_reg fsm_reg_0(.CP(n_63354), .D(n_5394), .CD(n_62728), .Q(fsm[0])
		);
	notech_mux2 i_3202(.S(n_1222), .A(n_8301), .B(fsm[0]), .Z(n_5394));
	notech_nao3 i_2022034(.A(n_2302), .B(n_2301), .C(n_1919), .Z(read_data[
		19]));
	notech_reg fsm_reg_1(.CP(n_63354), .D(n_5400), .CD(n_62728), .Q(fsm[1])
		);
	notech_mux2 i_3210(.S(n_1222), .A(n_1216), .B(fsm[1]), .Z(n_5400));
	notech_reg fsm_reg_2(.CP(n_63354), .D(n_5406), .CD(n_62728), .Q(fsm[2])
		);
	notech_mux2 i_3218(.S(n_1222), .A(n_1214), .B(fsm[2]), .Z(n_5406));
	notech_reg fsm_reg_3(.CP(n_63354), .D(n_5412), .CD(n_62728), .Q(fsm[3])
		);
	notech_mux2 i_3226(.S(n_1222), .A(n_8299), .B(fsm[3]), .Z(n_5412));
	notech_reg fsm_reg_4(.CP(n_63354), .D(n_5418), .CD(n_62728), .Q(fsm[4])
		);
	notech_mux2 i_3234(.S(n_1222), .A(n_1212), .B(fsm[4]), .Z(n_5418));
	notech_reg_set cacheD_reg_0(.CP(n_63354), .D(n_5424), .SD(1'b1), .Q(cacheD
		[0]));
	notech_mux2 i_3242(.S(n_1703), .A(n_1708), .B(cacheD[0]), .Z(n_5424));
	notech_and4 i_1341(.A(n_60785), .B(n_62810), .C(cacheQ[84]), .D(n_60720)
		, .Z(n_1925));
	notech_reg_set cacheD_reg_1(.CP(n_63318), .D(n_5430), .SD(1'b1), .Q(cacheD
		[1]));
	notech_mux2 i_3250(.S(n_1703), .A(n_1701), .B(cacheD[1]), .Z(n_5430));
	notech_nao3 i_2122035(.A(n_2305), .B(n_2304), .C(n_1925), .Z(read_data[
		20]));
	notech_reg_set cacheD_reg_2(.CP(n_63354), .D(n_5436), .SD(1'b1), .Q(cacheD
		[2]));
	notech_mux2 i_3258(.S(n_1703), .A(n_1697), .B(cacheD[2]), .Z(n_5436));
	notech_reg_set cacheD_reg_3(.CP(n_63342), .D(n_5442), .SD(1'b1), .Q(cacheD
		[3]));
	notech_mux2 i_3266(.S(n_1703), .A(n_1693), .B(cacheD[3]), .Z(n_5442));
	notech_reg_set cacheD_reg_4(.CP(n_63342), .D(n_5448), .SD(1'b1), .Q(cacheD
		[4]));
	notech_mux2 i_3274(.S(n_1703), .A(n_1689), .B(cacheD[4]), .Z(n_5448));
	notech_reg_set cacheD_reg_5(.CP(n_63342), .D(n_5454), .SD(1'b1), .Q(cacheD
		[5]));
	notech_mux2 i_3282(.S(n_1703), .A(n_1685), .B(cacheD[5]), .Z(n_5454));
	notech_reg_set cacheD_reg_6(.CP(n_63342), .D(n_5460), .SD(1'b1), .Q(cacheD
		[6]));
	notech_mux2 i_3290(.S(n_1703), .A(n_1681), .B(cacheD[6]), .Z(n_5460));
	notech_and4 i_1350(.A(n_60785), .B(n_62810), .C(cacheQ[85]), .D(n_60720)
		, .Z(n_1931));
	notech_reg_set cacheD_reg_7(.CP(n_63342), .D(n_5466), .SD(1'b1), .Q(cacheD
		[7]));
	notech_mux2 i_3298(.S(n_1703), .A(n_1677), .B(cacheD[7]), .Z(n_5466));
	notech_nao3 i_2222036(.A(n_2308), .B(n_2307), .C(n_1931), .Z(read_data[
		21]));
	notech_reg_set cacheD_reg_8(.CP(n_63342), .D(n_5472), .SD(1'b1), .Q(cacheD
		[8]));
	notech_mux2 i_3306(.S(n_1703), .A(n_1673), .B(cacheD[8]), .Z(n_5472));
	notech_reg_set cacheD_reg_9(.CP(n_63342), .D(n_5478), .SD(1'b1), .Q(cacheD
		[9]));
	notech_mux2 i_3314(.S(n_1703), .A(n_1669), .B(cacheD[9]), .Z(n_5478));
	notech_reg_set cacheD_reg_10(.CP(n_63342), .D(n_5484), .SD(1'b1), .Q(cacheD
		[10]));
	notech_mux2 i_3322(.S(n_1703), .A(n_1665), .B(cacheD[10]), .Z(n_5484));
	notech_reg_set cacheD_reg_11(.CP(n_63342), .D(n_5490), .SD(1'b1), .Q(cacheD
		[11]));
	notech_mux2 i_3330(.S(n_1703), .A(n_1661), .B(cacheD[11]), .Z(n_5490));
	notech_reg_set cacheD_reg_12(.CP(n_63342), .D(n_5496), .SD(1'b1), .Q(cacheD
		[12]));
	notech_mux2 i_3338(.S(n_1703), .A(n_1657), .B(cacheD[12]), .Z(n_5496));
	notech_and4 i_1359(.A(n_60785), .B(n_62810), .C(cacheQ[86]), .D(n_60717)
		, .Z(n_1937));
	notech_reg_set cacheD_reg_13(.CP(n_63342), .D(n_5502), .SD(1'b1), .Q(cacheD
		[13]));
	notech_mux2 i_3346(.S(n_1703), .A(n_1653), .B(cacheD[13]), .Z(n_5502));
	notech_nao3 i_2322037(.A(n_2311), .B(n_2310), .C(n_1937), .Z(read_data[
		22]));
	notech_reg_set cacheD_reg_14(.CP(n_63342), .D(n_5508), .SD(1'b1), .Q(cacheD
		[14]));
	notech_mux2 i_3354(.S(n_1703), .A(n_1649), .B(cacheD[14]), .Z(n_5508));
	notech_reg_set cacheD_reg_15(.CP(n_63342), .D(n_5514), .SD(1'b1), .Q(cacheD
		[15]));
	notech_mux2 i_3362(.S(n_1703), .A(n_1645), .B(cacheD[15]), .Z(n_5514));
	notech_reg_set cacheD_reg_16(.CP(n_63342), .D(n_5520), .SD(1'b1), .Q(cacheD
		[16]));
	notech_mux2 i_3370(.S(n_60649), .A(n_1641), .B(cacheD[16]), .Z(n_5520)
		);
	notech_reg_set cacheD_reg_17(.CP(n_63342), .D(n_5526), .SD(1'b1), .Q(cacheD
		[17]));
	notech_mux2 i_3378(.S(n_60649), .A(n_1637), .B(cacheD[17]), .Z(n_5526)
		);
	notech_reg_set cacheD_reg_18(.CP(n_63342), .D(n_5532), .SD(1'b1), .Q(cacheD
		[18]));
	notech_mux2 i_3386(.S(n_60649), .A(n_1633), .B(cacheD[18]), .Z(n_5532)
		);
	notech_and4 i_1368(.A(n_60789), .B(n_62810), .C(cacheQ[87]), .D(n_60717)
		, .Z(n_1943));
	notech_reg_set cacheD_reg_19(.CP(n_63342), .D(n_5538), .SD(1'b1), .Q(cacheD
		[19]));
	notech_mux2 i_3394(.S(n_60649), .A(n_1629), .B(cacheD[19]), .Z(n_5538)
		);
	notech_nao3 i_2422038(.A(n_2314), .B(n_2313), .C(n_1943), .Z(read_data[
		23]));
	notech_reg_set cacheD_reg_20(.CP(n_63342), .D(n_5544), .SD(1'b1), .Q(cacheD
		[20]));
	notech_mux2 i_3402(.S(n_60649), .A(n_1625), .B(cacheD[20]), .Z(n_5544)
		);
	notech_reg_set cacheD_reg_21(.CP(n_63320), .D(n_5550), .SD(1'b1), .Q(cacheD
		[21]));
	notech_mux2 i_3410(.S(n_60649), .A(n_1621), .B(cacheD[21]), .Z(n_5550)
		);
	notech_reg_set cacheD_reg_22(.CP(n_63294), .D(n_5556), .SD(1'b1), .Q(cacheD
		[22]));
	notech_mux2 i_3418(.S(n_60649), .A(n_1617), .B(cacheD[22]), .Z(n_5556)
		);
	notech_reg_set cacheD_reg_23(.CP(n_63294), .D(n_5562), .SD(1'b1), .Q(cacheD
		[23]));
	notech_mux2 i_3426(.S(n_60649), .A(n_1613), .B(cacheD[23]), .Z(n_5562)
		);
	notech_reg_set cacheD_reg_24(.CP(n_63294), .D(n_5568), .SD(1'b1), .Q(cacheD
		[24]));
	notech_mux2 i_3434(.S(n_60649), .A(n_1609), .B(cacheD[24]), .Z(n_5568)
		);
	notech_and4 i_1377(.A(n_60789), .B(n_62810), .C(cacheQ[88]), .D(n_60717)
		, .Z(n_1949));
	notech_reg_set cacheD_reg_25(.CP(n_63294), .D(n_5574), .SD(1'b1), .Q(cacheD
		[25]));
	notech_mux2 i_3442(.S(n_60649), .A(n_1605), .B(cacheD[25]), .Z(n_5574)
		);
	notech_nao3 i_2522039(.A(n_2317), .B(n_2316), .C(n_1949), .Z(read_data[
		24]));
	notech_reg_set cacheD_reg_26(.CP(n_63294), .D(n_5580), .SD(1'b1), .Q(cacheD
		[26]));
	notech_mux2 i_3450(.S(n_60649), .A(n_1601), .B(cacheD[26]), .Z(n_5580)
		);
	notech_reg_set cacheD_reg_27(.CP(n_63294), .D(n_5586), .SD(1'b1), .Q(cacheD
		[27]));
	notech_mux2 i_3458(.S(n_60649), .A(n_1597), .B(cacheD[27]), .Z(n_5586)
		);
	notech_reg_set cacheD_reg_28(.CP(n_63294), .D(n_5592), .SD(1'b1), .Q(cacheD
		[28]));
	notech_mux2 i_3466(.S(n_60649), .A(n_1593), .B(cacheD[28]), .Z(n_5592)
		);
	notech_reg_set cacheD_reg_29(.CP(n_63294), .D(n_5598), .SD(1'b1), .Q(cacheD
		[29]));
	notech_mux2 i_3474(.S(n_60649), .A(n_1589), .B(cacheD[29]), .Z(n_5598)
		);
	notech_reg_set cacheD_reg_30(.CP(n_63294), .D(n_5604), .SD(1'b1), .Q(cacheD
		[30]));
	notech_mux2 i_3482(.S(n_60649), .A(n_1585), .B(cacheD[30]), .Z(n_5604)
		);
	notech_and4 i_1386(.A(n_60785), .B(n_62810), .C(cacheQ[89]), .D(n_60717)
		, .Z(n_1955));
	notech_reg_set cacheD_reg_31(.CP(n_63294), .D(n_5610), .SD(1'b1), .Q(cacheD
		[31]));
	notech_mux2 i_3490(.S(n_60649), .A(n_1581), .B(cacheD[31]), .Z(n_5610)
		);
	notech_nao3 i_2622040(.A(n_2320), .B(n_2319), .C(n_1955), .Z(read_data[
		25]));
	notech_reg_set cacheD_reg_32(.CP(n_63294), .D(n_5616), .SD(1'b1), .Q(cacheD
		[32]));
	notech_mux2 i_3498(.S(n_1573), .A(n_1577), .B(cacheD[32]), .Z(n_5616));
	notech_reg_set cacheD_reg_33(.CP(n_63294), .D(n_5622), .SD(1'b1), .Q(cacheD
		[33]));
	notech_mux2 i_3506(.S(n_1573), .A(n_1571), .B(cacheD[33]), .Z(n_5622));
	notech_reg_set cacheD_reg_34(.CP(n_63294), .D(n_5628), .SD(1'b1), .Q(cacheD
		[34]));
	notech_mux2 i_3514(.S(n_1573), .A(n_1568), .B(cacheD[34]), .Z(n_5628));
	notech_reg_set cacheD_reg_35(.CP(n_63294), .D(n_5634), .SD(1'b1), .Q(cacheD
		[35]));
	notech_mux2 i_3522(.S(n_1573), .A(n_1565), .B(cacheD[35]), .Z(n_5634));
	notech_reg_set cacheD_reg_36(.CP(n_63294), .D(n_5640), .SD(1'b1), .Q(cacheD
		[36]));
	notech_mux2 i_3530(.S(n_1573), .A(n_1562), .B(cacheD[36]), .Z(n_5640));
	notech_and4 i_1395(.A(n_60785), .B(n_62810), .C(cacheQ[90]), .D(n_60717)
		, .Z(n_1961));
	notech_reg_set cacheD_reg_37(.CP(n_63294), .D(n_5646), .SD(1'b1), .Q(cacheD
		[37]));
	notech_mux2 i_3538(.S(n_1573), .A(n_1559), .B(cacheD[37]), .Z(n_5646));
	notech_nao3 i_2722041(.A(n_2323), .B(n_2322), .C(n_1961), .Z(read_data[
		26]));
	notech_reg_set cacheD_reg_38(.CP(n_63294), .D(n_5652), .SD(1'b1), .Q(cacheD
		[38]));
	notech_mux2 i_3546(.S(n_1573), .A(n_1556), .B(cacheD[38]), .Z(n_5652));
	notech_reg_set cacheD_reg_39(.CP(n_63294), .D(n_5658), .SD(1'b1), .Q(cacheD
		[39]));
	notech_mux2 i_3554(.S(n_1573), .A(n_1553), .B(cacheD[39]), .Z(n_5658));
	notech_reg_set cacheD_reg_40(.CP(n_63342), .D(n_5664), .SD(1'b1), .Q(cacheD
		[40]));
	notech_mux2 i_3562(.S(n_1573), .A(n_1550), .B(cacheD[40]), .Z(n_5664));
	notech_reg_set cacheD_reg_41(.CP(n_63312), .D(n_5670), .SD(1'b1), .Q(cacheD
		[41]));
	notech_mux2 i_3570(.S(n_1573), .A(n_1547), .B(cacheD[41]), .Z(n_5670));
	notech_reg_set cacheD_reg_42(.CP(n_63312), .D(n_5676), .SD(1'b1), .Q(cacheD
		[42]));
	notech_mux2 i_3578(.S(n_1573), .A(n_1544), .B(cacheD[42]), .Z(n_5676));
	notech_and4 i_1404(.A(n_60785), .B(n_62810), .C(cacheQ[91]), .D(n_60717)
		, .Z(n_1967));
	notech_reg_set cacheD_reg_43(.CP(n_63312), .D(n_5682), .SD(1'b1), .Q(cacheD
		[43]));
	notech_mux2 i_3586(.S(n_1573), .A(n_1541), .B(cacheD[43]), .Z(n_5682));
	notech_nao3 i_2822042(.A(n_2326), .B(n_2325), .C(n_1967), .Z(read_data[
		27]));
	notech_reg_set cacheD_reg_44(.CP(n_63312), .D(n_5688), .SD(1'b1), .Q(cacheD
		[44]));
	notech_mux2 i_3594(.S(n_1573), .A(n_1538), .B(cacheD[44]), .Z(n_5688));
	notech_reg_set cacheD_reg_45(.CP(n_63312), .D(n_5694), .SD(1'b1), .Q(cacheD
		[45]));
	notech_mux2 i_3602(.S(n_1573), .A(n_1535), .B(cacheD[45]), .Z(n_5694));
	notech_reg_set cacheD_reg_46(.CP(n_63312), .D(n_5700), .SD(1'b1), .Q(cacheD
		[46]));
	notech_mux2 i_3610(.S(n_1573), .A(n_1532), .B(cacheD[46]), .Z(n_5700));
	notech_reg_set cacheD_reg_47(.CP(n_63312), .D(n_5706), .SD(1'b1), .Q(cacheD
		[47]));
	notech_mux2 i_3618(.S(n_1573), .A(n_1529), .B(cacheD[47]), .Z(n_5706));
	notech_reg_set cacheD_reg_48(.CP(n_63312), .D(n_5712), .SD(1'b1), .Q(cacheD
		[48]));
	notech_mux2 i_3626(.S(n_60671), .A(n_1526), .B(cacheD[48]), .Z(n_5712)
		);
	notech_and4 i_1413(.A(n_60785), .B(n_62810), .C(cacheQ[92]), .D(n_60717)
		, .Z(n_1973));
	notech_reg_set cacheD_reg_49(.CP(n_63312), .D(n_5718), .SD(1'b1), .Q(cacheD
		[49]));
	notech_mux2 i_3634(.S(n_60671), .A(n_1523), .B(cacheD[49]), .Z(n_5718)
		);
	notech_nao3 i_2922043(.A(n_2329), .B(n_2328), .C(n_1973), .Z(read_data[
		28]));
	notech_reg_set cacheD_reg_50(.CP(n_63312), .D(n_5724), .SD(1'b1), .Q(cacheD
		[50]));
	notech_mux2 i_3642(.S(n_60671), .A(n_1520), .B(cacheD[50]), .Z(n_5724)
		);
	notech_reg_set cacheD_reg_51(.CP(n_63312), .D(n_5730), .SD(1'b1), .Q(cacheD
		[51]));
	notech_mux2 i_3650(.S(n_60671), .A(n_1517), .B(cacheD[51]), .Z(n_5730)
		);
	notech_reg_set cacheD_reg_52(.CP(n_63312), .D(n_5736), .SD(1'b1), .Q(cacheD
		[52]));
	notech_mux2 i_3658(.S(n_60671), .A(n_1514), .B(cacheD[52]), .Z(n_5736)
		);
	notech_reg_set cacheD_reg_53(.CP(n_63312), .D(n_5742), .SD(1'b1), .Q(cacheD
		[53]));
	notech_mux2 i_3666(.S(n_60671), .A(n_1511), .B(cacheD[53]), .Z(n_5742)
		);
	notech_reg_set cacheD_reg_54(.CP(n_63312), .D(n_5748), .SD(1'b1), .Q(cacheD
		[54]));
	notech_mux2 i_3674(.S(n_60671), .A(n_1508), .B(cacheD[54]), .Z(n_5748)
		);
	notech_and4 i_1422(.A(n_60785), .B(n_62810), .C(cacheQ[93]), .D(n_60720)
		, .Z(n_1979));
	notech_reg_set cacheD_reg_55(.CP(n_63312), .D(n_5754), .SD(1'b1), .Q(cacheD
		[55]));
	notech_mux2 i_3682(.S(n_60671), .A(n_1505), .B(cacheD[55]), .Z(n_5754)
		);
	notech_nao3 i_3022044(.A(n_2332), .B(n_2331), .C(n_1979), .Z(read_data[
		29]));
	notech_reg_set cacheD_reg_56(.CP(n_63312), .D(n_5760), .SD(1'b1), .Q(cacheD
		[56]));
	notech_mux2 i_3690(.S(n_60671), .A(n_1502), .B(cacheD[56]), .Z(n_5760)
		);
	notech_reg_set cacheD_reg_57(.CP(n_63312), .D(n_5766), .SD(1'b1), .Q(cacheD
		[57]));
	notech_mux2 i_3698(.S(n_60671), .A(n_1499), .B(cacheD[57]), .Z(n_5766)
		);
	notech_reg_set cacheD_reg_58(.CP(n_63312), .D(n_5772), .SD(1'b1), .Q(cacheD
		[58]));
	notech_mux2 i_3706(.S(n_60671), .A(n_1496), .B(cacheD[58]), .Z(n_5772)
		);
	notech_reg_set cacheD_reg_59(.CP(n_63312), .D(n_5778), .SD(1'b1), .Q(cacheD
		[59]));
	notech_mux2 i_3714(.S(n_60671), .A(n_1493), .B(cacheD[59]), .Z(n_5778)
		);
	notech_reg_set cacheD_reg_60(.CP(n_63350), .D(n_5784), .SD(1'b1), .Q(cacheD
		[60]));
	notech_mux2 i_3722(.S(n_60671), .A(n_1490), .B(cacheD[60]), .Z(n_5784)
		);
	notech_and4 i_1431(.A(n_60789), .B(n_62810), .C(cacheQ[94]), .D(n_60720)
		, .Z(n_1985));
	notech_reg_set cacheD_reg_61(.CP(n_63334), .D(n_5790), .SD(1'b1), .Q(cacheD
		[61]));
	notech_mux2 i_3730(.S(n_60671), .A(n_1487), .B(cacheD[61]), .Z(n_5790)
		);
	notech_nao3 i_3122045(.A(n_2335), .B(n_2334), .C(n_1985), .Z(read_data[
		30]));
	notech_reg_set cacheD_reg_62(.CP(n_63350), .D(n_5796), .SD(1'b1), .Q(cacheD
		[62]));
	notech_mux2 i_3738(.S(n_60671), .A(n_1484), .B(cacheD[62]), .Z(n_5796)
		);
	notech_reg_set cacheD_reg_63(.CP(n_63350), .D(n_5802), .SD(1'b1), .Q(cacheD
		[63]));
	notech_mux2 i_3746(.S(n_60671), .A(n_1481), .B(cacheD[63]), .Z(n_5802)
		);
	notech_reg_set cacheD_reg_64(.CP(n_63350), .D(n_5808), .SD(1'b1), .Q(cacheD
		[64]));
	notech_mux2 i_3754(.S(n_1474), .A(n_1478), .B(cacheD[64]), .Z(n_5808));
	notech_reg_set cacheD_reg_65(.CP(n_63350), .D(n_5814), .SD(1'b1), .Q(cacheD
		[65]));
	notech_mux2 i_3762(.S(n_1474), .A(n_1472), .B(cacheD[65]), .Z(n_5814));
	notech_reg_set cacheD_reg_66(.CP(n_63350), .D(n_5820), .SD(1'b1), .Q(cacheD
		[66]));
	notech_mux2 i_3770(.S(n_1474), .A(n_1469), .B(cacheD[66]), .Z(n_5820));
	notech_and4 i_1440(.A(n_60789), .B(n_62810), .C(cacheQ[95]), .D(n_60720)
		, .Z(n_1991));
	notech_reg_set cacheD_reg_67(.CP(n_63350), .D(n_5826), .SD(1'b1), .Q(cacheD
		[67]));
	notech_mux2 i_3778(.S(n_1474), .A(n_1466), .B(cacheD[67]), .Z(n_5826));
	notech_nao3 i_3222046(.A(n_2338), .B(n_2337), .C(n_1991), .Z(read_data[
		31]));
	notech_reg_set cacheD_reg_68(.CP(n_63350), .D(n_5832), .SD(1'b1), .Q(cacheD
		[68]));
	notech_mux2 i_3786(.S(n_1474), .A(n_1463), .B(cacheD[68]), .Z(n_5832));
	notech_reg_set cacheD_reg_69(.CP(n_63350), .D(n_5838), .SD(1'b1), .Q(cacheD
		[69]));
	notech_mux2 i_3794(.S(n_1474), .A(n_1460), .B(cacheD[69]), .Z(n_5838));
	notech_nand2 i_49(.A(n_8325), .B(fsm[3]), .Z(n_1994));
	notech_reg_set cacheD_reg_70(.CP(n_63350), .D(n_5844), .SD(1'b1), .Q(cacheD
		[70]));
	notech_mux2 i_3802(.S(n_1474), .A(n_1457), .B(cacheD[70]), .Z(n_5844));
	notech_nao3 i_117(.A(fsm[1]), .B(fsm[3]), .C(fsm[0]), .Z(n_1995));
	notech_reg_set cacheD_reg_71(.CP(n_63350), .D(n_5850), .SD(1'b1), .Q(cacheD
		[71]));
	notech_mux2 i_3810(.S(n_1474), .A(n_1454), .B(cacheD[71]), .Z(n_5850));
	notech_nao3 i_1329988(.A(fsm[4]), .B(fsm[2]), .C(n_1995), .Z(n_1996));
	notech_reg_set cacheD_reg_72(.CP(n_63350), .D(n_5856), .SD(1'b1), .Q(cacheD
		[72]));
	notech_mux2 i_3818(.S(n_1474), .A(n_1451), .B(cacheD[72]), .Z(n_5856));
	notech_reg_set cacheD_reg_73(.CP(n_63350), .D(n_5862), .SD(1'b1), .Q(cacheD
		[73]));
	notech_mux2 i_3826(.S(n_1474), .A(n_1448), .B(cacheD[73]), .Z(n_5862));
	notech_nand3 i_68(.A(fsm[1]), .B(fsm[3]), .C(fsm[0]), .Z(n_1998));
	notech_reg_set cacheD_reg_74(.CP(n_63350), .D(n_5868), .SD(1'b1), .Q(cacheD
		[74]));
	notech_mux2 i_3834(.S(n_1474), .A(n_1445), .B(cacheD[74]), .Z(n_5868));
	notech_and2 i_48(.A(n_8327), .B(n_8326), .Z(n_1999));
	notech_reg_set cacheD_reg_75(.CP(n_63350), .D(n_5874), .SD(1'b1), .Q(cacheD
		[75]));
	notech_mux2 i_3842(.S(n_1474), .A(n_1442), .B(cacheD[75]), .Z(n_5874));
	notech_nao3 i_31(.A(n_8327), .B(n_8326), .C(fsm[4]), .Z(n_2000));
	notech_reg_set cacheD_reg_76(.CP(n_63350), .D(n_5880), .SD(1'b1), .Q(cacheD
		[76]));
	notech_mux2 i_3850(.S(n_1474), .A(n_1439), .B(cacheD[76]), .Z(n_5880));
	notech_reg_set cacheD_reg_77(.CP(n_63350), .D(n_5886), .SD(1'b1), .Q(cacheD
		[77]));
	notech_mux2 i_3858(.S(n_1474), .A(n_1436), .B(cacheD[77]), .Z(n_5886));
	notech_or4 i_113(.A(fsm[0]), .B(fsm[3]), .C(n_2000), .D(n_970), .Z(n_2002
		));
	notech_reg_set cacheD_reg_78(.CP(n_63350), .D(n_5892), .SD(1'b1), .Q(cacheD
		[78]));
	notech_mux2 i_3866(.S(n_1474), .A(n_1433), .B(cacheD[78]), .Z(n_5892));
	notech_and2 i_56024(.A(write_req), .B(n_8563), .Z(n_2003));
	notech_reg_set cacheD_reg_79(.CP(n_63350), .D(n_5898), .SD(1'b1), .Q(cacheD
		[79]));
	notech_mux2 i_3874(.S(n_1474), .A(n_1430), .B(cacheD[79]), .Z(n_5898));
	notech_ao3 i_14(.A(n_62810), .B(n_8323), .C(n_1742), .Z(n_2004));
	notech_reg_set cacheD_reg_80(.CP(n_63348), .D(n_5904), .SD(1'b1), .Q(cacheD
		[80]));
	notech_mux2 i_3882(.S(n_60693), .A(n_1427), .B(cacheD[80]), .Z(n_5904)
		);
	notech_reg_set cacheD_reg_81(.CP(n_63356), .D(n_5910), .SD(1'b1), .Q(cacheD
		[81]));
	notech_mux2 i_3890(.S(n_60693), .A(n_1424), .B(cacheD[81]), .Z(n_5910)
		);
	notech_reg_set cacheD_reg_82(.CP(n_63356), .D(n_5916), .SD(1'b1), .Q(cacheD
		[82]));
	notech_mux2 i_3898(.S(n_60693), .A(n_1421), .B(cacheD[82]), .Z(n_5916)
		);
	notech_or4 i_140(.A(code_wack), .B(n_971), .C(n_2003), .D(n_8566), .Z(n_2007
		));
	notech_reg_set cacheD_reg_83(.CP(n_63356), .D(n_5922), .SD(1'b1), .Q(cacheD
		[83]));
	notech_mux2 i_3906(.S(n_60693), .A(n_1418), .B(cacheD[83]), .Z(n_5922)
		);
	notech_or2 i_56135(.A(n_2002), .B(n_2007), .Z(n_2008));
	notech_reg_set cacheD_reg_84(.CP(n_63356), .D(n_5928), .SD(1'b1), .Q(cacheD
		[84]));
	notech_mux2 i_3914(.S(n_60693), .A(n_1415), .B(cacheD[84]), .Z(n_5928)
		);
	notech_reg_set cacheD_reg_85(.CP(n_63356), .D(n_5934), .SD(1'b1), .Q(cacheD
		[85]));
	notech_mux2 i_3922(.S(n_60693), .A(n_1412), .B(cacheD[85]), .Z(n_5934)
		);
	notech_or4 i_56122(.A(code_ack), .B(n_2003), .C(n_2002), .D(n_8564), .Z(n_2010
		));
	notech_reg_set cacheD_reg_86(.CP(n_63356), .D(n_5940), .SD(1'b1), .Q(cacheD
		[86]));
	notech_mux2 i_3930(.S(n_60693), .A(n_1409), .B(cacheD[86]), .Z(n_5940)
		);
	notech_reg_set cacheD_reg_87(.CP(n_63356), .D(n_5946), .SD(1'b1), .Q(cacheD
		[87]));
	notech_mux2 i_3938(.S(n_60693), .A(n_1406), .B(cacheD[87]), .Z(n_5946)
		);
	notech_reg_set cacheD_reg_88(.CP(n_63356), .D(n_5952), .SD(1'b1), .Q(cacheD
		[88]));
	notech_mux2 i_3946(.S(n_60693), .A(n_1403), .B(cacheD[88]), .Z(n_5952)
		);
	notech_reg_set cacheD_reg_89(.CP(n_63356), .D(n_5958), .SD(1'b1), .Q(cacheD
		[89]));
	notech_mux2 i_3954(.S(n_60693), .A(n_1400), .B(cacheD[89]), .Z(n_5958)
		);
	notech_reg_set cacheD_reg_90(.CP(n_63356), .D(n_5964), .SD(1'b1), .Q(cacheD
		[90]));
	notech_mux2 i_3962(.S(n_60693), .A(n_1397), .B(cacheD[90]), .Z(n_5964)
		);
	notech_reg_set cacheD_reg_91(.CP(n_63356), .D(n_5970), .SD(1'b1), .Q(cacheD
		[91]));
	notech_mux2 i_3970(.S(n_60693), .A(n_1394), .B(cacheD[91]), .Z(n_5970)
		);
	notech_and2 i_27(.A(axi_RVALID), .B(axi_RLAST), .Z(n_2016));
	notech_reg_set cacheD_reg_92(.CP(n_63356), .D(n_5976), .SD(1'b1), .Q(cacheD
		[92]));
	notech_mux2 i_3978(.S(n_60693), .A(n_1391), .B(cacheD[92]), .Z(n_5976)
		);
	notech_or2 i_116(.A(fsm[4]), .B(fsm[2]), .Z(n_2017));
	notech_reg_set cacheD_reg_93(.CP(n_63356), .D(n_5982), .SD(1'b1), .Q(cacheD
		[93]));
	notech_mux2 i_3986(.S(n_60693), .A(n_1388), .B(cacheD[93]), .Z(n_5982)
		);
	notech_reg_set cacheD_reg_94(.CP(n_63356), .D(n_5988), .SD(1'b1), .Q(cacheD
		[94]));
	notech_mux2 i_3994(.S(n_60693), .A(n_1385), .B(cacheD[94]), .Z(n_5988)
		);
	notech_or4 i_56097(.A(n_2017), .B(n_2003), .C(n_1998), .D(n_8217), .Z(n_2019
		));
	notech_reg_set cacheD_reg_95(.CP(n_63356), .D(n_5994), .SD(1'b1), .Q(cacheD
		[95]));
	notech_mux2 i_4002(.S(n_60693), .A(n_1382), .B(cacheD[95]), .Z(n_5994)
		);
	notech_ao3 i_52(.A(n_62810), .B(n_2019), .C(n_1742), .Z(n_2020));
	notech_reg_set cacheD_reg_96(.CP(n_63356), .D(n_6000), .SD(1'b1), .Q(cacheD
		[96]));
	notech_mux2 i_4010(.S(n_1375), .A(n_1379), .B(cacheD[96]), .Z(n_6000));
	notech_and2 i_12(.A(axi_AR[30]), .B(n_8559), .Z(n_2021));
	notech_reg_set cacheD_reg_97(.CP(n_63356), .D(n_6006), .SD(1'b1), .Q(cacheD
		[97]));
	notech_mux2 i_4018(.S(n_1375), .A(n_1373), .B(cacheD[97]), .Z(n_6006));
	notech_and2 i_110(.A(n_1066), .B(n_62793), .Z(n_2022));
	notech_reg_set cacheD_reg_98(.CP(n_63356), .D(n_6012), .SD(1'b1), .Q(cacheD
		[98]));
	notech_mux2 i_4026(.S(n_1375), .A(n_1370), .B(cacheD[98]), .Z(n_6012));
	notech_ao3 i_56102(.A(n_8325), .B(fsm[3]), .C(n_2000), .Z(n_2023));
	notech_reg_set cacheD_reg_99(.CP(n_63356), .D(n_6018), .SD(1'b1), .Q(cacheD
		[99]));
	notech_mux2 i_4034(.S(n_1375), .A(n_1367), .B(cacheD[99]), .Z(n_6018));
	notech_and2 i_33(.A(n_8265), .B(n_62123), .Z(n_2024));
	notech_reg_set cacheD_reg_100(.CP(n_63356), .D(n_6024), .SD(1'b1), .Q(cacheD
		[100]));
	notech_mux2 i_4042(.S(n_1375), .A(n_1364), .B(cacheD[100]), .Z(n_6024)
		);
	notech_nand2 i_13(.A(burst_idx[0]), .B(burst_idx[1]), .Z(n_2025));
	notech_reg_set cacheD_reg_101(.CP(n_63332), .D(n_6030), .SD(1'b1), .Q(cacheD
		[101]));
	notech_mux2 i_4050(.S(n_1375), .A(n_1361), .B(cacheD[101]), .Z(n_6030)
		);
	notech_nand3 i_42(.A(burst_idx[0]), .B(burst_idx[1]), .C(burst_idx[2]), 
		.Z(n_2026));
	notech_reg_set cacheD_reg_102(.CP(n_63332), .D(n_6036), .SD(1'b1), .Q(cacheD
		[102]));
	notech_mux2 i_4058(.S(n_1375), .A(n_1358), .B(cacheD[102]), .Z(n_6036)
		);
	notech_nao3 i_72(.A(burst_idx[2]), .B(burst_idx[3]), .C(n_2025), .Z(n_2027
		));
	notech_reg_set cacheD_reg_103(.CP(n_63332), .D(n_6042), .SD(1'b1), .Q(cacheD
		[103]));
	notech_mux2 i_4066(.S(n_1375), .A(n_1355), .B(cacheD[103]), .Z(n_6042)
		);
	notech_nor2 i_120(.A(burst_idx[0]), .B(n_8302), .Z(n_2028));
	notech_reg_set cacheD_reg_104(.CP(n_63332), .D(n_6048), .SD(1'b1), .Q(cacheD
		[104]));
	notech_mux2 i_4074(.S(n_1375), .A(n_1352), .B(cacheD[104]), .Z(n_6048)
		);
	notech_and2 i_124(.A(burst_idx[0]), .B(n_8302), .Z(n_2029));
	notech_reg_set cacheD_reg_105(.CP(n_63332), .D(n_6054), .SD(1'b1), .Q(cacheD
		[105]));
	notech_mux2 i_4082(.S(n_1375), .A(n_1349), .B(cacheD[105]), .Z(n_6054)
		);
	notech_nand2 i_53(.A(axi_RVALID), .B(n_62728), .Z(n_2030));
	notech_reg_set cacheD_reg_106(.CP(n_63332), .D(n_6060), .SD(1'b1), .Q(cacheD
		[106]));
	notech_mux2 i_4090(.S(n_1375), .A(n_1346), .B(cacheD[106]), .Z(n_6060)
		);
	notech_reg_set cacheD_reg_107(.CP(n_63332), .D(n_6066), .SD(1'b1), .Q(cacheD
		[107]));
	notech_mux2 i_4098(.S(n_1375), .A(n_1343), .B(cacheD[107]), .Z(n_6066)
		);
	notech_nand2 i_343(.A(n_8328), .B(fsm[0]), .Z(n_2032));
	notech_reg_set cacheD_reg_108(.CP(n_63332), .D(n_6072), .SD(1'b1), .Q(cacheD
		[108]));
	notech_mux2 i_4106(.S(n_1375), .A(n_1340), .B(cacheD[108]), .Z(n_6072)
		);
	notech_ao3 i_1129979(.A(n_8328), .B(fsm[0]), .C(n_2000), .Z(n_2033));
	notech_reg_set cacheD_reg_109(.CP(n_63332), .D(n_6078), .SD(1'b1), .Q(cacheD
		[109]));
	notech_mux2 i_4114(.S(n_1375), .A(n_1337), .B(cacheD[109]), .Z(n_6078)
		);
	notech_reg_set cacheD_reg_110(.CP(n_63332), .D(n_6084), .SD(1'b1), .Q(cacheD
		[110]));
	notech_mux2 i_4122(.S(n_1375), .A(n_1334), .B(cacheD[110]), .Z(n_6084)
		);
	notech_ao3 i_56(.A(n_8303), .B(n_8304), .C(burst_idx[4]), .Z(n_2035));
	notech_reg_set cacheD_reg_111(.CP(n_63332), .D(n_6090), .SD(1'b1), .Q(cacheD
		[111]));
	notech_mux2 i_4130(.S(n_1375), .A(n_1331), .B(cacheD[111]), .Z(n_6090)
		);
	notech_or2 i_114(.A(burst_idx[0]), .B(burst_idx[1]), .Z(n_2036));
	notech_reg_set cacheD_reg_112(.CP(n_63332), .D(n_6096), .SD(1'b1), .Q(cacheD
		[112]));
	notech_mux2 i_4138(.S(n_60798), .A(n_1328), .B(cacheD[112]), .Z(n_6096)
		);
	notech_ao3 i_5780763(.A(n_910), .B(n_909), .C(n_894), .Z(n_2037));
	notech_reg_set cacheD_reg_113(.CP(n_63332), .D(n_6102), .SD(1'b1), .Q(cacheD
		[113]));
	notech_mux2 i_4146(.S(n_60798), .A(n_1325), .B(cacheD[113]), .Z(n_6102)
		);
	notech_reg_set cacheD_reg_114(.CP(n_63332), .D(n_6108), .SD(1'b1), .Q(cacheD
		[114]));
	notech_mux2 i_4154(.S(n_60798), .A(n_1322), .B(cacheD[114]), .Z(n_6108)
		);
	notech_reg_set cacheD_reg_115(.CP(n_63332), .D(n_6114), .SD(1'b1), .Q(cacheD
		[115]));
	notech_mux2 i_4162(.S(n_60798), .A(n_1319), .B(cacheD[115]), .Z(n_6114)
		);
	notech_or4 i_347(.A(axi_AWVALID), .B(n_2036), .C(n_8220), .D(n_8557), .Z
		(n_2040));
	notech_reg_set cacheD_reg_116(.CP(n_63332), .D(n_6120), .SD(1'b1), .Q(cacheD
		[116]));
	notech_mux2 i_4170(.S(n_60798), .A(n_1316), .B(cacheD[116]), .Z(n_6120)
		);
	notech_or4 i_21(.A(burst_idx[2]), .B(burst_idx[3]), .C(burst_idx[4]), .D
		(n_2040), .Z(n_2041));
	notech_reg_set cacheD_reg_117(.CP(n_63332), .D(n_6126), .SD(1'b1), .Q(cacheD
		[117]));
	notech_mux2 i_4178(.S(n_60798), .A(n_1313), .B(cacheD[117]), .Z(n_6126)
		);
	notech_nor2 i_15(.A(n_25047), .B(n_62170), .Z(n_2042));
	notech_reg_set cacheD_reg_118(.CP(n_63332), .D(n_6132), .SD(1'b1), .Q(cacheD
		[118]));
	notech_mux2 i_4186(.S(n_60798), .A(n_1310), .B(cacheD[118]), .Z(n_6132)
		);
	notech_reg_set cacheD_reg_119(.CP(n_63332), .D(n_6138), .SD(1'b1), .Q(cacheD
		[119]));
	notech_mux2 i_4194(.S(n_60798), .A(n_1307), .B(cacheD[119]), .Z(n_6138)
		);
	notech_reg_set cacheD_reg_120(.CP(n_63352), .D(n_6144), .SD(1'b1), .Q(cacheD
		[120]));
	notech_mux2 i_4202(.S(n_60798), .A(n_1304), .B(cacheD[120]), .Z(n_6144)
		);
	notech_or4 i_56114(.A(fsm[4]), .B(fsm[1]), .C(n_1994), .D(n_8327), .Z(n_2045
		));
	notech_reg_set cacheD_reg_121(.CP(n_63314), .D(n_6150), .SD(1'b1), .Q(cacheD
		[121]));
	notech_mux2 i_4210(.S(n_60798), .A(n_1301), .B(cacheD[121]), .Z(n_6150)
		);
	notech_ao4 i_385(.A(code_req), .B(n_8265), .C(n_2045), .D(read_req), .Z(n_2046
		));
	notech_reg_set cacheD_reg_122(.CP(n_63314), .D(n_6156), .SD(1'b1), .Q(cacheD
		[122]));
	notech_mux2 i_4218(.S(n_60798), .A(n_1298), .B(cacheD[122]), .Z(n_6156)
		);
	notech_reg_set cacheD_reg_123(.CP(n_63314), .D(n_6162), .SD(1'b1), .Q(cacheD
		[123]));
	notech_mux2 i_4226(.S(n_60798), .A(n_1295), .B(cacheD[123]), .Z(n_6162)
		);
	notech_reg_set cacheD_reg_124(.CP(n_63314), .D(n_6168), .SD(1'b1), .Q(cacheD
		[124]));
	notech_mux2 i_4234(.S(n_60798), .A(n_1292), .B(cacheD[124]), .Z(n_6168)
		);
	notech_or4 i_47(.A(n_928), .B(n_944), .C(n_943), .D(n_8557), .Z(n_2049)
		);
	notech_reg_set cacheD_reg_125(.CP(n_63314), .D(n_6174), .SD(1'b1), .Q(cacheD
		[125]));
	notech_mux2 i_4242(.S(n_60798), .A(n_1289), .B(cacheD[125]), .Z(n_6174)
		);
	notech_nor2 i_125(.A(n_2019), .B(n_2021), .Z(n_2050));
	notech_reg_set cacheD_reg_126(.CP(n_63314), .D(n_6180), .SD(1'b1), .Q(cacheD
		[126]));
	notech_mux2 i_4250(.S(n_60798), .A(n_1286), .B(cacheD[126]), .Z(n_6180)
		);
	notech_ao4 i_46(.A(n_2049), .B(n_8216), .C(n_1995), .D(n_2017), .Z(n_2051
		));
	notech_reg_set cacheD_reg_127(.CP(n_63314), .D(n_6186), .SD(1'b1), .Q(cacheD
		[127]));
	notech_mux2 i_4258(.S(n_60798), .A(n_1283), .B(cacheD[127]), .Z(n_6186)
		);
	notech_and2 i_30(.A(axi_RREADY), .B(axi_RVALID), .Z(n_2052));
	notech_reg_set cacheD_reg_128(.CP(n_63314), .D(n_6192), .SD(1'b1), .Q(cacheD
		[128]));
	notech_mux2 i_4266(.S(n_1277), .A(n_8324), .B(cacheD[128]), .Z(n_6192)
		);
	notech_reg_set cacheD_reg_129(.CP(n_63314), .D(n_6198), .SD(1'b1), .Q(cacheD
		[129]));
	notech_mux2 i_4274(.S(n_1277), .A(n_8322), .B(cacheD[129]), .Z(n_6198)
		);
	notech_reg_set cacheD_reg_130(.CP(n_63314), .D(n_6204), .SD(1'b1), .Q(cacheD
		[130]));
	notech_mux2 i_4282(.S(n_1277), .A(n_8321), .B(cacheD[130]), .Z(n_6204)
		);
	notech_reg_set cacheD_reg_131(.CP(n_63314), .D(n_6210), .SD(1'b1), .Q(cacheD
		[131]));
	notech_mux2 i_4290(.S(n_1277), .A(n_8320), .B(cacheD[131]), .Z(n_6210)
		);
	notech_and2 i_57(.A(n_2045), .B(n_2042), .Z(n_2056));
	notech_reg_set cacheD_reg_132(.CP(n_63314), .D(n_6216), .SD(1'b1), .Q(cacheD
		[132]));
	notech_mux2 i_4298(.S(n_1277), .A(n_8319), .B(cacheD[132]), .Z(n_6216)
		);
	notech_and3 i_73(.A(n_2045), .B(n_2051), .C(n_2042), .Z(n_2057));
	notech_reg_set cacheD_reg_133(.CP(n_63314), .D(n_6222), .SD(1'b1), .Q(cacheD
		[133]));
	notech_mux2 i_4306(.S(n_1277), .A(n_8318), .B(cacheD[133]), .Z(n_6222)
		);
	notech_and2 i_119(.A(n_2057), .B(n_8265), .Z(n_2058));
	notech_reg_set cacheD_reg_134(.CP(n_63314), .D(n_6228), .SD(1'b1), .Q(cacheD
		[134]));
	notech_mux2 i_4314(.S(n_1277), .A(n_8317), .B(cacheD[134]), .Z(n_6228)
		);
	notech_reg_set cacheD_reg_135(.CP(n_63314), .D(n_6234), .SD(1'b1), .Q(cacheD
		[135]));
	notech_mux2 i_4322(.S(n_1277), .A(n_8316), .B(cacheD[135]), .Z(n_6234)
		);
	notech_reg_set cacheD_reg_136(.CP(n_63314), .D(n_6240), .SD(1'b1), .Q(cacheD
		[136]));
	notech_mux2 i_4330(.S(n_1277), .A(n_8315), .B(cacheD[136]), .Z(n_6240)
		);
	notech_and4 i_402(.A(n_2019), .B(n_1205), .C(n_1215), .D(n_8300), .Z(n_2061
		));
	notech_reg_set cacheD_reg_137(.CP(n_63314), .D(n_6246), .SD(1'b1), .Q(cacheD
		[137]));
	notech_mux2 i_4338(.S(n_1277), .A(n_8314), .B(cacheD[137]), .Z(n_6246)
		);
	notech_reg_set cacheD_reg_138(.CP(n_63352), .D(n_6252), .SD(1'b1), .Q(cacheD
		[138]));
	notech_mux2 i_4346(.S(n_1277), .A(n_8313), .B(cacheD[138]), .Z(n_6252)
		);
	notech_reg_set cacheD_reg_139(.CP(n_63336), .D(n_6258), .SD(1'b1), .Q(cacheD
		[139]));
	notech_mux2 i_4354(.S(n_60809), .A(n_8312), .B(cacheD[139]), .Z(n_6258)
		);
	notech_ao4 i_71(.A(n_2045), .B(n_8213), .C(n_2024), .D(n_8214), .Z(n_2064
		));
	notech_reg_set cacheD_reg_140(.CP(n_63352), .D(n_6264), .SD(1'b1), .Q(cacheD
		[140]));
	notech_mux2 i_4362(.S(n_60809), .A(n_8311), .B(cacheD[140]), .Z(n_6264)
		);
	notech_reg_set cacheD_reg_141(.CP(n_63352), .D(n_6270), .SD(1'b1), .Q(cacheD
		[141]));
	notech_mux2 i_4370(.S(n_60809), .A(n_8310), .B(cacheD[141]), .Z(n_6270)
		);
	notech_and4 i_415(.A(n_2019), .B(n_1205), .C(n_973), .D(n_8300), .Z(n_2066
		));
	notech_reg_set cacheD_reg_142(.CP(n_63352), .D(n_6276), .SD(1'b1), .Q(cacheD
		[142]));
	notech_mux2 i_4378(.S(n_60809), .A(n_8309), .B(cacheD[142]), .Z(n_6276)
		);
	notech_reg_set cacheD_reg_143(.CP(n_63352), .D(n_6282), .SD(1'b1), .Q(cacheD
		[143]));
	notech_mux2 i_4386(.S(n_60809), .A(n_8308), .B(cacheD[143]), .Z(n_6282)
		);
	notech_reg_set cacheD_reg_144(.CP(n_63352), .D(n_6288), .SD(1'b1), .Q(cacheD
		[144]));
	notech_mux2 i_4394(.S(n_60809), .A(n_8306), .B(cacheD[144]), .Z(n_6288)
		);
	notech_and2 i_0(.A(n_62170), .B(n_8562), .Z(n_2069));
	notech_reg_set cacheD_reg_145(.CP(n_63352), .D(n_6294), .SD(1'b1), .Q(cacheD
		[145]));
	notech_mux2 i_4402(.S(n_60809), .A(n_8305), .B(cacheD[145]), .Z(n_6294)
		);
	notech_and2 i_51(.A(n_62820), .B(n_1167), .Z(n_2070));
	notech_reg_set cacheD_reg_146(.CP(n_63352), .D(n_6300), .SD(1'b1), .Q(cacheD
		[146]));
	notech_mux2 i_4410(.S(n_1277), .A(n_23512), .B(cacheD[146]), .Z(n_6300)
		);
	notech_nand3 i_474(.A(axi_RVALID), .B(axi_RLAST), .C(n_62728), .Z(n_2071
		));
	notech_reg_set cacheD_reg_147(.CP(n_63352), .D(n_6306), .SD(1'b1), .Q(cacheD
		[147]));
	notech_mux2 i_4418(.S(n_60809), .A(n_23517), .B(cacheD[147]), .Z(n_6306)
		);
	notech_ao3 i_67(.A(n_62170), .B(n_60789), .C(n_21466), .Z(n_2072));
	notech_reg_set cacheD_reg_148(.CP(n_63352), .D(n_6312), .SD(1'b1), .Q(cacheD
		[148]));
	notech_mux2 i_4426(.S(n_60809), .A(n_1224), .B(cacheD[148]), .Z(n_6312)
		);
	notech_nand3 i_37(.A(n_60789), .B(n_2069), .C(n_60717), .Z(n_2073));
	notech_reg_set cacheD_reg_149(.CP(n_63352), .D(n_6318), .SD(1'b1), .Q(cacheD
		[149]));
	notech_mux2 i_4434(.S(n_60809), .A(n_23527), .B(cacheD[149]), .Z(n_6318)
		);
	notech_or4 i_65(.A(n_21466), .B(n_60789), .C(n_2032), .D(n_2000), .Z(n_2074
		));
	notech_reg axi_WSTRB_reg_0(.CP(n_63352), .D(n_6324), .CD(n_62727), .Q(axi_WSTRB
		[0]));
	notech_mux2 i_4442(.S(n_62777), .A(n_8332), .B(axi_WSTRB[0]), .Z(n_6324)
		);
	notech_nand3 i_35(.A(n_60789), .B(n_2069), .C(n_60755), .Z(n_2075));
	notech_reg axi_WSTRB_reg_1(.CP(n_63352), .D(n_6330), .CD(n_62727), .Q(axi_WSTRB
		[1]));
	notech_mux2 i_4450(.S(n_62777), .A(n_25326), .B(axi_WSTRB[1]), .Z(n_6330
		));
	notech_reg axi_WSTRB_reg_2(.CP(n_63352), .D(n_6336), .CD(n_62727), .Q(axi_WSTRB
		[2]));
	notech_mux2 i_4458(.S(n_62777), .A(n_25332), .B(axi_WSTRB[2]), .Z(n_6336
		));
	notech_reg axi_WSTRB_reg_3(.CP(n_63352), .D(n_6342), .CD(n_62727), .Q(axi_WSTRB
		[3]));
	notech_mux2 i_4466(.S(n_62777), .A(n_25338), .B(axi_WSTRB[3]), .Z(n_6342
		));
	notech_reg_set cacheM_reg_0(.CP(n_63352), .D(n_6348), .SD(n_62728), .Q(cacheM
		[0]));
	notech_mux2 i_4474(.S(n_1744), .A(n_1746), .B(cacheM[0]), .Z(n_6348));
	notech_reg_set cacheM_reg_1(.CP(n_63352), .D(n_6354), .SD(n_62728), .Q(cacheM
		[1]));
	notech_mux2 i_4482(.S(n_1744), .A(n_1741), .B(cacheM[1]), .Z(n_6354));
	notech_reg_set cacheM_reg_2(.CP(n_63352), .D(n_6360), .SD(n_62727), .Q(cacheM
		[2]));
	notech_mux2 i_4490(.S(n_1744), .A(n_1739), .B(cacheM[2]), .Z(n_6360));
	notech_reg_set cacheM_reg_3(.CP(n_63314), .D(n_6366), .SD(n_62728), .Q(cacheM
		[3]));
	notech_mux2 i_4498(.S(n_1744), .A(n_1737), .B(cacheM[3]), .Z(n_6366));
	notech_reg_set cacheM_reg_4(.CP(n_63314), .D(n_6372), .SD(n_62728), .Q(cacheM
		[4]));
	notech_mux2 i_4506(.S(n_1744), .A(n_1735), .B(cacheM[4]), .Z(n_6372));
	notech_reg_set cacheM_reg_5(.CP(n_63338), .D(n_6378), .SD(n_62729), .Q(cacheM
		[5]));
	notech_mux2 i_4514(.S(n_1744), .A(n_1733), .B(cacheM[5]), .Z(n_6378));
	notech_reg_set cacheM_reg_6(.CP(n_63338), .D(n_6384), .SD(n_62729), .Q(cacheM
		[6]));
	notech_mux2 i_4522(.S(n_1744), .A(n_1731), .B(cacheM[6]), .Z(n_6384));
	notech_reg_set cacheM_reg_7(.CP(n_63338), .D(n_6390), .SD(n_62729), .Q(cacheM
		[7]));
	notech_mux2 i_4530(.S(n_1744), .A(n_1729), .B(cacheM[7]), .Z(n_6390));
	notech_reg_set cacheM_reg_8(.CP(n_63338), .D(n_6396), .SD(n_62729), .Q(cacheM
		[8]));
	notech_mux2 i_4538(.S(n_1744), .A(n_1727), .B(cacheM[8]), .Z(n_6396));
	notech_reg_set cacheM_reg_9(.CP(n_63338), .D(n_6402), .SD(n_62729), .Q(cacheM
		[9]));
	notech_mux2 i_4546(.S(n_1744), .A(n_1725), .B(cacheM[9]), .Z(n_6402));
	notech_reg_set cacheM_reg_10(.CP(n_63338), .D(n_6408), .SD(n_62729), .Q(cacheM
		[10]));
	notech_mux2 i_4554(.S(n_1744), .A(n_1723), .B(cacheM[10]), .Z(n_6408));
	notech_reg_set cacheM_reg_11(.CP(n_63338), .D(n_6414), .SD(n_62729), .Q(cacheM
		[11]));
	notech_mux2 i_4562(.S(n_1744), .A(n_1721), .B(cacheM[11]), .Z(n_6414));
	notech_reg_set cacheM_reg_12(.CP(n_63338), .D(n_6420), .SD(n_62729), .Q(cacheM
		[12]));
	notech_mux2 i_4570(.S(n_1744), .A(n_1719), .B(cacheM[12]), .Z(n_6420));
	notech_reg_set cacheM_reg_13(.CP(n_63338), .D(n_6426), .SD(n_62729), .Q(cacheM
		[13]));
	notech_mux2 i_4578(.S(n_1744), .A(n_1717), .B(cacheM[13]), .Z(n_6426));
	notech_reg_set cacheM_reg_14(.CP(n_63338), .D(n_6432), .SD(n_62729), .Q(cacheM
		[14]));
	notech_mux2 i_4586(.S(n_1744), .A(n_1715), .B(cacheM[14]), .Z(n_6432));
	notech_reg_set cacheM_reg_15(.CP(n_63338), .D(n_6438), .SD(n_62728), .Q(cacheM
		[15]));
	notech_mux2 i_4594(.S(n_1744), .A(n_1713), .B(cacheM[15]), .Z(n_6438));
	notech_reg_set cacheWEN_reg(.CP(n_63338), .D(n_6444), .SD(n_62728), .Q(cacheWEN
		));
	notech_mux2 i_4602(.S(n_1749), .A(n_1751), .B(cacheWEN), .Z(n_6444));
	notech_reg axi_RREADY_reg(.CP(n_63338), .D(n_6450), .CD(n_62729), .Q(axi_RREADY
		));
	notech_mux2 i_4610(.S(n_1755), .A(n_1756), .B(axi_RREADY), .Z(n_6450));
	notech_reg axi_ARVALID_reg(.CP(n_63338), .D(n_6456), .CD(n_62729), .Q(axi_ARVALID
		));
	notech_mux2 i_4618(.S(n_1759), .A(n_1760), .B(axi_ARVALID), .Z(n_6456)
		);
	notech_reg axi_io_WVALID_reg(.CP(n_63338), .D(n_6462), .CD(n_62729), .Q(axi_io_WVALID
		));
	notech_mux2 i_4626(.S(n_1763), .A(n_23624), .B(axi_io_WVALID), .Z(n_6462
		));
	notech_reg wf_reg(.CP(n_63338), .D(writeio_req), .CD(n_62729), .Q(wf));
	notech_reg rf_reg(.CP(n_63338), .D(readio_req), .CD(n_62722), .Q(rf));
	notech_reg axi_io_ARVALID_reg(.CP(n_63338), .D(n_6472), .CD(n_62715), .Q
		(axi_io_ARVALID));
	notech_mux2 i_4642(.S(n_1765), .A(n_8330), .B(axi_io_ARVALID), .Z(n_6472
		));
	notech_reg axi_io_RREADY_reg(.CP(n_63316), .D(n_6478), .CD(n_62715), .Q(axi_io_RREADY
		));
	notech_mux2 i_4650(.S(n_1766), .A(n_23569), .B(axi_io_RREADY), .Z(n_6478
		));
	notech_reg readio_ack_reg(.CP(n_63338), .D(n_6486), .CD(n_62714), .Q(readio_ack
		));
	notech_ao3 i_4659(.A(n_222956487), .B(n_222856486), .C(readio_ack), .Z(n_6486
		));
	notech_reg writeio_ack_reg(.CP(n_63292), .D(n_6490), .CD(n_62714), .Q(writeio_ack
		));
	notech_xor2 i_4666(.A(n_8560), .B(n_1769), .Z(n_6490));
	notech_reg axi_io_AWVALID_reg(.CP(n_63292), .D(n_6496), .CD(n_62715), .Q
		(axi_io_AWVALID));
	notech_mux2 i_4674(.S(n_1770), .A(n_8333), .B(axi_io_AWVALID), .Z(n_6496
		));
	notech_reg axi_ARSIZE_reg_0(.CP(n_63292), .D(n_6505), .CD(n_62715), .Q(axi_ARSIZE
		[0]));
	notech_and2 i_4684(.A(n_62793), .B(axi_ARSIZE[0]), .Z(n_6505));
	notech_reg_set axi_ARSIZE_reg_1(.CP(n_63292), .D(n_6513), .SD(n_62715), 
		.Q(axi_ARSIZE[1]));
	notech_nao3 i_4695(.A(n_62793), .B(1'b1), .C(axi_ARSIZE[1]), .Z(n_6513)
		);
	notech_reg axi_ARSIZE_reg_2(.CP(n_63292), .D(n_6517), .CD(n_62715), .Q(axi_ARSIZE
		[2]));
	notech_and2 i_4700(.A(n_62793), .B(axi_ARSIZE[2]), .Z(n_6517));
	notech_reg axi_AWLEN_reg_0(.CP(n_63292), .D(n_6523), .CD(n_62714), .Q(axi_AWLEN
		[0]));
	notech_and4 i_4708(.A(n_62793), .B(n_8323), .C(n_62820), .D(axi_AWLEN[0]
		), .Z(n_6523));
	notech_and3 i_44(.A(axi_RVALID), .B(n_2035), .C(n_62714), .Z(n_210756365
		));
	notech_reg axi_AWLEN_reg_1(.CP(n_63292), .D(n_6529), .CD(n_62714), .Q(axi_AWLEN
		[1]));
	notech_and4 i_4716(.A(n_62793), .B(n_8323), .C(n_62820), .D(axi_AWLEN[1]
		), .Z(n_6529));
	notech_nao3 i_109(.A(n_2035), .B(n_62132), .C(n_2030), .Z(n_210856366)
		);
	notech_reg axi_AWLEN_reg_2(.CP(n_63292), .D(n_6535), .CD(n_62714), .Q(axi_AWLEN
		[2]));
	notech_and4 i_4724(.A(n_62793), .B(n_8323), .C(n_62820), .D(axi_AWLEN[2]
		), .Z(n_6535));
	notech_reg axi_AWLEN_reg_3(.CP(n_63292), .D(n_6541), .CD(n_62714), .Q(axi_AWLEN
		[3]));
	notech_and4 i_4732(.A(n_62788), .B(n_8323), .C(n_62820), .D(axi_AWLEN[3]
		), .Z(n_6541));
	notech_reg axi_AWLEN_reg_4(.CP(n_63292), .D(n_6547), .CD(n_62714), .Q(axi_AWLEN
		[4]));
	notech_and4 i_4740(.A(n_62788), .B(n_8323), .C(n_62820), .D(axi_AWLEN[4]
		), .Z(n_6547));
	notech_reg axi_AWLEN_reg_5(.CP(n_63292), .D(n_6553), .CD(n_62714), .Q(axi_AWLEN
		[5]));
	notech_and4 i_4748(.A(n_62788), .B(n_8323), .C(n_62820), .D(axi_AWLEN[5]
		), .Z(n_6553));
	notech_reg axi_AWLEN_reg_6(.CP(n_63292), .D(n_6559), .CD(n_62714), .Q(axi_AWLEN
		[6]));
	notech_and4 i_4756(.A(n_62788), .B(n_8323), .C(n_62820), .D(axi_AWLEN[6]
		), .Z(n_6559));
	notech_reg axi_AWLEN_reg_7(.CP(n_63292), .D(n_6565), .CD(n_62715), .Q(axi_AWLEN
		[7]));
	notech_and4 i_4764(.A(n_62788), .B(n_8323), .C(n_62820), .D(axi_AWLEN[7]
		), .Z(n_6565));
	notech_reg axi_WLAST_reg(.CP(n_63292), .D(n_6568), .CD(n_62716), .Q(axi_WLAST
		));
	notech_mux2 i_4770(.S(n_62777), .A(n_1176), .B(axi_WLAST), .Z(n_6568));
	notech_reg axi_ARLEN_reg_0(.CP(n_63292), .D(n_6574), .CD(n_62716), .Q(axi_ARLEN
		[0]));
	notech_mux2 i_4778(.S(n_62150), .A(n_8226), .B(axi_ARLEN[0]), .Z(n_6574)
		);
	notech_reg axi_ARLEN_reg_1(.CP(n_63292), .D(n_6580), .CD(n_62716), .Q(axi_ARLEN
		[1]));
	notech_mux2 i_4786(.S(n_62150), .A(n_8226), .B(axi_ARLEN[1]), .Z(n_6580)
		);
	notech_reg axi_ARLEN_reg_2(.CP(n_63292), .D(n_6589), .CD(n_62716), .Q(axi_ARLEN
		[2]));
	notech_and4 i_4796(.A(n_62788), .B(n_1066), .C(axi_ARLEN[2]), .D(n_973),
		 .Z(n_6589));
	notech_reg axi_ARLEN_reg_3(.CP(n_63292), .D(n_6595), .CD(n_62716), .Q(axi_ARLEN
		[3]));
	notech_and4 i_4804(.A(n_62788), .B(n_1066), .C(axi_ARLEN[3]), .D(n_973),
		 .Z(n_6595));
	notech_reg axi_ARLEN_reg_4(.CP(n_63292), .D(n_6601), .CD(n_62716), .Q(axi_ARLEN
		[4]));
	notech_and4 i_4812(.A(n_62788), .B(n_1066), .C(axi_ARLEN[4]), .D(n_973),
		 .Z(n_6601));
	notech_reg axi_ARLEN_reg_5(.CP(n_63300), .D(n_6607), .CD(n_62716), .Q(axi_ARLEN
		[5]));
	notech_and4 i_4820(.A(n_62788), .B(n_1066), .C(axi_ARLEN[5]), .D(n_973),
		 .Z(n_6607));
	notech_reg axi_ARLEN_reg_6(.CP(n_63284), .D(n_6613), .CD(n_62716), .Q(axi_ARLEN
		[6]));
	notech_and4 i_4828(.A(n_62788), .B(n_1066), .C(axi_ARLEN[6]), .D(n_973),
		 .Z(n_6613));
	notech_reg axi_ARLEN_reg_7(.CP(n_63284), .D(n_6619), .CD(n_62715), .Q(axi_ARLEN
		[7]));
	notech_and4 i_4836(.A(n_62788), .B(n_1066), .C(axi_ARLEN[7]), .D(n_973),
		 .Z(n_6619));
	notech_reg axi_io_AR_reg_0(.CP(n_63284), .D(n_6625), .CD(n_62715), .Q(axi_io_AR
		[0]));
	notech_and2 i_4844(.A(axi_io_AR[0]), .B(n_8331), .Z(n_6625));
	notech_reg axi_io_AR_reg_1(.CP(n_63284), .D(n_6631), .CD(n_62715), .Q(axi_io_AR
		[1]));
	notech_and2 i_4852(.A(n_8331), .B(axi_io_AR[1]), .Z(n_6631));
	notech_reg axi_io_AR_reg_2(.CP(n_63284), .D(n_6634), .CD(n_62715), .Q(axi_io_AR
		[2]));
	notech_mux2 i_4858(.S(\nbus_11673[0] ), .A(axi_io_AR[2]), .B(io_add[0]),
		 .Z(n_6634));
	notech_reg axi_io_AR_reg_3(.CP(n_63284), .D(n_6640), .CD(n_62715), .Q(axi_io_AR
		[3]));
	notech_mux2 i_4866(.S(\nbus_11673[0] ), .A(axi_io_AR[3]), .B(io_add[1]),
		 .Z(n_6640));
	notech_reg axi_io_AR_reg_4(.CP(n_63284), .D(n_6646), .CD(n_62715), .Q(axi_io_AR
		[4]));
	notech_mux2 i_4874(.S(\nbus_11673[0] ), .A(axi_io_AR[4]), .B(io_add[2]),
		 .Z(n_6646));
	notech_reg axi_io_AR_reg_5(.CP(n_63284), .D(n_6652), .CD(n_62715), .Q(axi_io_AR
		[5]));
	notech_mux2 i_4882(.S(\nbus_11673[0] ), .A(axi_io_AR[5]), .B(io_add[3]),
		 .Z(n_6652));
	notech_reg axi_io_AR_reg_6(.CP(n_63284), .D(n_6658), .CD(n_62715), .Q(axi_io_AR
		[6]));
	notech_mux2 i_4890(.S(\nbus_11673[0] ), .A(axi_io_AR[6]), .B(io_add[4]),
		 .Z(n_6658));
	notech_reg axi_io_AR_reg_7(.CP(n_63284), .D(n_6664), .CD(n_62714), .Q(axi_io_AR
		[7]));
	notech_mux2 i_4898(.S(\nbus_11673[0] ), .A(axi_io_AR[7]), .B(io_add[5]),
		 .Z(n_6664));
	notech_reg axi_io_AR_reg_8(.CP(n_63284), .D(n_6670), .CD(n_62712), .Q(axi_io_AR
		[8]));
	notech_mux2 i_4906(.S(\nbus_11673[0] ), .A(axi_io_AR[8]), .B(io_add[6]),
		 .Z(n_6670));
	notech_reg axi_io_AR_reg_9(.CP(n_63284), .D(n_6676), .CD(n_62712), .Q(axi_io_AR
		[9]));
	notech_mux2 i_4914(.S(\nbus_11673[0] ), .A(axi_io_AR[9]), .B(io_add[7]),
		 .Z(n_6676));
	notech_reg axi_io_AR_reg_10(.CP(n_63284), .D(n_6682), .CD(n_62712), .Q(axi_io_AR
		[10]));
	notech_mux2 i_4922(.S(\nbus_11673[0] ), .A(axi_io_AR[10]), .B(io_add[8])
		, .Z(n_6682));
	notech_reg axi_io_AR_reg_11(.CP(n_63284), .D(n_6688), .CD(n_62712), .Q(axi_io_AR
		[11]));
	notech_mux2 i_4930(.S(\nbus_11673[0] ), .A(axi_io_AR[11]), .B(io_add[9])
		, .Z(n_6688));
	notech_reg axi_io_AR_reg_12(.CP(n_63284), .D(n_6694), .CD(n_62713), .Q(axi_io_AR
		[12]));
	notech_mux2 i_4938(.S(\nbus_11673[0] ), .A(axi_io_AR[12]), .B(io_add[10]
		), .Z(n_6694));
	notech_reg axi_io_AR_reg_13(.CP(n_63304), .D(n_6700), .CD(n_62713), .Q(axi_io_AR
		[13]));
	notech_mux2 i_4946(.S(\nbus_11673[0] ), .A(axi_io_AR[13]), .B(io_add[11]
		), .Z(n_6700));
	notech_reg axi_io_AR_reg_14(.CP(n_63304), .D(n_6706), .CD(n_62712), .Q(axi_io_AR
		[14]));
	notech_mux2 i_4954(.S(\nbus_11673[0] ), .A(axi_io_AR[14]), .B(io_add[12]
		), .Z(n_6706));
	notech_reg axi_io_AR_reg_15(.CP(n_63304), .D(n_6712), .CD(n_62712), .Q(axi_io_AR
		[15]));
	notech_mux2 i_4962(.S(\nbus_11673[0] ), .A(axi_io_AR[15]), .B(io_add[13]
		), .Z(n_6712));
	notech_reg axi_io_AR_reg_16(.CP(n_63304), .D(n_6718), .CD(n_62712), .Q(axi_io_AR
		[16]));
	notech_mux2 i_4970(.S(\nbus_11673[0] ), .A(axi_io_AR[16]), .B(io_add[14]
		), .Z(n_6718));
	notech_reg axi_io_AR_reg_17(.CP(n_63304), .D(n_6724), .CD(n_62712), .Q(axi_io_AR
		[17]));
	notech_mux2 i_4978(.S(\nbus_11673[0] ), .A(axi_io_AR[17]), .B(io_add[15]
		), .Z(n_6724));
	notech_reg axi_io_AR_reg_18(.CP(n_63304), .D(n_6733), .CD(n_62712), .Q(axi_io_AR
		[18]));
	notech_and2 i_4988(.A(axi_io_AR[18]), .B(n_8331), .Z(n_6733));
	notech_ao3 i_36(.A(n_2069), .B(n_60720), .C(n_60789), .Z(n_214256400));
	notech_reg axi_io_AR_reg_19(.CP(n_63304), .D(n_6739), .CD(n_62712), .Q(axi_io_AR
		[19]));
	notech_and2 i_4996(.A(axi_io_AR[19]), .B(n_8331), .Z(n_6739));
	notech_ao3 i_34(.A(n_2069), .B(n_60755), .C(n_60789), .Z(n_214356401));
	notech_reg axi_io_AR_reg_20(.CP(n_63304), .D(n_6745), .CD(n_62712), .Q(axi_io_AR
		[20]));
	notech_and2 i_5004(.A(axi_io_AR[20]), .B(n_8331), .Z(n_6745));
	notech_reg axi_io_AR_reg_21(.CP(n_63304), .D(n_6751), .CD(n_62712), .Q(axi_io_AR
		[21]));
	notech_and2 i_5012(.A(axi_io_AR[21]), .B(n_8331), .Z(n_6751));
	notech_reg axi_io_AR_reg_22(.CP(n_63304), .D(n_6757), .CD(n_62712), .Q(axi_io_AR
		[22]));
	notech_and2 i_5020(.A(axi_io_AR[22]), .B(n_8331), .Z(n_6757));
	notech_reg axi_io_AR_reg_23(.CP(n_63304), .D(n_6763), .CD(n_62712), .Q(axi_io_AR
		[23]));
	notech_and2 i_5028(.A(axi_io_AR[23]), .B(n_8331), .Z(n_6763));
	notech_reg axi_io_AR_reg_24(.CP(n_63304), .D(n_6769), .CD(n_62713), .Q(axi_io_AR
		[24]));
	notech_and2 i_5036(.A(axi_io_AR[24]), .B(n_8331), .Z(n_6769));
	notech_reg axi_io_AR_reg_25(.CP(n_63304), .D(n_6775), .CD(n_62713), .Q(axi_io_AR
		[25]));
	notech_and2 i_5044(.A(axi_io_AR[25]), .B(n_8331), .Z(n_6775));
	notech_reg axi_io_AR_reg_26(.CP(n_63304), .D(n_6781), .CD(n_62713), .Q(axi_io_AR
		[26]));
	notech_and2 i_5052(.A(axi_io_AR[26]), .B(n_8331), .Z(n_6781));
	notech_reg axi_io_AR_reg_27(.CP(n_63304), .D(n_6787), .CD(n_62713), .Q(axi_io_AR
		[27]));
	notech_and2 i_5060(.A(axi_io_AR[27]), .B(n_8331), .Z(n_6787));
	notech_reg axi_io_AR_reg_28(.CP(n_63304), .D(n_6793), .CD(n_62713), .Q(axi_io_AR
		[28]));
	notech_and2 i_5068(.A(axi_io_AR[28]), .B(n_8331), .Z(n_6793));
	notech_reg axi_io_AR_reg_29(.CP(n_63304), .D(n_6799), .CD(n_62714), .Q(axi_io_AR
		[29]));
	notech_and2 i_5076(.A(axi_io_AR[29]), .B(n_8331), .Z(n_6799));
	notech_reg axi_io_AR_reg_30(.CP(n_63304), .D(n_6805), .CD(n_62714), .Q(axi_io_AR
		[30]));
	notech_and2 i_5084(.A(axi_io_AR[30]), .B(n_8331), .Z(n_6805));
	notech_reg axi_io_AR_reg_31(.CP(n_63304), .D(n_6811), .CD(n_62714), .Q(axi_io_AR
		[31]));
	notech_and2 i_5092(.A(axi_io_AR[31]), .B(n_8331), .Z(n_6811));
	notech_reg_set readio_data_reg_0(.CP(n_63302), .D(n_6814), .SD(1'b1), .Q
		(readio_data[0]));
	notech_mux2 i_5098(.S(\nbus_11671[0] ), .A(readio_data[0]), .B(axi_io_R[
		0]), .Z(n_6814));
	notech_reg_set readio_data_reg_1(.CP(n_63302), .D(n_6820), .SD(1'b1), .Q
		(readio_data[1]));
	notech_mux2 i_5106(.S(\nbus_11671[0] ), .A(readio_data[1]), .B(axi_io_R[
		1]), .Z(n_6820));
	notech_reg_set readio_data_reg_2(.CP(n_63328), .D(n_6826), .SD(1'b1), .Q
		(readio_data[2]));
	notech_mux2 i_5114(.S(\nbus_11671[0] ), .A(readio_data[2]), .B(axi_io_R[
		2]), .Z(n_6826));
	notech_reg_set readio_data_reg_3(.CP(n_63328), .D(n_6832), .SD(1'b1), .Q
		(readio_data[3]));
	notech_mux2 i_5122(.S(\nbus_11671[0] ), .A(readio_data[3]), .B(axi_io_R[
		3]), .Z(n_6832));
	notech_reg_set readio_data_reg_4(.CP(n_63328), .D(n_6838), .SD(1'b1), .Q
		(readio_data[4]));
	notech_mux2 i_5130(.S(\nbus_11671[0] ), .A(readio_data[4]), .B(axi_io_R[
		4]), .Z(n_6838));
	notech_reg_set readio_data_reg_5(.CP(n_63328), .D(n_6844), .SD(1'b1), .Q
		(readio_data[5]));
	notech_mux2 i_5138(.S(\nbus_11671[0] ), .A(readio_data[5]), .B(axi_io_R[
		5]), .Z(n_6844));
	notech_reg_set readio_data_reg_6(.CP(n_63328), .D(n_6850), .SD(1'b1), .Q
		(readio_data[6]));
	notech_mux2 i_5146(.S(\nbus_11671[0] ), .A(readio_data[6]), .B(axi_io_R[
		6]), .Z(n_6850));
	notech_reg_set readio_data_reg_7(.CP(n_63328), .D(n_6856), .SD(1'b1), .Q
		(readio_data[7]));
	notech_mux2 i_5154(.S(\nbus_11671[0] ), .A(readio_data[7]), .B(axi_io_R[
		7]), .Z(n_6856));
	notech_reg_set readio_data_reg_8(.CP(n_63328), .D(n_6862), .SD(1'b1), .Q
		(readio_data[8]));
	notech_mux2 i_5162(.S(\nbus_11671[0] ), .A(readio_data[8]), .B(axi_io_R[
		8]), .Z(n_6862));
	notech_reg_set readio_data_reg_9(.CP(n_63328), .D(n_6868), .SD(1'b1), .Q
		(readio_data[9]));
	notech_mux2 i_5170(.S(\nbus_11671[0] ), .A(readio_data[9]), .B(axi_io_R[
		9]), .Z(n_6868));
	notech_reg_set readio_data_reg_10(.CP(n_63328), .D(n_6874), .SD(1'b1), .Q
		(readio_data[10]));
	notech_mux2 i_5178(.S(\nbus_11671[0] ), .A(readio_data[10]), .B(axi_io_R
		[10]), .Z(n_6874));
	notech_reg_set readio_data_reg_11(.CP(n_63328), .D(n_6880), .SD(1'b1), .Q
		(readio_data[11]));
	notech_mux2 i_5186(.S(\nbus_11671[0] ), .A(readio_data[11]), .B(axi_io_R
		[11]), .Z(n_6880));
	notech_reg_set readio_data_reg_12(.CP(n_63328), .D(n_6886), .SD(1'b1), .Q
		(readio_data[12]));
	notech_mux2 i_5194(.S(\nbus_11671[0] ), .A(readio_data[12]), .B(axi_io_R
		[12]), .Z(n_6886));
	notech_reg_set readio_data_reg_13(.CP(n_63328), .D(n_6892), .SD(1'b1), .Q
		(readio_data[13]));
	notech_mux2 i_5202(.S(\nbus_11671[0] ), .A(readio_data[13]), .B(axi_io_R
		[13]), .Z(n_6892));
	notech_reg_set readio_data_reg_14(.CP(n_63328), .D(n_6898), .SD(1'b1), .Q
		(readio_data[14]));
	notech_mux2 i_5210(.S(\nbus_11671[0] ), .A(readio_data[14]), .B(axi_io_R
		[14]), .Z(n_6898));
	notech_reg_set readio_data_reg_15(.CP(n_63328), .D(n_6904), .SD(1'b1), .Q
		(readio_data[15]));
	notech_mux2 i_5218(.S(\nbus_11671[0] ), .A(readio_data[15]), .B(axi_io_R
		[15]), .Z(n_6904));
	notech_reg_set readio_data_reg_16(.CP(n_63328), .D(n_6910), .SD(1'b1), .Q
		(readio_data[16]));
	notech_mux2 i_5226(.S(n_56052), .A(readio_data[16]), .B(axi_io_R[16]), .Z
		(n_6910));
	notech_reg_set readio_data_reg_17(.CP(n_63328), .D(n_6916), .SD(1'b1), .Q
		(readio_data[17]));
	notech_mux2 i_5234(.S(n_56052), .A(readio_data[17]), .B(axi_io_R[17]), .Z
		(n_6916));
	notech_reg_set readio_data_reg_18(.CP(n_63328), .D(n_6922), .SD(1'b1), .Q
		(readio_data[18]));
	notech_mux2 i_5242(.S(n_56052), .A(readio_data[18]), .B(axi_io_R[18]), .Z
		(n_6922));
	notech_reg_set readio_data_reg_19(.CP(n_63328), .D(n_6928), .SD(1'b1), .Q
		(readio_data[19]));
	notech_mux2 i_5250(.S(n_56052), .A(readio_data[19]), .B(axi_io_R[19]), .Z
		(n_6928));
	notech_reg_set readio_data_reg_20(.CP(n_63302), .D(n_6934), .SD(1'b1), .Q
		(readio_data[20]));
	notech_mux2 i_5258(.S(n_56052), .A(readio_data[20]), .B(axi_io_R[20]), .Z
		(n_6934));
	notech_reg_set readio_data_reg_21(.CP(n_63302), .D(n_6940), .SD(1'b1), .Q
		(readio_data[21]));
	notech_mux2 i_5266(.S(n_56052), .A(readio_data[21]), .B(axi_io_R[21]), .Z
		(n_6940));
	notech_reg_set readio_data_reg_22(.CP(n_63302), .D(n_6946), .SD(1'b1), .Q
		(readio_data[22]));
	notech_mux2 i_5274(.S(n_56052), .A(readio_data[22]), .B(axi_io_R[22]), .Z
		(n_6946));
	notech_reg_set readio_data_reg_23(.CP(n_63302), .D(n_6952), .SD(1'b1), .Q
		(readio_data[23]));
	notech_mux2 i_5282(.S(n_56052), .A(readio_data[23]), .B(axi_io_R[23]), .Z
		(n_6952));
	notech_reg_set readio_data_reg_24(.CP(n_63302), .D(n_6958), .SD(1'b1), .Q
		(readio_data[24]));
	notech_mux2 i_5290(.S(n_56052), .A(readio_data[24]), .B(axi_io_R[24]), .Z
		(n_6958));
	notech_reg_set readio_data_reg_25(.CP(n_63302), .D(n_6964), .SD(1'b1), .Q
		(readio_data[25]));
	notech_mux2 i_5298(.S(n_56052), .A(readio_data[25]), .B(axi_io_R[25]), .Z
		(n_6964));
	notech_reg_set readio_data_reg_26(.CP(n_63302), .D(n_6970), .SD(1'b1), .Q
		(readio_data[26]));
	notech_mux2 i_5306(.S(n_56052), .A(readio_data[26]), .B(axi_io_R[26]), .Z
		(n_6970));
	notech_reg_set readio_data_reg_27(.CP(n_63302), .D(n_6976), .SD(1'b1), .Q
		(readio_data[27]));
	notech_mux2 i_5314(.S(n_56052), .A(readio_data[27]), .B(axi_io_R[27]), .Z
		(n_6976));
	notech_reg_set readio_data_reg_28(.CP(n_63302), .D(n_6982), .SD(1'b1), .Q
		(readio_data[28]));
	notech_mux2 i_5322(.S(n_56052), .A(readio_data[28]), .B(axi_io_R[28]), .Z
		(n_6982));
	notech_reg_set readio_data_reg_29(.CP(n_63302), .D(n_6988), .SD(1'b1), .Q
		(readio_data[29]));
	notech_mux2 i_5330(.S(n_56052), .A(readio_data[29]), .B(axi_io_R[29]), .Z
		(n_6988));
	notech_reg_set readio_data_reg_30(.CP(n_63302), .D(n_6994), .SD(1'b1), .Q
		(readio_data[30]));
	notech_mux2 i_5338(.S(n_56052), .A(readio_data[30]), .B(axi_io_R[30]), .Z
		(n_6994));
	notech_reg_set readio_data_reg_31(.CP(n_63302), .D(n_7000), .SD(1'b1), .Q
		(readio_data[31]));
	notech_mux2 i_5346(.S(n_56052), .A(readio_data[31]), .B(axi_io_R[31]), .Z
		(n_7000));
	notech_reg axi_AWSIZE_reg_0(.CP(n_63302), .D(n_7009), .CD(n_62714), .Q(axi_AWSIZE
		[0]));
	notech_and2 i_5356(.A(n_62793), .B(axi_AWSIZE[0]), .Z(n_7009));
	notech_reg_set axi_AWSIZE_reg_1(.CP(n_63302), .D(n_7017), .SD(n_62713), 
		.Q(axi_AWSIZE[1]));
	notech_nao3 i_5367(.A(n_62788), .B(1'b1), .C(axi_AWSIZE[1]), .Z(n_7017)
		);
	notech_reg axi_AWSIZE_reg_2(.CP(n_63302), .D(n_7021), .CD(n_62713), .Q(axi_AWSIZE
		[2]));
	notech_and2 i_5372(.A(n_62788), .B(axi_AWSIZE[2]), .Z(n_7021));
	notech_reg_set axi_AWBURST_reg_0(.CP(n_63328), .D(n_7029), .SD(n_62713),
		 .Q(axi_AWBURST[0]));
	notech_nao3 i_5383(.A(n_62788), .B(1'b1), .C(axi_AWBURST[0]), .Z(n_7029)
		);
	notech_reg axi_AWBURST_reg_1(.CP(n_63324), .D(n_7033), .CD(n_62713), .Q(axi_AWBURST
		[1]));
	notech_and2 i_5388(.A(n_62788), .B(axi_AWBURST[1]), .Z(n_7033));
	notech_reg_set code_data_reg_0(.CP(n_63300), .D(n_7036), .SD(1'b1), .Q(\nbus_14547[0] 
		));
	notech_mux2 i_5394(.S(\nbus_11667[0] ), .A(n_61573), .B(axi_R[0]), .Z(n_7036
		));
	notech_reg_set code_data_reg_1(.CP(n_63324), .D(n_7042), .SD(1'b1), .Q(code_data
		[1]));
	notech_mux2 i_5402(.S(\nbus_11667[0] ), .A(code_data[1]), .B(axi_R[1]), 
		.Z(n_7042));
	notech_reg_set code_data_reg_2(.CP(n_63324), .D(n_7048), .SD(1'b1), .Q(code_data
		[2]));
	notech_mux2 i_5410(.S(\nbus_11667[0] ), .A(code_data[2]), .B(axi_R[2]), 
		.Z(n_7048));
	notech_reg_set code_data_reg_3(.CP(n_63324), .D(n_7054), .SD(1'b1), .Q(code_data
		[3]));
	notech_mux2 i_5418(.S(\nbus_11667[0] ), .A(code_data[3]), .B(axi_R[3]), 
		.Z(n_7054));
	notech_reg_set code_data_reg_4(.CP(n_63324), .D(n_7060), .SD(1'b1), .Q(code_data
		[4]));
	notech_mux2 i_5426(.S(\nbus_11667[0] ), .A(code_data[4]), .B(axi_R[4]), 
		.Z(n_7060));
	notech_reg_set code_data_reg_5(.CP(n_63324), .D(n_7066), .SD(1'b1), .Q(code_data
		[5]));
	notech_mux2 i_5434(.S(\nbus_11667[0] ), .A(code_data[5]), .B(axi_R[5]), 
		.Z(n_7066));
	notech_reg_set code_data_reg_6(.CP(n_63324), .D(n_7072), .SD(1'b1), .Q(code_data
		[6]));
	notech_mux2 i_5442(.S(\nbus_11667[0] ), .A(code_data[6]), .B(axi_R[6]), 
		.Z(n_7072));
	notech_reg_set code_data_reg_7(.CP(n_63324), .D(n_7078), .SD(1'b1), .Q(code_data
		[7]));
	notech_mux2 i_5450(.S(\nbus_11667[0] ), .A(code_data[7]), .B(axi_R[7]), 
		.Z(n_7078));
	notech_reg_set code_data_reg_8(.CP(n_63324), .D(n_7084), .SD(1'b1), .Q(code_data
		[8]));
	notech_mux2 i_5458(.S(\nbus_11667[0] ), .A(code_data[8]), .B(axi_R[8]), 
		.Z(n_7084));
	notech_reg_set code_data_reg_9(.CP(n_63324), .D(n_7090), .SD(1'b1), .Q(code_data
		[9]));
	notech_mux2 i_5466(.S(\nbus_11667[0] ), .A(code_data[9]), .B(axi_R[9]), 
		.Z(n_7090));
	notech_reg_set code_data_reg_10(.CP(n_63324), .D(n_7096), .SD(1'b1), .Q(code_data
		[10]));
	notech_mux2 i_5474(.S(\nbus_11667[0] ), .A(code_data[10]), .B(axi_R[10])
		, .Z(n_7096));
	notech_reg_set code_data_reg_11(.CP(n_63324), .D(n_7102), .SD(1'b1), .Q(code_data
		[11]));
	notech_mux2 i_5482(.S(\nbus_11667[0] ), .A(code_data[11]), .B(axi_R[11])
		, .Z(n_7102));
	notech_reg_set code_data_reg_12(.CP(n_63324), .D(n_7108), .SD(1'b1), .Q(code_data
		[12]));
	notech_mux2 i_5490(.S(\nbus_11667[0] ), .A(code_data[12]), .B(axi_R[12])
		, .Z(n_7108));
	notech_reg_set code_data_reg_13(.CP(n_63324), .D(n_7114), .SD(1'b1), .Q(code_data
		[13]));
	notech_mux2 i_5498(.S(\nbus_11667[0] ), .A(code_data[13]), .B(axi_R[13])
		, .Z(n_7114));
	notech_reg_set code_data_reg_14(.CP(n_63324), .D(n_7120), .SD(1'b1), .Q(code_data
		[14]));
	notech_mux2 i_5506(.S(\nbus_11667[0] ), .A(code_data[14]), .B(axi_R[14])
		, .Z(n_7120));
	notech_reg_set code_data_reg_15(.CP(n_63324), .D(n_7126), .SD(1'b1), .Q(code_data
		[15]));
	notech_mux2 i_5514(.S(\nbus_11667[0] ), .A(code_data[15]), .B(axi_R[15])
		, .Z(n_7126));
	notech_reg_set code_data_reg_16(.CP(n_63346), .D(n_7132), .SD(1'b1), .Q(code_data
		[16]));
	notech_mux2 i_5522(.S(n_57733), .A(code_data[16]), .B(axi_R[16]), .Z(n_7132
		));
	notech_ao3 i_1013(.A(n_2019), .B(n_1711), .C(n_1742), .Z(n_220956467));
	notech_reg_set code_data_reg_17(.CP(n_63346), .D(n_7138), .SD(1'b1), .Q(code_data
		[17]));
	notech_mux2 i_5530(.S(n_57733), .A(code_data[17]), .B(axi_R[17]), .Z(n_7138
		));
	notech_reg_set code_data_reg_18(.CP(n_63346), .D(n_7144), .SD(1'b1), .Q(code_data
		[18]));
	notech_mux2 i_5538(.S(n_57733), .A(code_data[18]), .B(axi_R[18]), .Z(n_7144
		));
	notech_reg_set code_data_reg_19(.CP(n_63346), .D(n_7150), .SD(1'b1), .Q(code_data
		[19]));
	notech_mux2 i_5546(.S(n_57733), .A(code_data[19]), .B(axi_R[19]), .Z(n_7150
		));
	notech_reg_set code_data_reg_20(.CP(n_63346), .D(n_7156), .SD(1'b1), .Q(code_data
		[20]));
	notech_mux2 i_5554(.S(n_57733), .A(code_data[20]), .B(axi_R[20]), .Z(n_7156
		));
	notech_reg_set code_data_reg_21(.CP(n_63346), .D(n_7162), .SD(1'b1), .Q(code_data
		[21]));
	notech_mux2 i_5562(.S(n_57733), .A(code_data[21]), .B(axi_R[21]), .Z(n_7162
		));
	notech_reg_set code_data_reg_22(.CP(n_63346), .D(n_7168), .SD(1'b1), .Q(code_data
		[22]));
	notech_mux2 i_5570(.S(n_57733), .A(code_data[22]), .B(axi_R[22]), .Z(n_7168
		));
	notech_reg_set code_data_reg_23(.CP(n_63346), .D(n_7174), .SD(1'b1), .Q(code_data
		[23]));
	notech_mux2 i_5578(.S(n_57733), .A(code_data[23]), .B(axi_R[23]), .Z(n_7174
		));
	notech_or4 i_1058(.A(n_1221), .B(n_974), .C(n_1748), .D(n_2033), .Z(n_221656474
		));
	notech_reg_set code_data_reg_24(.CP(n_63346), .D(n_7180), .SD(1'b1), .Q(code_data
		[24]));
	notech_mux2 i_5586(.S(n_57733), .A(code_data[24]), .B(axi_R[24]), .Z(n_7180
		));
	notech_reg_set code_data_reg_25(.CP(n_63346), .D(n_7186), .SD(1'b1), .Q(code_data
		[25]));
	notech_mux2 i_5594(.S(n_57733), .A(code_data[25]), .B(axi_R[25]), .Z(n_7186
		));
	notech_reg_set code_data_reg_26(.CP(n_63346), .D(n_7192), .SD(1'b1), .Q(code_data
		[26]));
	notech_mux2 i_5602(.S(n_57733), .A(code_data[26]), .B(axi_R[26]), .Z(n_7192
		));
	notech_ao4 i_58(.A(n_2045), .B(n_2052), .C(n_62123), .D(n_2016), .Z(n_221956477
		));
	notech_reg_set code_data_reg_27(.CP(n_63346), .D(n_7198), .SD(1'b1), .Q(code_data
		[27]));
	notech_mux2 i_5610(.S(n_57733), .A(code_data[27]), .B(axi_R[27]), .Z(n_7198
		));
	notech_reg_set code_data_reg_28(.CP(n_63346), .D(n_7204), .SD(1'b1), .Q(code_data
		[28]));
	notech_mux2 i_5618(.S(n_57733), .A(code_data[28]), .B(axi_R[28]), .Z(n_7204
		));
	notech_reg_set code_data_reg_29(.CP(n_63346), .D(n_7210), .SD(1'b1), .Q(code_data
		[29]));
	notech_mux2 i_5626(.S(n_57733), .A(code_data[29]), .B(axi_R[29]), .Z(n_7210
		));
	notech_reg_set code_data_reg_30(.CP(n_63346), .D(n_7216), .SD(1'b1), .Q(code_data
		[30]));
	notech_mux2 i_5634(.S(n_57733), .A(code_data[30]), .B(axi_R[30]), .Z(n_7216
		));
	notech_reg_set code_data_reg_31(.CP(n_63346), .D(n_7222), .SD(1'b1), .Q(code_data
		[31]));
	notech_mux2 i_5642(.S(n_57733), .A(code_data[31]), .B(axi_R[31]), .Z(n_7222
		));
	notech_or2 i_55(.A(readio_ack), .B(writeio_ack), .Z(n_222456482));
	notech_reg_set code_data_reg_32(.CP(n_63346), .D(n_7228), .SD(1'b1), .Q(code_data
		[32]));
	notech_mux2 i_5650(.S(\nbus_11667[32] ), .A(code_data[32]), .B(axi_R[0])
		, .Z(n_7228));
	notech_nao3 i_118(.A(n_8560), .B(n_8333), .C(readio_ack), .Z(n_222556483
		));
	notech_reg_set code_data_reg_33(.CP(n_63346), .D(n_7234), .SD(1'b1), .Q(code_data
		[33]));
	notech_mux2 i_5658(.S(\nbus_11667[32] ), .A(code_data[33]), .B(axi_R[1])
		, .Z(n_7234));
	notech_nand2 i_122(.A(axi_io_WVALID), .B(axi_io_WREADY), .Z(n_222656484)
		);
	notech_reg_set code_data_reg_34(.CP(n_63324), .D(n_7240), .SD(1'b1), .Q(code_data
		[34]));
	notech_mux2 i_5666(.S(\nbus_11667[32] ), .A(code_data[34]), .B(axi_R[2])
		, .Z(n_7240));
	notech_nao3 i_54(.A(n_222656484), .B(n_8333), .C(n_222456482), .Z(n_222756485
		));
	notech_reg_set code_data_reg_35(.CP(n_63346), .D(n_7246), .SD(1'b1), .Q(code_data
		[35]));
	notech_mux2 i_5674(.S(\nbus_11667[32] ), .A(code_data[35]), .B(axi_R[3])
		, .Z(n_7246));
	notech_ao3 i_63(.A(n_222656484), .B(n_8330), .C(n_222556483), .Z(n_222856486
		));
	notech_reg_set code_data_reg_36(.CP(n_63326), .D(n_7252), .SD(1'b1), .Q(code_data
		[36]));
	notech_mux2 i_5682(.S(\nbus_11667[32] ), .A(code_data[36]), .B(axi_R[4])
		, .Z(n_7252));
	notech_and2 i_75(.A(axi_io_RREADY), .B(axi_io_RVALID), .Z(n_222956487)
		);
	notech_reg_set code_data_reg_37(.CP(n_63326), .D(n_7258), .SD(1'b1), .Q(code_data
		[37]));
	notech_mux2 i_5690(.S(\nbus_11667[32] ), .A(code_data[37]), .B(axi_R[5])
		, .Z(n_7258));
	notech_nao3 i_66(.A(n_8330), .B(n_8219), .C(n_222756485), .Z(n_223056488
		));
	notech_reg_set code_data_reg_38(.CP(n_63326), .D(n_7264), .SD(1'b1), .Q(code_data
		[38]));
	notech_mux2 i_5698(.S(\nbus_11667[32] ), .A(code_data[38]), .B(axi_R[6])
		, .Z(n_7264));
	notech_nand2 i_23(.A(writeio_req), .B(n_8329), .Z(n_223156489));
	notech_reg_set code_data_reg_39(.CP(n_63326), .D(n_7270), .SD(1'b1), .Q(code_data
		[39]));
	notech_mux2 i_5706(.S(\nbus_11667[32] ), .A(code_data[39]), .B(axi_R[7])
		, .Z(n_7270));
	notech_reg_set code_data_reg_40(.CP(n_63326), .D(n_7276), .SD(1'b1), .Q(code_data
		[40]));
	notech_mux2 i_5714(.S(\nbus_11667[32] ), .A(code_data[40]), .B(axi_R[8])
		, .Z(n_7276));
	notech_nao3 i_1112(.A(readio_req), .B(n_223156489), .C(rf), .Z(n_223356491
		));
	notech_reg_set code_data_reg_41(.CP(n_63326), .D(n_7282), .SD(1'b1), .Q(code_data
		[41]));
	notech_mux2 i_5722(.S(\nbus_11667[32] ), .A(code_data[41]), .B(axi_R[9])
		, .Z(n_7282));
	notech_reg_set code_data_reg_42(.CP(n_63326), .D(n_7288), .SD(1'b1), .Q(code_data
		[42]));
	notech_mux2 i_5730(.S(\nbus_11667[32] ), .A(code_data[42]), .B(axi_R[10]
		), .Z(n_7288));
	notech_reg_set code_data_reg_43(.CP(n_63326), .D(n_7294), .SD(1'b1), .Q(code_data
		[43]));
	notech_mux2 i_5738(.S(\nbus_11667[32] ), .A(code_data[43]), .B(axi_R[11]
		), .Z(n_7294));
	notech_reg_set code_data_reg_44(.CP(n_63326), .D(n_7300), .SD(1'b1), .Q(code_data
		[44]));
	notech_mux2 i_5746(.S(\nbus_11667[32] ), .A(code_data[44]), .B(axi_R[12]
		), .Z(n_7300));
	notech_nand3 i_40(.A(n_60789), .B(n_62799), .C(n_60755), .Z(n_2237));
	notech_reg_set code_data_reg_45(.CP(n_63326), .D(n_7306), .SD(1'b1), .Q(code_data
		[45]));
	notech_mux2 i_5754(.S(\nbus_11667[32] ), .A(code_data[45]), .B(axi_R[13]
		), .Z(n_7306));
	notech_reg_set code_data_reg_46(.CP(n_63326), .D(n_7312), .SD(1'b1), .Q(code_data
		[46]));
	notech_mux2 i_5762(.S(\nbus_11667[32] ), .A(code_data[46]), .B(axi_R[14]
		), .Z(n_7312));
	notech_nao3 i_41(.A(n_62799), .B(n_60755), .C(n_60789), .Z(n_2239));
	notech_reg_set code_data_reg_47(.CP(n_63326), .D(n_7318), .SD(1'b1), .Q(code_data
		[47]));
	notech_mux2 i_5770(.S(\nbus_11667[32] ), .A(code_data[47]), .B(axi_R[15]
		), .Z(n_7318));
	notech_ao4 i_1164(.A(n_2239), .B(n_8475), .C(n_2237), .D(n_8507), .Z(n_2240
		));
	notech_reg_set code_data_reg_48(.CP(n_63326), .D(n_7324), .SD(1'b1), .Q(code_data
		[48]));
	notech_mux2 i_5778(.S(n_55679), .A(code_data[48]), .B(axi_R[16]), .Z(n_7324
		));
	notech_reg_set code_data_reg_49(.CP(n_63326), .D(n_7330), .SD(1'b1), .Q(code_data
		[49]));
	notech_mux2 i_5786(.S(n_55679), .A(code_data[49]), .B(axi_R[17]), .Z(n_7330
		));
	notech_reg_set code_data_reg_50(.CP(n_63326), .D(n_7336), .SD(1'b1), .Q(code_data
		[50]));
	notech_mux2 i_5794(.S(n_55679), .A(code_data[50]), .B(axi_R[18]), .Z(n_7336
		));
	notech_reg_set code_data_reg_51(.CP(n_63326), .D(n_7342), .SD(1'b1), .Q(code_data
		[51]));
	notech_mux2 i_5802(.S(n_55679), .A(code_data[51]), .B(axi_R[19]), .Z(n_7342
		));
	notech_nao3 i_38(.A(n_62799), .B(n_60720), .C(n_60789), .Z(n_2244));
	notech_reg_set code_data_reg_52(.CP(n_63326), .D(n_7348), .SD(1'b1), .Q(code_data
		[52]));
	notech_mux2 i_5810(.S(n_55679), .A(code_data[52]), .B(axi_R[20]), .Z(n_7348
		));
	notech_ao4 i_1163(.A(n_62799), .B(n_8335), .C(n_2244), .D(n_8443), .Z(n_2245
		));
	notech_reg_set code_data_reg_53(.CP(n_63326), .D(n_7354), .SD(1'b1), .Q(code_data
		[53]));
	notech_mux2 i_5818(.S(n_55679), .A(code_data[53]), .B(axi_R[21]), .Z(n_7354
		));
	notech_reg_set code_data_reg_54(.CP(n_63326), .D(n_7360), .SD(1'b1), .Q(code_data
		[54]));
	notech_mux2 i_5826(.S(n_55679), .A(code_data[54]), .B(axi_R[22]), .Z(n_7360
		));
	notech_ao4 i_1173(.A(n_2239), .B(n_8476), .C(n_2237), .D(n_8508), .Z(n_2247
		));
	notech_reg_set code_data_reg_55(.CP(n_63300), .D(n_7366), .SD(1'b1), .Q(code_data
		[55]));
	notech_mux2 i_5834(.S(n_55679), .A(code_data[55]), .B(axi_R[23]), .Z(n_7366
		));
	notech_ao4 i_1172(.A(n_62799), .B(n_8336), .C(n_2244), .D(n_8444), .Z(n_2248
		));
	notech_reg_set code_data_reg_56(.CP(n_63300), .D(n_7372), .SD(1'b1), .Q(code_data
		[56]));
	notech_mux2 i_5842(.S(n_55679), .A(code_data[56]), .B(axi_R[24]), .Z(n_7372
		));
	notech_reg_set code_data_reg_57(.CP(n_63300), .D(n_7378), .SD(1'b1), .Q(code_data
		[57]));
	notech_mux2 i_5850(.S(n_55679), .A(code_data[57]), .B(axi_R[25]), .Z(n_7378
		));
	notech_ao4 i_1182(.A(n_2239), .B(n_8477), .C(n_2237), .D(n_8509), .Z(n_2250
		));
	notech_reg_set code_data_reg_58(.CP(n_63300), .D(n_7384), .SD(1'b1), .Q(code_data
		[58]));
	notech_mux2 i_5858(.S(n_55679), .A(code_data[58]), .B(axi_R[26]), .Z(n_7384
		));
	notech_ao4 i_1181(.A(n_62804), .B(n_8337), .C(n_2244), .D(n_8445), .Z(n_2251
		));
	notech_reg_set code_data_reg_59(.CP(n_63300), .D(n_7390), .SD(1'b1), .Q(code_data
		[59]));
	notech_mux2 i_5866(.S(n_55679), .A(code_data[59]), .B(axi_R[27]), .Z(n_7390
		));
	notech_reg_set code_data_reg_60(.CP(n_63300), .D(n_7396), .SD(1'b1), .Q(code_data
		[60]));
	notech_mux2 i_5874(.S(n_55679), .A(code_data[60]), .B(axi_R[28]), .Z(n_7396
		));
	notech_ao4 i_1191(.A(n_2239), .B(n_8478), .C(n_2237), .D(n_8510), .Z(n_2253
		));
	notech_reg_set code_data_reg_61(.CP(n_63284), .D(n_7402), .SD(1'b1), .Q(code_data
		[61]));
	notech_mux2 i_5882(.S(n_55679), .A(code_data[61]), .B(axi_R[29]), .Z(n_7402
		));
	notech_ao4 i_1190(.A(n_62799), .B(n_8338), .C(n_2244), .D(n_8446), .Z(n_2254
		));
	notech_reg_set code_data_reg_62(.CP(n_63300), .D(n_7408), .SD(1'b1), .Q(code_data
		[62]));
	notech_mux2 i_5890(.S(n_55679), .A(code_data[62]), .B(axi_R[30]), .Z(n_7408
		));
	notech_reg_set code_data_reg_63(.CP(n_63300), .D(n_7414), .SD(1'b1), .Q(code_data
		[63]));
	notech_mux2 i_5898(.S(n_55679), .A(code_data[63]), .B(axi_R[31]), .Z(n_7414
		));
	notech_ao4 i_1200(.A(n_2239), .B(n_8479), .C(n_2237), .D(n_8511), .Z(n_2256
		));
	notech_reg_set code_data_reg_64(.CP(n_63300), .D(n_7420), .SD(1'b1), .Q(code_data
		[64]));
	notech_mux2 i_5906(.S(\nbus_11667[64] ), .A(code_data[64]), .B(axi_R[0])
		, .Z(n_7420));
	notech_ao4 i_1199(.A(n_62799), .B(n_8339), .C(n_2244), .D(n_8447), .Z(n_2257
		));
	notech_reg_set code_data_reg_65(.CP(n_63300), .D(n_7426), .SD(1'b1), .Q(code_data
		[65]));
	notech_mux2 i_5914(.S(\nbus_11667[64] ), .A(code_data[65]), .B(axi_R[1])
		, .Z(n_7426));
	notech_reg_set code_data_reg_66(.CP(n_63300), .D(n_7432), .SD(1'b1), .Q(code_data
		[66]));
	notech_mux2 i_5922(.S(\nbus_11667[64] ), .A(code_data[66]), .B(axi_R[2])
		, .Z(n_7432));
	notech_ao4 i_1209(.A(n_2239), .B(n_8480), .C(n_2237), .D(n_8512), .Z(n_2259
		));
	notech_reg_set code_data_reg_67(.CP(n_63300), .D(n_7438), .SD(1'b1), .Q(code_data
		[67]));
	notech_mux2 i_5930(.S(\nbus_11667[64] ), .A(code_data[67]), .B(axi_R[3])
		, .Z(n_7438));
	notech_ao4 i_1208(.A(n_62799), .B(n_8340), .C(n_2244), .D(n_8448), .Z(n_2260
		));
	notech_reg_set code_data_reg_68(.CP(n_63300), .D(n_7444), .SD(1'b1), .Q(code_data
		[68]));
	notech_mux2 i_5938(.S(\nbus_11667[64] ), .A(code_data[68]), .B(axi_R[4])
		, .Z(n_7444));
	notech_reg_set code_data_reg_69(.CP(n_63300), .D(n_7450), .SD(1'b1), .Q(code_data
		[69]));
	notech_mux2 i_5946(.S(\nbus_11667[64] ), .A(code_data[69]), .B(axi_R[5])
		, .Z(n_7450));
	notech_ao4 i_1218(.A(n_2239), .B(n_8481), .C(n_2237), .D(n_8513), .Z(n_2262
		));
	notech_reg_set code_data_reg_70(.CP(n_63284), .D(n_7456), .SD(1'b1), .Q(code_data
		[70]));
	notech_mux2 i_5954(.S(\nbus_11667[64] ), .A(code_data[70]), .B(axi_R[6])
		, .Z(n_7456));
	notech_ao4 i_1217(.A(n_62799), .B(n_8341), .C(n_2244), .D(n_8449), .Z(n_2263
		));
	notech_reg_set code_data_reg_71(.CP(n_63300), .D(n_7462), .SD(1'b1), .Q(code_data
		[71]));
	notech_mux2 i_5962(.S(\nbus_11667[64] ), .A(code_data[71]), .B(axi_R[7])
		, .Z(n_7462));
	notech_reg_set code_data_reg_72(.CP(n_63306), .D(n_7468), .SD(1'b1), .Q(code_data
		[72]));
	notech_mux2 i_5970(.S(\nbus_11667[64] ), .A(code_data[72]), .B(axi_R[8])
		, .Z(n_7468));
	notech_ao4 i_1227(.A(n_2239), .B(n_8482), .C(n_2237), .D(n_8514), .Z(n_2265
		));
	notech_reg_set code_data_reg_73(.CP(n_63286), .D(n_7474), .SD(1'b1), .Q(code_data
		[73]));
	notech_mux2 i_5978(.S(\nbus_11667[64] ), .A(code_data[73]), .B(axi_R[9])
		, .Z(n_7474));
	notech_ao4 i_1226(.A(n_62799), .B(n_8342), .C(n_2244), .D(n_8450), .Z(n_2266
		));
	notech_reg_set code_data_reg_74(.CP(n_63286), .D(n_7480), .SD(1'b1), .Q(code_data
		[74]));
	notech_mux2 i_5986(.S(\nbus_11667[64] ), .A(code_data[74]), .B(axi_R[10]
		), .Z(n_7480));
	notech_reg_set code_data_reg_75(.CP(n_63286), .D(n_7486), .SD(1'b1), .Q(code_data
		[75]));
	notech_mux2 i_5994(.S(\nbus_11667[64] ), .A(code_data[75]), .B(axi_R[11]
		), .Z(n_7486));
	notech_ao4 i_1236(.A(n_2239), .B(n_8483), .C(n_2237), .D(n_8515), .Z(n_2268
		));
	notech_reg_set code_data_reg_76(.CP(n_63286), .D(n_7492), .SD(1'b1), .Q(code_data
		[76]));
	notech_mux2 i_6002(.S(\nbus_11667[64] ), .A(code_data[76]), .B(axi_R[12]
		), .Z(n_7492));
	notech_ao4 i_1235(.A(n_62799), .B(n_8343), .C(n_2244), .D(n_8451), .Z(n_2269
		));
	notech_reg_set code_data_reg_77(.CP(n_63286), .D(n_7498), .SD(1'b1), .Q(code_data
		[77]));
	notech_mux2 i_6010(.S(\nbus_11667[64] ), .A(code_data[77]), .B(axi_R[13]
		), .Z(n_7498));
	notech_reg_set code_data_reg_78(.CP(n_63286), .D(n_7504), .SD(1'b1), .Q(code_data
		[78]));
	notech_mux2 i_6018(.S(\nbus_11667[64] ), .A(code_data[78]), .B(axi_R[14]
		), .Z(n_7504));
	notech_ao4 i_1245(.A(n_2239), .B(n_8484), .C(n_2237), .D(n_8516), .Z(n_2271
		));
	notech_reg_set code_data_reg_79(.CP(n_63286), .D(n_7510), .SD(1'b1), .Q(code_data
		[79]));
	notech_mux2 i_6026(.S(\nbus_11667[64] ), .A(code_data[79]), .B(axi_R[15]
		), .Z(n_7510));
	notech_ao4 i_1244(.A(n_62799), .B(n_8344), .C(n_2244), .D(n_8452), .Z(n_2272
		));
	notech_reg_set code_data_reg_80(.CP(n_63286), .D(n_7516), .SD(1'b1), .Q(code_data
		[80]));
	notech_mux2 i_6034(.S(n_55668), .A(code_data[80]), .B(axi_R[16]), .Z(n_7516
		));
	notech_reg_set code_data_reg_81(.CP(n_63286), .D(n_7522), .SD(1'b1), .Q(code_data
		[81]));
	notech_mux2 i_6042(.S(n_55668), .A(code_data[81]), .B(axi_R[17]), .Z(n_7522
		));
	notech_ao4 i_1254(.A(n_2239), .B(n_8485), .C(n_2237), .D(n_8517), .Z(n_2274
		));
	notech_reg_set code_data_reg_82(.CP(n_63286), .D(n_7528), .SD(1'b1), .Q(code_data
		[82]));
	notech_mux2 i_6050(.S(n_55668), .A(code_data[82]), .B(axi_R[18]), .Z(n_7528
		));
	notech_ao4 i_1253(.A(n_62799), .B(n_8345), .C(n_2244), .D(n_8453), .Z(n_2275
		));
	notech_reg_set code_data_reg_83(.CP(n_63308), .D(n_7534), .SD(1'b1), .Q(code_data
		[83]));
	notech_mux2 i_6058(.S(n_55668), .A(code_data[83]), .B(axi_R[19]), .Z(n_7534
		));
	notech_reg_set code_data_reg_84(.CP(n_63308), .D(n_7540), .SD(1'b1), .Q(code_data
		[84]));
	notech_mux2 i_6066(.S(n_55668), .A(code_data[84]), .B(axi_R[20]), .Z(n_7540
		));
	notech_ao4 i_1263(.A(n_2239), .B(n_8486), .C(n_2237), .D(n_8518), .Z(n_2277
		));
	notech_reg_set code_data_reg_85(.CP(n_63308), .D(n_7546), .SD(1'b1), .Q(code_data
		[85]));
	notech_mux2 i_6074(.S(n_55668), .A(code_data[85]), .B(axi_R[21]), .Z(n_7546
		));
	notech_ao4 i_1262(.A(n_62799), .B(n_8346), .C(n_2244), .D(n_8454), .Z(n_2278
		));
	notech_reg_set code_data_reg_86(.CP(n_63308), .D(n_7552), .SD(1'b1), .Q(code_data
		[86]));
	notech_mux2 i_6082(.S(n_55668), .A(code_data[86]), .B(axi_R[22]), .Z(n_7552
		));
	notech_reg_set code_data_reg_87(.CP(n_63308), .D(n_7558), .SD(1'b1), .Q(code_data
		[87]));
	notech_mux2 i_6090(.S(n_55668), .A(code_data[87]), .B(axi_R[23]), .Z(n_7558
		));
	notech_ao4 i_1272(.A(n_2239), .B(n_8487), .C(n_2237), .D(n_8519), .Z(n_2280
		));
	notech_reg_set code_data_reg_88(.CP(n_63308), .D(n_7564), .SD(1'b1), .Q(code_data
		[88]));
	notech_mux2 i_6098(.S(n_55668), .A(code_data[88]), .B(axi_R[24]), .Z(n_7564
		));
	notech_ao4 i_1271(.A(n_62799), .B(n_8347), .C(n_2244), .D(n_8455), .Z(n_2281
		));
	notech_reg_set code_data_reg_89(.CP(n_63308), .D(n_7570), .SD(1'b1), .Q(code_data
		[89]));
	notech_mux2 i_6106(.S(n_55668), .A(code_data[89]), .B(axi_R[25]), .Z(n_7570
		));
	notech_reg_set code_data_reg_90(.CP(n_63308), .D(n_7576), .SD(1'b1), .Q(code_data
		[90]));
	notech_mux2 i_6114(.S(n_55668), .A(code_data[90]), .B(axi_R[26]), .Z(n_7576
		));
	notech_ao4 i_1281(.A(n_2239), .B(n_8488), .C(n_2237), .D(n_8520), .Z(n_2283
		));
	notech_reg_set code_data_reg_91(.CP(n_63308), .D(n_7582), .SD(1'b1), .Q(code_data
		[91]));
	notech_mux2 i_6122(.S(n_55668), .A(code_data[91]), .B(axi_R[27]), .Z(n_7582
		));
	notech_ao4 i_1280(.A(n_62799), .B(n_8348), .C(n_2244), .D(n_8456), .Z(n_2284
		));
	notech_reg_set code_data_reg_92(.CP(n_63308), .D(n_7588), .SD(1'b1), .Q(code_data
		[92]));
	notech_mux2 i_6130(.S(n_55668), .A(code_data[92]), .B(axi_R[28]), .Z(n_7588
		));
	notech_reg_set code_data_reg_93(.CP(n_63308), .D(n_7594), .SD(1'b1), .Q(code_data
		[93]));
	notech_mux2 i_6138(.S(n_55668), .A(code_data[93]), .B(axi_R[29]), .Z(n_7594
		));
	notech_ao4 i_1290(.A(n_2239), .B(n_8489), .C(n_2237), .D(n_8521), .Z(n_2286
		));
	notech_reg_set code_data_reg_94(.CP(n_63308), .D(n_7600), .SD(1'b1), .Q(code_data
		[94]));
	notech_mux2 i_6146(.S(n_55668), .A(code_data[94]), .B(axi_R[30]), .Z(n_7600
		));
	notech_ao4 i_1289(.A(n_62804), .B(n_8349), .C(n_2244), .D(n_8457), .Z(n_2287
		));
	notech_reg_set code_data_reg_95(.CP(n_63308), .D(n_7606), .SD(1'b1), .Q(code_data
		[95]));
	notech_mux2 i_6154(.S(n_55668), .A(code_data[95]), .B(axi_R[31]), .Z(n_7606
		));
	notech_reg_set code_data_reg_96(.CP(n_63308), .D(n_7612), .SD(1'b1), .Q(code_data
		[96]));
	notech_mux2 i_6162(.S(\nbus_11667[96] ), .A(code_data[96]), .B(axi_R[0])
		, .Z(n_7612));
	notech_ao4 i_1299(.A(n_2239), .B(n_8490), .C(n_2237), .D(n_8522), .Z(n_2289
		));
	notech_reg_set code_data_reg_97(.CP(n_63308), .D(n_7618), .SD(1'b1), .Q(code_data
		[97]));
	notech_mux2 i_6170(.S(\nbus_11667[96] ), .A(code_data[97]), .B(axi_R[1])
		, .Z(n_7618));
	notech_ao4 i_1298(.A(n_62804), .B(n_8350), .C(n_2244), .D(n_8458), .Z(n_2290
		));
	notech_reg_set code_data_reg_98(.CP(n_63308), .D(n_7624), .SD(1'b1), .Q(code_data
		[98]));
	notech_mux2 i_6178(.S(\nbus_11667[96] ), .A(code_data[98]), .B(axi_R[2])
		, .Z(n_7624));
	notech_reg_set code_data_reg_99(.CP(n_63308), .D(n_7630), .SD(1'b1), .Q(code_data
		[99]));
	notech_mux2 i_6186(.S(\nbus_11667[96] ), .A(code_data[99]), .B(axi_R[3])
		, .Z(n_7630));
	notech_ao4 i_1308(.A(n_55475), .B(n_8491), .C(n_55422), .D(n_8523), .Z(n_2292
		));
	notech_reg_set code_data_reg_100(.CP(n_63308), .D(n_7636), .SD(1'b1), .Q
		(code_data[100]));
	notech_mux2 i_6194(.S(\nbus_11667[96] ), .A(code_data[100]), .B(axi_R[4]
		), .Z(n_7636));
	notech_ao4 i_1307(.A(n_62804), .B(n_8351), .C(n_55486), .D(n_8459), .Z(n_2293
		));
	notech_reg_set code_data_reg_101(.CP(n_63308), .D(n_7642), .SD(1'b1), .Q
		(code_data[101]));
	notech_mux2 i_6202(.S(\nbus_11667[96] ), .A(code_data[101]), .B(axi_R[5]
		), .Z(n_7642));
	notech_reg_set code_data_reg_102(.CP(n_63330), .D(n_7648), .SD(1'b1), .Q
		(code_data[102]));
	notech_mux2 i_6210(.S(\nbus_11667[96] ), .A(code_data[102]), .B(axi_R[6]
		), .Z(n_7648));
	notech_ao4 i_1317(.A(n_55475), .B(n_8492), .C(n_55422), .D(n_8524), .Z(n_2295
		));
	notech_reg_set code_data_reg_103(.CP(n_63306), .D(n_7654), .SD(1'b1), .Q
		(code_data[103]));
	notech_mux2 i_6218(.S(\nbus_11667[96] ), .A(code_data[103]), .B(axi_R[7]
		), .Z(n_7654));
	notech_ao4 i_1316(.A(n_62804), .B(n_8352), .C(n_55486), .D(n_8460), .Z(n_2296
		));
	notech_reg_set code_data_reg_104(.CP(n_63330), .D(n_7660), .SD(1'b1), .Q
		(code_data[104]));
	notech_mux2 i_6226(.S(\nbus_11667[96] ), .A(code_data[104]), .B(axi_R[8]
		), .Z(n_7660));
	notech_reg_set code_data_reg_105(.CP(n_63330), .D(n_7666), .SD(1'b1), .Q
		(code_data[105]));
	notech_mux2 i_6234(.S(\nbus_11667[96] ), .A(code_data[105]), .B(axi_R[9]
		), .Z(n_7666));
	notech_ao4 i_1326(.A(n_55475), .B(n_8493), .C(n_55422), .D(n_8525), .Z(n_2298
		));
	notech_reg_set code_data_reg_106(.CP(n_63330), .D(n_7672), .SD(1'b1), .Q
		(code_data[106]));
	notech_mux2 i_6242(.S(\nbus_11667[96] ), .A(code_data[106]), .B(axi_R[10
		]), .Z(n_7672));
	notech_ao4 i_1325(.A(n_62804), .B(n_8353), .C(n_55486), .D(n_8461), .Z(n_2299
		));
	notech_reg_set code_data_reg_107(.CP(n_63330), .D(n_7678), .SD(1'b1), .Q
		(code_data[107]));
	notech_mux2 i_6250(.S(\nbus_11667[96] ), .A(code_data[107]), .B(axi_R[11
		]), .Z(n_7678));
	notech_reg_set code_data_reg_108(.CP(n_63330), .D(n_7684), .SD(1'b1), .Q
		(code_data[108]));
	notech_mux2 i_6258(.S(\nbus_11667[96] ), .A(code_data[108]), .B(axi_R[12
		]), .Z(n_7684));
	notech_ao4 i_1335(.A(n_55475), .B(n_8494), .C(n_55422), .D(n_8526), .Z(n_2301
		));
	notech_reg_set code_data_reg_109(.CP(n_63330), .D(n_7690), .SD(1'b1), .Q
		(code_data[109]));
	notech_mux2 i_6266(.S(\nbus_11667[96] ), .A(code_data[109]), .B(axi_R[13
		]), .Z(n_7690));
	notech_ao4 i_1334(.A(n_62804), .B(n_8354), .C(n_55486), .D(n_8462), .Z(n_2302
		));
	notech_reg_set code_data_reg_110(.CP(n_63330), .D(n_7696), .SD(1'b1), .Q
		(code_data[110]));
	notech_mux2 i_6274(.S(\nbus_11667[96] ), .A(code_data[110]), .B(axi_R[14
		]), .Z(n_7696));
	notech_reg_set code_data_reg_111(.CP(n_63330), .D(n_7702), .SD(1'b1), .Q
		(code_data[111]));
	notech_mux2 i_6282(.S(\nbus_11667[96] ), .A(code_data[111]), .B(axi_R[15
		]), .Z(n_7702));
	notech_ao4 i_1344(.A(n_55475), .B(n_8495), .C(n_55422), .D(n_8527), .Z(n_2304
		));
	notech_reg_set code_data_reg_112(.CP(n_63330), .D(n_7708), .SD(1'b1), .Q
		(code_data[112]));
	notech_mux2 i_6290(.S(n_55690), .A(code_data[112]), .B(axi_R[16]), .Z(n_7708
		));
	notech_ao4 i_1343(.A(n_62809), .B(n_8355), .C(n_55486), .D(n_8463), .Z(n_2305
		));
	notech_reg_set code_data_reg_113(.CP(n_63330), .D(n_7714), .SD(1'b1), .Q
		(code_data[113]));
	notech_mux2 i_6298(.S(n_55690), .A(code_data[113]), .B(axi_R[17]), .Z(n_7714
		));
	notech_reg_set code_data_reg_114(.CP(n_63330), .D(n_7720), .SD(1'b1), .Q
		(code_data[114]));
	notech_mux2 i_6306(.S(n_55690), .A(code_data[114]), .B(axi_R[18]), .Z(n_7720
		));
	notech_ao4 i_1353(.A(n_55475), .B(n_8496), .C(n_55422), .D(n_8528), .Z(n_2307
		));
	notech_reg_set code_data_reg_115(.CP(n_63330), .D(n_7726), .SD(1'b1), .Q
		(code_data[115]));
	notech_mux2 i_6314(.S(n_55690), .A(code_data[115]), .B(axi_R[19]), .Z(n_7726
		));
	notech_ao4 i_1352(.A(n_62804), .B(n_8356), .C(n_55486), .D(n_8464), .Z(n_2308
		));
	notech_reg_set code_data_reg_116(.CP(n_63330), .D(n_7732), .SD(1'b1), .Q
		(code_data[116]));
	notech_mux2 i_6322(.S(n_55690), .A(code_data[116]), .B(axi_R[20]), .Z(n_7732
		));
	notech_reg_set code_data_reg_117(.CP(n_63330), .D(n_7738), .SD(1'b1), .Q
		(code_data[117]));
	notech_mux2 i_6330(.S(n_55690), .A(code_data[117]), .B(axi_R[21]), .Z(n_7738
		));
	notech_ao4 i_1362(.A(n_55475), .B(n_8497), .C(n_55422), .D(n_8529), .Z(n_2310
		));
	notech_reg_set code_data_reg_118(.CP(n_63330), .D(n_7744), .SD(1'b1), .Q
		(code_data[118]));
	notech_mux2 i_6338(.S(n_55690), .A(code_data[118]), .B(axi_R[22]), .Z(n_7744
		));
	notech_ao4 i_1361(.A(n_62804), .B(n_8357), .C(n_55486), .D(n_8465), .Z(n_2311
		));
	notech_reg_set code_data_reg_119(.CP(n_63330), .D(n_7750), .SD(1'b1), .Q
		(code_data[119]));
	notech_mux2 i_6346(.S(n_55690), .A(code_data[119]), .B(axi_R[23]), .Z(n_7750
		));
	notech_reg_set code_data_reg_120(.CP(n_63330), .D(n_7756), .SD(1'b1), .Q
		(code_data[120]));
	notech_mux2 i_6354(.S(n_55690), .A(code_data[120]), .B(axi_R[24]), .Z(n_7756
		));
	notech_ao4 i_1371(.A(n_55475), .B(n_8498), .C(n_55422), .D(n_8530), .Z(n_2313
		));
	notech_reg_set code_data_reg_121(.CP(n_63330), .D(n_7762), .SD(1'b1), .Q
		(code_data[121]));
	notech_mux2 i_6362(.S(n_55690), .A(code_data[121]), .B(axi_R[25]), .Z(n_7762
		));
	notech_ao4 i_1370(.A(n_62804), .B(n_8358), .C(n_55486), .D(n_8466), .Z(n_2314
		));
	notech_reg_set code_data_reg_122(.CP(n_63306), .D(n_7768), .SD(1'b1), .Q
		(code_data[122]));
	notech_mux2 i_6370(.S(n_55690), .A(code_data[122]), .B(axi_R[26]), .Z(n_7768
		));
	notech_reg_set code_data_reg_123(.CP(n_63306), .D(n_7774), .SD(1'b1), .Q
		(code_data[123]));
	notech_mux2 i_6378(.S(n_55690), .A(code_data[123]), .B(axi_R[27]), .Z(n_7774
		));
	notech_ao4 i_1380(.A(n_55475), .B(n_8499), .C(n_55422), .D(n_8531), .Z(n_2316
		));
	notech_reg_set code_data_reg_124(.CP(n_63306), .D(n_7780), .SD(1'b1), .Q
		(code_data[124]));
	notech_mux2 i_6386(.S(n_55690), .A(code_data[124]), .B(axi_R[28]), .Z(n_7780
		));
	notech_ao4 i_1379(.A(n_62804), .B(n_8359), .C(n_55486), .D(n_8467), .Z(n_2317
		));
	notech_reg_set code_data_reg_125(.CP(n_63306), .D(n_7786), .SD(1'b1), .Q
		(code_data[125]));
	notech_mux2 i_6394(.S(n_55690), .A(code_data[125]), .B(axi_R[29]), .Z(n_7786
		));
	notech_reg_set code_data_reg_126(.CP(n_63306), .D(n_7792), .SD(1'b1), .Q
		(code_data[126]));
	notech_mux2 i_6402(.S(n_55690), .A(code_data[126]), .B(axi_R[30]), .Z(n_7792
		));
	notech_ao4 i_1389(.A(n_55475), .B(n_8500), .C(n_55422), .D(n_8532), .Z(n_2319
		));
	notech_reg_set code_data_reg_127(.CP(n_63306), .D(n_7798), .SD(1'b1), .Q
		(code_data[127]));
	notech_mux2 i_6410(.S(n_55690), .A(code_data[127]), .B(axi_R[31]), .Z(n_7798
		));
	notech_ao4 i_1388(.A(n_62804), .B(n_8360), .C(n_55486), .D(n_8468), .Z(n_2320
		));
	notech_reg axi_io_WLAST_reg(.CP(n_63306), .D(n_7804), .CD(n_62713), .Q(axi_io_WLAST
		));
	notech_mux2 i_6418(.S(n_1763), .A(n_23624), .B(axi_io_WLAST), .Z(n_7804)
		);
	notech_reg axi_WVALID_reg(.CP(n_63306), .D(n_7810), .CD(n_62713), .Q(axi_WVALID
		));
	notech_mux2 i_6426(.S(n_1218), .A(n_1176), .B(axi_WVALID), .Z(n_7810));
	notech_ao4 i_1398(.A(n_55475), .B(n_8501), .C(n_2237), .D(n_8533), .Z(n_2322
		));
	notech_reg_set axi_ARBURST_reg_0(.CP(n_63306), .D(n_7816), .SD(n_62713),
		 .Q(axi_ARBURST[0]));
	notech_or2 i_6434(.A(axi_ARBURST[0]), .B(n_8224), .Z(n_7816));
	notech_ao4 i_1397(.A(n_62804), .B(n_8361), .C(n_2244), .D(n_8469), .Z(n_2323
		));
	notech_reg axi_ARBURST_reg_1(.CP(n_63306), .D(n_7825), .CD(n_62713), .Q(axi_ARBURST
		[1]));
	notech_and2 i_6444(.A(axi_ARBURST[1]), .B(n_62788), .Z(n_7825));
	notech_reg axi_io_AW_reg_0(.CP(n_63286), .D(n_7831), .CD(n_62720), .Q(axi_io_AW
		[0]));
	notech_and2 i_6452(.A(n_8334), .B(axi_io_AW[0]), .Z(n_7831));
	notech_ao4 i_1407(.A(n_55475), .B(n_8502), .C(n_55422), .D(n_8534), .Z(n_2325
		));
	notech_reg axi_io_AW_reg_1(.CP(n_63286), .D(n_7837), .CD(n_62720), .Q(axi_io_AW
		[1]));
	notech_and2 i_6460(.A(n_8334), .B(axi_io_AW[1]), .Z(n_7837));
	notech_ao4 i_1406(.A(n_62804), .B(n_8362), .C(n_55486), .D(n_8470), .Z(n_2326
		));
	notech_reg axi_io_AW_reg_2(.CP(n_63310), .D(n_7840), .CD(n_62720), .Q(axi_io_AW
		[2]));
	notech_mux2 i_6466(.S(\nbus_11662[0] ), .A(axi_io_AW[2]), .B(io_add[0]),
		 .Z(n_7840));
	notech_reg axi_io_AW_reg_3(.CP(n_63288), .D(n_7846), .CD(n_62720), .Q(axi_io_AW
		[3]));
	notech_mux2 i_6474(.S(\nbus_11662[0] ), .A(axi_io_AW[3]), .B(io_add[1]),
		 .Z(n_7846));
	notech_ao4 i_1416(.A(n_55475), .B(n_8503), .C(n_55422), .D(n_8535), .Z(n_2328
		));
	notech_reg axi_io_AW_reg_4(.CP(n_63288), .D(n_7852), .CD(n_62720), .Q(axi_io_AW
		[4]));
	notech_mux2 i_6482(.S(\nbus_11662[0] ), .A(axi_io_AW[4]), .B(io_add[2]),
		 .Z(n_7852));
	notech_ao4 i_1415(.A(n_62804), .B(n_8363), .C(n_55486), .D(n_8471), .Z(n_2329
		));
	notech_reg axi_io_AW_reg_5(.CP(n_63288), .D(n_7858), .CD(n_62720), .Q(axi_io_AW
		[5]));
	notech_mux2 i_6490(.S(\nbus_11662[0] ), .A(axi_io_AW[5]), .B(io_add[3]),
		 .Z(n_7858));
	notech_reg axi_io_AW_reg_6(.CP(n_63288), .D(n_7864), .CD(n_62720), .Q(axi_io_AW
		[6]));
	notech_mux2 i_6498(.S(\nbus_11662[0] ), .A(axi_io_AW[6]), .B(io_add[4]),
		 .Z(n_7864));
	notech_ao4 i_1425(.A(n_55475), .B(n_8504), .C(n_55422), .D(n_8536), .Z(n_2331
		));
	notech_reg axi_io_AW_reg_7(.CP(n_63288), .D(n_7870), .CD(n_62720), .Q(axi_io_AW
		[7]));
	notech_mux2 i_6506(.S(\nbus_11662[0] ), .A(axi_io_AW[7]), .B(io_add[5]),
		 .Z(n_7870));
	notech_ao4 i_1424(.A(n_62804), .B(n_8364), .C(n_55486), .D(n_8472), .Z(n_2332
		));
	notech_reg axi_io_AW_reg_8(.CP(n_63288), .D(n_7876), .CD(n_62720), .Q(axi_io_AW
		[8]));
	notech_mux2 i_6514(.S(n_62105), .A(axi_io_AW[8]), .B(io_add[6]), .Z(n_7876
		));
	notech_reg axi_io_AW_reg_9(.CP(n_63288), .D(n_7882), .CD(n_62720), .Q(axi_io_AW
		[9]));
	notech_mux2 i_6522(.S(n_62105), .A(axi_io_AW[9]), .B(io_add[7]), .Z(n_7882
		));
	notech_ao4 i_1434(.A(n_55475), .B(n_8505), .C(n_55422), .D(n_8537), .Z(n_2334
		));
	notech_reg axi_io_AW_reg_10(.CP(n_63288), .D(n_7888), .CD(n_62719), .Q(axi_io_AW
		[10]));
	notech_mux2 i_6530(.S(n_62105), .A(axi_io_AW[10]), .B(io_add[8]), .Z(n_7888
		));
	notech_ao4 i_1433(.A(n_62804), .B(n_8365), .C(n_55486), .D(n_8473), .Z(n_2335
		));
	notech_reg axi_io_AW_reg_11(.CP(n_63288), .D(n_7894), .CD(n_62719), .Q(axi_io_AW
		[11]));
	notech_mux2 i_6538(.S(n_62105), .A(axi_io_AW[11]), .B(io_add[9]), .Z(n_7894
		));
	notech_reg axi_io_AW_reg_12(.CP(n_63288), .D(n_7900), .CD(n_62720), .Q(axi_io_AW
		[12]));
	notech_mux2 i_6546(.S(n_62105), .A(axi_io_AW[12]), .B(io_add[10]), .Z(n_7900
		));
	notech_ao4 i_1443(.A(n_55475), .B(n_8506), .C(n_55422), .D(n_8538), .Z(n_2337
		));
	notech_reg axi_io_AW_reg_13(.CP(n_63310), .D(n_7906), .CD(n_62720), .Q(axi_io_AW
		[13]));
	notech_mux2 i_6554(.S(n_62105), .A(axi_io_AW[13]), .B(io_add[11]), .Z(n_7906
		));
	notech_ao4 i_1442(.A(n_62804), .B(n_8366), .C(n_55486), .D(n_8474), .Z(n_2338
		));
	notech_reg axi_io_AW_reg_14(.CP(n_63310), .D(n_7912), .CD(n_62720), .Q(axi_io_AW
		[14]));
	notech_mux2 i_6562(.S(\nbus_11662[0] ), .A(axi_io_AW[14]), .B(io_add[12]
		), .Z(n_7912));
	notech_reg axi_io_AW_reg_15(.CP(n_63310), .D(n_7918), .CD(n_62720), .Q(axi_io_AW
		[15]));
	notech_mux2 i_6570(.S(\nbus_11662[0] ), .A(axi_io_AW[15]), .B(io_add[13]
		), .Z(n_7918));
	notech_and2 i_1098(.A(n_62720), .B(n_963), .Z(\nbus_11672[0] ));
	notech_reg axi_io_AW_reg_16(.CP(n_63310), .D(n_7924), .CD(n_62721), .Q(axi_io_AW
		[16]));
	notech_mux2 i_6578(.S(\nbus_11662[0] ), .A(axi_io_AW[16]), .B(io_add[14]
		), .Z(n_7924));
	notech_nor2 i_900(.A(n_223056488), .B(n_223356491), .Z(\nbus_11673[0] )
		);
	notech_reg axi_io_AW_reg_17(.CP(n_63310), .D(n_7930), .CD(n_62721), .Q(axi_io_AW
		[17]));
	notech_mux2 i_6586(.S(\nbus_11662[0] ), .A(axi_io_AW[17]), .B(io_add[15]
		), .Z(n_7930));
	notech_nor2 i_899(.A(n_223156489), .B(n_223056488), .Z(\nbus_11662[0] )
		);
	notech_reg axi_io_AW_reg_18(.CP(n_63310), .D(n_7939), .CD(n_62721), .Q(axi_io_AW
		[18]));
	notech_and2 i_6596(.A(axi_io_AW[18]), .B(n_8334), .Z(n_7939));
	notech_and4 i_898(.A(axi_io_RREADY), .B(axi_io_RVALID), .C(n_222856486),
		 .D(n_62721), .Z(\nbus_11671[0] ));
	notech_reg axi_io_AW_reg_19(.CP(n_63310), .D(n_7945), .CD(n_62722), .Q(axi_io_AW
		[19]));
	notech_and2 i_6604(.A(axi_io_AW[19]), .B(n_8334), .Z(n_7945));
	notech_and4 i_896(.A(burst_idx[0]), .B(burst_idx[1]), .C(n_22714), .D(n_210756365
		), .Z(\nbus_11667[96] ));
	notech_reg axi_io_AW_reg_20(.CP(n_63310), .D(n_7951), .CD(n_62722), .Q(axi_io_AW
		[20]));
	notech_and2 i_6612(.A(axi_io_AW[20]), .B(n_8334), .Z(n_7951));
	notech_and3 i_894(.A(n_210756365), .B(n_22714), .C(n_2028), .Z(\nbus_11667[64] 
		));
	notech_reg axi_io_AW_reg_21(.CP(n_63310), .D(n_7957), .CD(n_62721), .Q(axi_io_AW
		[21]));
	notech_and2 i_6620(.A(axi_io_AW[21]), .B(n_8334), .Z(n_7957));
	notech_and3 i_893(.A(n_210756365), .B(n_22714), .C(n_2029), .Z(\nbus_11667[32] 
		));
	notech_reg axi_io_AW_reg_22(.CP(n_63310), .D(n_7963), .CD(n_62721), .Q(axi_io_AW
		[22]));
	notech_and2 i_6628(.A(axi_io_AW[22]), .B(n_8334), .Z(n_7963));
	notech_ao3 i_891(.A(n_210756365), .B(n_22714), .C(n_2036), .Z(\nbus_11667[0] 
		));
	notech_reg axi_io_AW_reg_23(.CP(n_63310), .D(n_7969), .CD(n_62721), .Q(axi_io_AW
		[23]));
	notech_and2 i_6636(.A(axi_io_AW[23]), .B(n_8334), .Z(n_7969));
	notech_ao3 i_26(.A(n_8217), .B(n_2003), .C(busy), .Z(n_23557));
	notech_reg axi_io_AW_reg_24(.CP(n_63310), .D(n_7975), .CD(n_62721), .Q(axi_io_AW
		[24]));
	notech_and2 i_6644(.A(axi_io_AW[24]), .B(n_8334), .Z(n_7975));
	notech_and2 i_211(.A(axi_io_AWVALID), .B(axi_io_AWREADY), .Z(n_23624));
	notech_reg axi_io_AW_reg_25(.CP(n_63310), .D(n_7981), .CD(n_62721), .Q(axi_io_AW
		[25]));
	notech_and2 i_6652(.A(axi_io_AW[25]), .B(n_8334), .Z(n_7981));
	notech_and2 i_29(.A(axi_io_ARVALID), .B(axi_io_ARREADY), .Z(n_23569));
	notech_reg axi_io_AW_reg_26(.CP(n_63310), .D(n_7987), .CD(n_62721), .Q(axi_io_AW
		[26]));
	notech_and2 i_6660(.A(axi_io_AW[26]), .B(n_8334), .Z(n_7987));
	notech_ao3 i_918(.A(n_2003), .B(write_msk[1]), .C(n_2002), .Z(n_25326)
		);
	notech_reg axi_io_AW_reg_27(.CP(n_63310), .D(n_7993), .CD(n_62721), .Q(axi_io_AW
		[27]));
	notech_and2 i_6668(.A(axi_io_AW[27]), .B(n_8334), .Z(n_7993));
	notech_ao3 i_919(.A(n_2003), .B(write_msk[2]), .C(n_2002), .Z(n_25332)
		);
	notech_reg axi_io_AW_reg_28(.CP(n_63310), .D(n_7999), .CD(n_62721), .Q(axi_io_AW
		[28]));
	notech_and2 i_6676(.A(axi_io_AW[28]), .B(n_8334), .Z(n_7999));
	notech_ao3 i_920(.A(n_2003), .B(write_msk[3]), .C(n_2002), .Z(n_25338)
		);
	notech_reg axi_io_AW_reg_29(.CP(n_63310), .D(n_8005), .CD(n_62721), .Q(axi_io_AW
		[29]));
	notech_and2 i_6684(.A(axi_io_AW[29]), .B(n_8334), .Z(n_8005));
	notech_ao3 i_1053(.A(n_62170), .B(cacheQ[146]), .C(n_21466), .Z(n_23512)
		);
	notech_reg axi_io_AW_reg_30(.CP(n_63310), .D(n_8011), .CD(n_62721), .Q(axi_io_AW
		[30]));
	notech_and2 i_6692(.A(axi_io_AW[30]), .B(n_8334), .Z(n_8011));
	notech_ao3 i_1054(.A(n_62170), .B(cacheQ[147]), .C(n_21466), .Z(n_23517)
		);
	notech_reg axi_io_AW_reg_31(.CP(n_63288), .D(n_8017), .CD(n_62719), .Q(axi_io_AW
		[31]));
	notech_and2 i_6700(.A(axi_io_AW[31]), .B(n_8334), .Z(n_8017));
	notech_ao3 i_1055(.A(n_62170), .B(cacheQ[149]), .C(n_21466), .Z(n_23527)
		);
	notech_reg axi_io_W_reg_0(.CP(n_63288), .D(n_8020), .CD(n_62717), .Q(axi_io_W
		[0]));
	notech_mux2 i_6706(.S(\nbus_11662[0] ), .A(axi_io_W[0]), .B(writeio_data
		[0]), .Z(n_8020));
	notech_and4 i_56126(.A(fsm[4]), .B(fsm[0]), .C(n_1999), .D(n_8328), .Z(n_22714
		));
	notech_reg axi_io_W_reg_1(.CP(n_63290), .D(n_8026), .CD(n_62717), .Q(axi_io_W
		[1]));
	notech_mux2 i_6714(.S(\nbus_11662[0] ), .A(axi_io_W[1]), .B(writeio_data
		[1]), .Z(n_8026));
	notech_and2 i_1074(.A(write_data[8]), .B(n_8233), .Z(n_24828));
	notech_reg axi_io_W_reg_2(.CP(n_63290), .D(n_8032), .CD(n_62717), .Q(axi_io_W
		[2]));
	notech_mux2 i_6722(.S(\nbus_11662[0] ), .A(axi_io_W[2]), .B(writeio_data
		[2]), .Z(n_8032));
	notech_and2 i_1075(.A(write_data[9]), .B(n_8233), .Z(n_24834));
	notech_reg axi_io_W_reg_3(.CP(n_63290), .D(n_8038), .CD(n_62717), .Q(axi_io_W
		[3]));
	notech_mux2 i_6730(.S(\nbus_11662[0] ), .A(axi_io_W[3]), .B(writeio_data
		[3]), .Z(n_8038));
	notech_and2 i_1076(.A(write_data[10]), .B(n_8233), .Z(n_24840));
	notech_reg axi_io_W_reg_4(.CP(n_63290), .D(n_8044), .CD(n_62717), .Q(axi_io_W
		[4]));
	notech_mux2 i_6738(.S(\nbus_11662[0] ), .A(axi_io_W[4]), .B(writeio_data
		[4]), .Z(n_8044));
	notech_and2 i_1077(.A(write_data[11]), .B(n_8233), .Z(n_24846));
	notech_reg axi_io_W_reg_5(.CP(n_63290), .D(n_8050), .CD(n_62717), .Q(axi_io_W
		[5]));
	notech_mux2 i_6746(.S(\nbus_11662[0] ), .A(axi_io_W[5]), .B(writeio_data
		[5]), .Z(n_8050));
	notech_and2 i_1078(.A(write_data[12]), .B(n_8233), .Z(n_24852));
	notech_reg axi_io_W_reg_6(.CP(n_63290), .D(n_8056), .CD(n_62717), .Q(axi_io_W
		[6]));
	notech_mux2 i_6754(.S(\nbus_11662[0] ), .A(axi_io_W[6]), .B(writeio_data
		[6]), .Z(n_8056));
	notech_and2 i_1079(.A(write_data[13]), .B(n_8233), .Z(n_24858));
	notech_reg axi_io_W_reg_7(.CP(n_63290), .D(n_8062), .CD(n_62717), .Q(axi_io_W
		[7]));
	notech_mux2 i_6762(.S(\nbus_11662[0] ), .A(axi_io_W[7]), .B(writeio_data
		[7]), .Z(n_8062));
	notech_and2 i_1080(.A(write_data[14]), .B(n_8233), .Z(n_24864));
	notech_reg axi_io_W_reg_8(.CP(n_63290), .D(n_8068), .CD(n_62716), .Q(axi_io_W
		[8]));
	notech_mux2 i_6770(.S(n_62105), .A(axi_io_W[8]), .B(writeio_data[8]), .Z
		(n_8068));
	notech_and2 i_1081(.A(write_data[15]), .B(n_8233), .Z(n_24870));
	notech_reg axi_io_W_reg_9(.CP(n_63290), .D(n_8074), .CD(n_62716), .Q(axi_io_W
		[9]));
	notech_mux2 i_6778(.S(n_62101), .A(axi_io_W[9]), .B(writeio_data[9]), .Z
		(n_8074));
	notech_and2 i_1082(.A(write_data[16]), .B(n_8233), .Z(n_24876));
	notech_reg axi_io_W_reg_10(.CP(n_63290), .D(n_8080), .CD(n_62716), .Q(axi_io_W
		[10]));
	notech_mux2 i_6786(.S(n_62101), .A(axi_io_W[10]), .B(writeio_data[10]), 
		.Z(n_8080));
	notech_and2 i_1083(.A(write_data[17]), .B(n_8233), .Z(n_24882));
	notech_reg axi_io_W_reg_11(.CP(n_63290), .D(n_8086), .CD(n_62716), .Q(axi_io_W
		[11]));
	notech_mux2 i_6794(.S(n_62101), .A(axi_io_W[11]), .B(writeio_data[11]), 
		.Z(n_8086));
	notech_and2 i_1084(.A(write_data[18]), .B(n_8233), .Z(n_24888));
	notech_reg axi_io_W_reg_12(.CP(n_63290), .D(n_8092), .CD(n_62716), .Q(axi_io_W
		[12]));
	notech_mux2 i_6802(.S(n_62101), .A(axi_io_W[12]), .B(writeio_data[12]), 
		.Z(n_8092));
	notech_and2 i_1085(.A(write_data[19]), .B(n_8233), .Z(n_24894));
	notech_reg axi_io_W_reg_13(.CP(n_63290), .D(n_8098), .CD(n_62717), .Q(axi_io_W
		[13]));
	notech_mux2 i_6810(.S(n_62101), .A(axi_io_W[13]), .B(writeio_data[13]), 
		.Z(n_8098));
	notech_and2 i_1086(.A(write_data[20]), .B(n_62114), .Z(n_24900));
	notech_reg axi_io_W_reg_14(.CP(n_63290), .D(n_8104), .CD(n_62716), .Q(axi_io_W
		[14]));
	notech_mux2 i_6818(.S(n_62101), .A(axi_io_W[14]), .B(writeio_data[14]), 
		.Z(n_8104));
	notech_and2 i_1087(.A(write_data[21]), .B(n_62114), .Z(n_24906));
	notech_reg axi_io_W_reg_15(.CP(n_63290), .D(n_8110), .CD(n_62716), .Q(axi_io_W
		[15]));
	notech_mux2 i_6826(.S(n_62101), .A(axi_io_W[15]), .B(writeio_data[15]), 
		.Z(n_8110));
	notech_and2 i_1088(.A(write_data[22]), .B(n_62114), .Z(n_24912));
	notech_reg axi_io_W_reg_16(.CP(n_63290), .D(n_8116), .CD(n_62717), .Q(axi_io_W
		[16]));
	notech_mux2 i_6834(.S(n_62101), .A(axi_io_W[16]), .B(writeio_data[16]), 
		.Z(n_8116));
	notech_and2 i_1089(.A(write_data[23]), .B(n_62114), .Z(n_24918));
	notech_reg axi_io_W_reg_17(.CP(n_63290), .D(n_8122), .CD(n_62719), .Q(axi_io_W
		[17]));
	notech_mux2 i_6842(.S(n_62101), .A(axi_io_W[17]), .B(writeio_data[17]), 
		.Z(n_8122));
	notech_and2 i_1090(.A(write_data[24]), .B(n_62114), .Z(n_24924));
	notech_reg axi_io_W_reg_18(.CP(n_63290), .D(n_8128), .CD(n_62719), .Q(axi_io_W
		[18]));
	notech_mux2 i_6850(.S(n_62101), .A(axi_io_W[18]), .B(writeio_data[18]), 
		.Z(n_8128));
	notech_and2 i_1091(.A(write_data[25]), .B(n_62114), .Z(n_24930));
	notech_reg axi_io_W_reg_19(.CP(n_63290), .D(n_8134), .CD(n_62719), .Q(axi_io_W
		[19]));
	notech_mux2 i_6858(.S(n_62101), .A(axi_io_W[19]), .B(writeio_data[19]), 
		.Z(n_8134));
	notech_and2 i_1092(.A(write_data[26]), .B(n_62114), .Z(n_24936));
	notech_reg axi_io_W_reg_20(.CP(clk), .D(n_8140), .CD(n_62719), .Q(axi_io_W
		[20]));
	notech_mux2 i_6866(.S(n_62101), .A(axi_io_W[20]), .B(writeio_data[20]), 
		.Z(n_8140));
	notech_and2 i_1093(.A(write_data[27]), .B(n_62114), .Z(n_24942));
	notech_reg axi_io_W_reg_21(.CP(clk), .D(n_8146), .CD(n_62719), .Q(axi_io_W
		[21]));
	notech_mux2 i_6874(.S(n_62105), .A(axi_io_W[21]), .B(writeio_data[21]), 
		.Z(n_8146));
	notech_and2 i_1094(.A(write_data[28]), .B(n_62114), .Z(n_24948));
	notech_reg axi_io_W_reg_22(.CP(clk), .D(n_8152), .CD(n_62719), .Q(axi_io_W
		[22]));
	notech_mux2 i_6882(.S(n_62105), .A(axi_io_W[22]), .B(writeio_data[22]), 
		.Z(n_8152));
	notech_and2 i_1095(.A(write_data[29]), .B(n_62114), .Z(n_24954));
	notech_reg axi_io_W_reg_23(.CP(clk), .D(n_8158), .CD(n_62719), .Q(axi_io_W
		[23]));
	notech_mux2 i_6890(.S(n_62105), .A(axi_io_W[23]), .B(writeio_data[23]), 
		.Z(n_8158));
	notech_and2 i_1096(.A(write_data[30]), .B(n_62114), .Z(n_24960));
	notech_reg axi_io_W_reg_24(.CP(clk), .D(n_8164), .CD(n_62719), .Q(axi_io_W
		[24]));
	notech_mux2 i_6898(.S(n_62105), .A(axi_io_W[24]), .B(writeio_data[24]), 
		.Z(n_8164));
	notech_and2 i_1097(.A(write_data[31]), .B(n_62114), .Z(n_24966));
	notech_reg axi_io_W_reg_25(.CP(clk), .D(n_8170), .CD(n_62717), .Q(axi_io_W
		[25]));
	notech_mux2 i_6906(.S(n_62105), .A(axi_io_W[25]), .B(writeio_data[25]), 
		.Z(n_8170));
	notech_ao4 i_1104(.A(n_2029), .B(n_2028), .C(n_22714), .D(n_62132), .Z(n_25495
		));
	notech_reg axi_io_W_reg_26(.CP(clk), .D(n_8176), .CD(n_62717), .Q(axi_io_W
		[26]));
	notech_mux2 i_6914(.S(n_62105), .A(axi_io_W[26]), .B(writeio_data[26]), 
		.Z(n_8176));
	notech_nor2 i_1105(.A(n_965), .B(n_2024), .Z(n_25500));
	notech_reg axi_io_W_reg_27(.CP(clk), .D(n_8182), .CD(n_62717), .Q(axi_io_W
		[27]));
	notech_mux2 i_6922(.S(n_62101), .A(axi_io_W[27]), .B(writeio_data[27]), 
		.Z(n_8182));
	notech_nor2 i_1106(.A(n_2024), .B(n_966), .Z(n_25505));
	notech_reg axi_io_W_reg_28(.CP(clk), .D(n_8188), .CD(n_62717), .Q(axi_io_W
		[28]));
	notech_mux2 i_6930(.S(n_62101), .A(axi_io_W[28]), .B(writeio_data[28]), 
		.Z(n_8188));
	notech_nor2 i_1107(.A(n_2024), .B(n_967), .Z(n_25510));
	notech_reg axi_io_W_reg_29(.CP(clk), .D(n_8194), .CD(n_62719), .Q(axi_io_W
		[29]));
	notech_mux2 i_6938(.S(n_62101), .A(axi_io_W[29]), .B(writeio_data[29]), 
		.Z(n_8194));
	notech_and4 i_56139(.A(fsm[4]), .B(n_1999), .C(fsm[3]), .D(n_8325), .Z(n_25047
		));
	notech_reg axi_io_W_reg_30(.CP(clk), .D(n_8200), .CD(n_62719), .Q(axi_io_W
		[30]));
	notech_mux2 i_6946(.S(n_62105), .A(axi_io_W[30]), .B(writeio_data[30]), 
		.Z(n_8200));
	notech_reg axi_io_W_reg_31(.CP(clk), .D(n_8206), .CD(n_62717), .Q(axi_io_W
		[31]));
	notech_mux2 i_6954(.S(n_62105), .A(axi_io_W[31]), .B(writeio_data[31]), 
		.Z(n_8206));
	notech_inv i_9031(.A(n_62132), .Z(n_8212));
	notech_inv i_9032(.A(n_2052), .Z(n_8213));
	notech_inv i_9033(.A(n_2016), .Z(n_8214));
	notech_inv i_9034(.A(n_221956477), .Z(n_8215));
	notech_inv i_9035(.A(n_2050), .Z(n_8216));
	notech_inv i_9036(.A(n_970), .Z(n_8217));
	notech_inv i_9037(.A(n_222856486), .Z(n_8218));
	notech_inv i_9038(.A(n_222956487), .Z(n_8219));
	notech_inv i_9039(.A(n_2037), .Z(n_8220));
	notech_inv i_9040(.A(n_2069), .Z(n_8221));
	notech_inv i_9041(.A(n_2029), .Z(n_8222));
	notech_inv i_9042(.A(n_2028), .Z(n_8223));
	notech_inv i_9043(.A(n_62788), .Z(n_8224));
	notech_inv i_9044(.A(n_1742), .Z(n_8225));
	notech_inv i_9045(.A(n_973), .Z(n_8226));
	notech_inv i_9046(.A(n_980), .Z(n_8227));
	notech_inv i_9047(.A(n_983), .Z(n_8228));
	notech_inv i_9048(.A(n_2042), .Z(n_8229));
	notech_inv i_9049(.A(n_986), .Z(n_8230));
	notech_inv i_9050(.A(n_989), .Z(n_8231));
	notech_inv i_9051(.A(n_992), .Z(n_8232));
	notech_inv i_9052(.A(n_62734), .Z(n_8233));
	notech_inv i_9053(.A(n_995), .Z(n_8234));
	notech_inv i_9054(.A(n_998), .Z(n_8235));
	notech_inv i_9055(.A(n_1001), .Z(n_8236));
	notech_inv i_9056(.A(n_1004), .Z(n_8237));
	notech_inv i_9057(.A(n_1007), .Z(n_8238));
	notech_inv i_9058(.A(n_1010), .Z(n_8239));
	notech_inv i_9059(.A(n_1013), .Z(n_8240));
	notech_inv i_9060(.A(n_1016), .Z(n_8241));
	notech_inv i_9061(.A(n_1019), .Z(n_8242));
	notech_inv i_9062(.A(n_1022), .Z(n_8243));
	notech_inv i_9063(.A(n_1025), .Z(n_8244));
	notech_inv i_9064(.A(n_1028), .Z(n_8245));
	notech_inv i_9065(.A(n_1031), .Z(n_8246));
	notech_inv i_9066(.A(n_1034), .Z(n_8247));
	notech_inv i_9067(.A(n_1037), .Z(n_8248));
	notech_inv i_9068(.A(n_1040), .Z(n_8249));
	notech_inv i_9069(.A(n_1043), .Z(n_8250));
	notech_inv i_9070(.A(n_1046), .Z(n_8251));
	notech_inv i_9071(.A(n_1049), .Z(n_8252));
	notech_inv i_9072(.A(n_1052), .Z(n_8253));
	notech_inv i_9073(.A(n_1055), .Z(n_8254));
	notech_inv i_9074(.A(n_1058), .Z(n_8255));
	notech_inv i_9075(.A(n_1062), .Z(n_8256));
	notech_inv i_9076(.A(n_1065), .Z(n_8257));
	notech_inv i_9077(.A(n_1070), .Z(n_8258));
	notech_inv i_9078(.A(n_1073), .Z(n_8259));
	notech_inv i_9079(.A(n_1076), .Z(n_8260));
	notech_inv i_9080(.A(n_1079), .Z(n_8261));
	notech_inv i_9081(.A(n_1082), .Z(n_8262));
	notech_inv i_9082(.A(n_1085), .Z(n_8263));
	notech_inv i_9083(.A(n_1088), .Z(n_8264));
	notech_inv i_9084(.A(n_22714), .Z(n_8265));
	notech_inv i_9085(.A(n_1091), .Z(n_8266));
	notech_inv i_9086(.A(n_1094), .Z(n_8267));
	notech_inv i_9087(.A(n_1097), .Z(n_8268));
	notech_inv i_9088(.A(n_1100), .Z(n_8269));
	notech_inv i_9089(.A(n_1103), .Z(n_8270));
	notech_inv i_9090(.A(n_1106), .Z(n_8271));
	notech_inv i_9091(.A(n_1109), .Z(n_8272));
	notech_inv i_9092(.A(n_1112), .Z(n_8273));
	notech_inv i_9093(.A(n_1115), .Z(n_8274));
	notech_inv i_9094(.A(n_1118), .Z(n_8275));
	notech_inv i_9095(.A(n_1121), .Z(n_8276));
	notech_inv i_9096(.A(n_1124), .Z(n_8277));
	notech_inv i_9097(.A(n_1127), .Z(n_8278));
	notech_inv i_9098(.A(n_1130), .Z(n_8279));
	notech_inv i_9099(.A(n_1133), .Z(n_8280));
	notech_inv i_9100(.A(n_1136), .Z(n_8281));
	notech_inv i_9101(.A(n_1139), .Z(n_8282));
	notech_inv i_9102(.A(n_1142), .Z(n_8283));
	notech_inv i_9103(.A(n_1145), .Z(n_8284));
	notech_inv i_9104(.A(n_1148), .Z(n_8285));
	notech_inv i_9105(.A(n_1151), .Z(n_8286));
	notech_inv i_9106(.A(n_1154), .Z(n_8287));
	notech_inv i_9107(.A(n_1157), .Z(n_8288));
	notech_inv i_9108(.A(n_1160), .Z(n_8289));
	notech_inv i_9109(.A(n_1173), .Z(n_8290));
	notech_inv i_9110(.A(n_1179), .Z(n_8291));
	notech_inv i_9111(.A(n_1182), .Z(n_8292));
	notech_inv i_9112(.A(n_1185), .Z(n_8293));
	notech_inv i_9113(.A(n_1188), .Z(n_8294));
	notech_inv i_9114(.A(n_1191), .Z(n_8295));
	notech_inv i_9115(.A(n_1194), .Z(n_8296));
	notech_inv i_9116(.A(n_1197), .Z(n_8297));
	notech_inv i_9117(.A(n_1200), .Z(n_8298));
	notech_inv i_9118(.A(n_1213), .Z(n_8299));
	notech_inv i_9119(.A(n_1221), .Z(n_8300));
	notech_inv i_9120(.A(n_1223), .Z(n_8301));
	notech_inv i_9121(.A(burst_idx[1]), .Z(n_8302));
	notech_inv i_9122(.A(burst_idx[2]), .Z(n_8303));
	notech_inv i_9123(.A(burst_idx[3]), .Z(n_8304));
	notech_inv i_9124(.A(n_1227), .Z(n_8305));
	notech_inv i_9125(.A(n_1230), .Z(n_8306));
	notech_inv i_9127(.A(n_1233), .Z(n_8308));
	notech_inv i_9128(.A(n_1236), .Z(n_8309));
	notech_inv i_9129(.A(n_1239), .Z(n_8310));
	notech_inv i_9130(.A(n_1242), .Z(n_8311));
	notech_inv i_9131(.A(n_1245), .Z(n_8312));
	notech_inv i_9132(.A(n_1248), .Z(n_8313));
	notech_inv i_9133(.A(n_1251), .Z(n_8314));
	notech_inv i_9134(.A(n_1254), .Z(n_8315));
	notech_inv i_9135(.A(n_1257), .Z(n_8316));
	notech_inv i_9136(.A(n_1260), .Z(n_8317));
	notech_inv i_9137(.A(n_1263), .Z(n_8318));
	notech_inv i_9138(.A(n_1266), .Z(n_8319));
	notech_inv i_9139(.A(n_1269), .Z(n_8320));
	notech_inv i_9140(.A(n_1272), .Z(n_8321));
	notech_inv i_9141(.A(n_1275), .Z(n_8322));
	notech_inv i_9142(.A(n_23557), .Z(n_8323));
	notech_inv i_9143(.A(n_1280), .Z(n_8324));
	notech_inv i_9144(.A(fsm[0]), .Z(n_8325));
	notech_inv i_9145(.A(fsm[1]), .Z(n_8326));
	notech_inv i_9146(.A(fsm[2]), .Z(n_8327));
	notech_inv i_9147(.A(fsm[3]), .Z(n_8328));
	notech_inv i_9148(.A(wf), .Z(n_8329));
	notech_inv i_9149(.A(n_23569), .Z(n_8330));
	notech_inv i_9150(.A(\nbus_11673[0] ), .Z(n_8331));
	notech_inv i_9151(.A(n_1710), .Z(n_8332));
	notech_inv i_9152(.A(n_23624), .Z(n_8333));
	notech_inv i_9153(.A(n_62105), .Z(n_8334));
	notech_inv i_9154(.A(axi_R[0]), .Z(n_8335));
	notech_inv i_9155(.A(axi_R[1]), .Z(n_8336));
	notech_inv i_9156(.A(axi_R[2]), .Z(n_8337));
	notech_inv i_9157(.A(axi_R[3]), .Z(n_8338));
	notech_inv i_9158(.A(axi_R[4]), .Z(n_8339));
	notech_inv i_9159(.A(axi_R[5]), .Z(n_8340));
	notech_inv i_9160(.A(axi_R[6]), .Z(n_8341));
	notech_inv i_9161(.A(axi_R[7]), .Z(n_8342));
	notech_inv i_9162(.A(axi_R[8]), .Z(n_8343));
	notech_inv i_9163(.A(axi_R[9]), .Z(n_8344));
	notech_inv i_9164(.A(axi_R[10]), .Z(n_8345));
	notech_inv i_9165(.A(axi_R[11]), .Z(n_8346));
	notech_inv i_9166(.A(axi_R[12]), .Z(n_8347));
	notech_inv i_9167(.A(axi_R[13]), .Z(n_8348));
	notech_inv i_9168(.A(axi_R[14]), .Z(n_8349));
	notech_inv i_9169(.A(axi_R[15]), .Z(n_8350));
	notech_inv i_9170(.A(axi_R[16]), .Z(n_8351));
	notech_inv i_9171(.A(axi_R[17]), .Z(n_8352));
	notech_inv i_9172(.A(axi_R[18]), .Z(n_8353));
	notech_inv i_9173(.A(axi_R[19]), .Z(n_8354));
	notech_inv i_9174(.A(axi_R[20]), .Z(n_8355));
	notech_inv i_9175(.A(axi_R[21]), .Z(n_8356));
	notech_inv i_9176(.A(axi_R[22]), .Z(n_8357));
	notech_inv i_9177(.A(axi_R[23]), .Z(n_8358));
	notech_inv i_9178(.A(axi_R[24]), .Z(n_8359));
	notech_inv i_9179(.A(axi_R[25]), .Z(n_8360));
	notech_inv i_9180(.A(axi_R[26]), .Z(n_8361));
	notech_inv i_9181(.A(axi_R[27]), .Z(n_8362));
	notech_inv i_9182(.A(axi_R[28]), .Z(n_8363));
	notech_inv i_9183(.A(axi_R[29]), .Z(n_8364));
	notech_inv i_9184(.A(axi_R[30]), .Z(n_8365));
	notech_inv i_9185(.A(axi_R[31]), .Z(n_8366));
	notech_inv i_9186(.A(Daddr[2]), .Z(n_8367));
	notech_inv i_9187(.A(Daddr[3]), .Z(n_8368));
	notech_inv i_9188(.A(Daddr[13]), .Z(n_8369));
	notech_inv i_9189(.A(Daddr[12]), .Z(n_8370));
	notech_inv i_9190(.A(Daddr[11]), .Z(n_8371));
	notech_inv i_9191(.A(Daddr[10]), .Z(n_8372));
	notech_inv i_9192(.A(Daddr[9]), .Z(n_8373));
	notech_inv i_9193(.A(Daddr[8]), .Z(n_8374));
	notech_inv i_9194(.A(Daddr[7]), .Z(n_8375));
	notech_inv i_9195(.A(Daddr[6]), .Z(n_8376));
	notech_inv i_9196(.A(Daddr[5]), .Z(n_8377));
	notech_inv i_9197(.A(Daddr[4]), .Z(n_8378));
	notech_inv i_9198(.A(Daddr[14]), .Z(n_8379));
	notech_inv i_9199(.A(Daddr[15]), .Z(n_8380));
	notech_inv i_9200(.A(Daddr[16]), .Z(n_8381));
	notech_inv i_9201(.A(Daddr[17]), .Z(n_8382));
	notech_inv i_9202(.A(Daddr[18]), .Z(n_8383));
	notech_inv i_9203(.A(Daddr[19]), .Z(n_8384));
	notech_inv i_9204(.A(Daddr[20]), .Z(n_8385));
	notech_inv i_9205(.A(Daddr[21]), .Z(n_8386));
	notech_inv i_9206(.A(Daddr[22]), .Z(n_8387));
	notech_inv i_9207(.A(Daddr[23]), .Z(n_8388));
	notech_inv i_9208(.A(Daddr[24]), .Z(n_8389));
	notech_inv i_9209(.A(Daddr[25]), .Z(n_8390));
	notech_inv i_9210(.A(Daddr[26]), .Z(n_8391));
	notech_inv i_9211(.A(Daddr[27]), .Z(n_8392));
	notech_inv i_9212(.A(Daddr[28]), .Z(n_8393));
	notech_inv i_9213(.A(Daddr[29]), .Z(n_8394));
	notech_inv i_9214(.A(Daddr[30]), .Z(n_8395));
	notech_inv i_9215(.A(Daddr[31]), .Z(n_8396));
	notech_inv i_9216(.A(code_wdata[0]), .Z(n_8397));
	notech_inv i_9217(.A(code_wdata[1]), .Z(n_8398));
	notech_inv i_9218(.A(code_wdata[2]), .Z(n_8399));
	notech_inv i_9219(.A(code_wdata[3]), .Z(n_8400));
	notech_inv i_9220(.A(code_wdata[4]), .Z(n_8401));
	notech_inv i_9221(.A(code_wdata[5]), .Z(n_8402));
	notech_inv i_9222(.A(code_wdata[6]), .Z(n_8403));
	notech_inv i_9223(.A(code_wdata[7]), .Z(n_8404));
	notech_inv i_9224(.A(code_addr[2]), .Z(n_8405));
	notech_inv i_9225(.A(code_addr[3]), .Z(n_8406));
	notech_inv i_9226(.A(code_addr[4]), .Z(n_8407));
	notech_inv i_9227(.A(code_addr[5]), .Z(n_8408));
	notech_inv i_9228(.A(code_addr[6]), .Z(n_8409));
	notech_inv i_9229(.A(code_addr[7]), .Z(n_8410));
	notech_inv i_9230(.A(code_addr[8]), .Z(n_8411));
	notech_inv i_9231(.A(code_addr[9]), .Z(n_8412));
	notech_inv i_9232(.A(code_addr[10]), .Z(n_8413));
	notech_inv i_9233(.A(code_addr[11]), .Z(n_8414));
	notech_inv i_9234(.A(code_addr[12]), .Z(n_8415));
	notech_inv i_9235(.A(code_addr[13]), .Z(n_8416));
	notech_inv i_9236(.A(code_addr[14]), .Z(n_8417));
	notech_inv i_9237(.A(code_addr[15]), .Z(n_8418));
	notech_inv i_9238(.A(code_addr[16]), .Z(n_8419));
	notech_inv i_9239(.A(code_addr[17]), .Z(n_8420));
	notech_inv i_9240(.A(code_addr[18]), .Z(n_8421));
	notech_inv i_9241(.A(code_addr[19]), .Z(n_8422));
	notech_inv i_9242(.A(code_addr[20]), .Z(n_8423));
	notech_inv i_9243(.A(code_addr[21]), .Z(n_8424));
	notech_inv i_9244(.A(code_addr[22]), .Z(n_8425));
	notech_inv i_9245(.A(code_addr[23]), .Z(n_8426));
	notech_inv i_9246(.A(code_addr[24]), .Z(n_8427));
	notech_inv i_9247(.A(code_addr[25]), .Z(n_8428));
	notech_inv i_9248(.A(code_addr[26]), .Z(n_8429));
	notech_inv i_9249(.A(code_addr[27]), .Z(n_8430));
	notech_inv i_9250(.A(code_addr[28]), .Z(n_8431));
	notech_inv i_9251(.A(code_addr[29]), .Z(n_8432));
	notech_inv i_9252(.A(code_addr[30]), .Z(n_8433));
	notech_inv i_9253(.A(code_addr[31]), .Z(n_8434));
	notech_inv i_9254(.A(write_data[0]), .Z(n_8435));
	notech_inv i_9255(.A(write_data[1]), .Z(n_8436));
	notech_inv i_9256(.A(write_data[2]), .Z(n_8437));
	notech_inv i_9257(.A(write_data[3]), .Z(n_8438));
	notech_inv i_9258(.A(write_data[4]), .Z(n_8439));
	notech_inv i_9259(.A(write_data[5]), .Z(n_8440));
	notech_inv i_9260(.A(write_data[6]), .Z(n_8441));
	notech_inv i_9261(.A(write_data[7]), .Z(n_8442));
	notech_inv i_9262(.A(cacheQ[0]), .Z(n_8443));
	notech_inv i_9263(.A(cacheQ[1]), .Z(n_8444));
	notech_inv i_9264(.A(cacheQ[2]), .Z(n_8445));
	notech_inv i_9265(.A(cacheQ[3]), .Z(n_8446));
	notech_inv i_9266(.A(cacheQ[4]), .Z(n_8447));
	notech_inv i_9267(.A(cacheQ[5]), .Z(n_8448));
	notech_inv i_9268(.A(cacheQ[6]), .Z(n_8449));
	notech_inv i_9269(.A(cacheQ[7]), .Z(n_8450));
	notech_inv i_9270(.A(cacheQ[8]), .Z(n_8451));
	notech_inv i_9271(.A(cacheQ[9]), .Z(n_8452));
	notech_inv i_9272(.A(cacheQ[10]), .Z(n_8453));
	notech_inv i_9273(.A(cacheQ[11]), .Z(n_8454));
	notech_inv i_9274(.A(cacheQ[12]), .Z(n_8455));
	notech_inv i_9275(.A(cacheQ[13]), .Z(n_8456));
	notech_inv i_9276(.A(cacheQ[14]), .Z(n_8457));
	notech_inv i_9277(.A(cacheQ[15]), .Z(n_8458));
	notech_inv i_9278(.A(cacheQ[16]), .Z(n_8459));
	notech_inv i_9279(.A(cacheQ[17]), .Z(n_8460));
	notech_inv i_9280(.A(cacheQ[18]), .Z(n_8461));
	notech_inv i_9281(.A(cacheQ[19]), .Z(n_8462));
	notech_inv i_9282(.A(cacheQ[20]), .Z(n_8463));
	notech_inv i_9283(.A(cacheQ[21]), .Z(n_8464));
	notech_inv i_9284(.A(cacheQ[22]), .Z(n_8465));
	notech_inv i_9285(.A(cacheQ[23]), .Z(n_8466));
	notech_inv i_9286(.A(cacheQ[24]), .Z(n_8467));
	notech_inv i_9287(.A(cacheQ[25]), .Z(n_8468));
	notech_inv i_9288(.A(cacheQ[26]), .Z(n_8469));
	notech_inv i_9289(.A(cacheQ[27]), .Z(n_8470));
	notech_inv i_9290(.A(cacheQ[28]), .Z(n_8471));
	notech_inv i_9291(.A(cacheQ[29]), .Z(n_8472));
	notech_inv i_9292(.A(cacheQ[30]), .Z(n_8473));
	notech_inv i_9293(.A(cacheQ[31]), .Z(n_8474));
	notech_inv i_9294(.A(cacheQ[32]), .Z(n_8475));
	notech_inv i_9295(.A(cacheQ[33]), .Z(n_8476));
	notech_inv i_9296(.A(cacheQ[34]), .Z(n_8477));
	notech_inv i_9297(.A(cacheQ[35]), .Z(n_8478));
	notech_inv i_9298(.A(cacheQ[36]), .Z(n_8479));
	notech_inv i_9299(.A(cacheQ[37]), .Z(n_8480));
	notech_inv i_9300(.A(cacheQ[38]), .Z(n_8481));
	notech_inv i_9301(.A(cacheQ[39]), .Z(n_8482));
	notech_inv i_9302(.A(cacheQ[40]), .Z(n_8483));
	notech_inv i_9303(.A(cacheQ[41]), .Z(n_8484));
	notech_inv i_9304(.A(cacheQ[42]), .Z(n_8485));
	notech_inv i_9305(.A(cacheQ[43]), .Z(n_8486));
	notech_inv i_9306(.A(cacheQ[44]), .Z(n_8487));
	notech_inv i_9307(.A(cacheQ[45]), .Z(n_8488));
	notech_inv i_9308(.A(cacheQ[46]), .Z(n_8489));
	notech_inv i_9309(.A(cacheQ[47]), .Z(n_8490));
	notech_inv i_9310(.A(cacheQ[48]), .Z(n_8491));
	notech_inv i_9311(.A(cacheQ[49]), .Z(n_8492));
	notech_inv i_9312(.A(cacheQ[50]), .Z(n_8493));
	notech_inv i_9313(.A(cacheQ[51]), .Z(n_8494));
	notech_inv i_9314(.A(cacheQ[52]), .Z(n_8495));
	notech_inv i_9315(.A(cacheQ[53]), .Z(n_8496));
	notech_inv i_9316(.A(cacheQ[54]), .Z(n_8497));
	notech_inv i_9317(.A(cacheQ[55]), .Z(n_8498));
	notech_inv i_9318(.A(cacheQ[56]), .Z(n_8499));
	notech_inv i_9319(.A(cacheQ[57]), .Z(n_8500));
	notech_inv i_9320(.A(cacheQ[58]), .Z(n_8501));
	notech_inv i_9321(.A(cacheQ[59]), .Z(n_8502));
	notech_inv i_9322(.A(cacheQ[60]), .Z(n_8503));
	notech_inv i_9323(.A(cacheQ[61]), .Z(n_8504));
	notech_inv i_9324(.A(cacheQ[62]), .Z(n_8505));
	notech_inv i_9325(.A(cacheQ[63]), .Z(n_8506));
	notech_inv i_9326(.A(cacheQ[96]), .Z(n_8507));
	notech_inv i_9327(.A(cacheQ[97]), .Z(n_8508));
	notech_inv i_9328(.A(cacheQ[98]), .Z(n_8509));
	notech_inv i_9329(.A(cacheQ[99]), .Z(n_8510));
	notech_inv i_9330(.A(cacheQ[100]), .Z(n_8511));
	notech_inv i_9331(.A(cacheQ[101]), .Z(n_8512));
	notech_inv i_9332(.A(cacheQ[102]), .Z(n_8513));
	notech_inv i_9333(.A(cacheQ[103]), .Z(n_8514));
	notech_inv i_9334(.A(cacheQ[104]), .Z(n_8515));
	notech_inv i_9335(.A(cacheQ[105]), .Z(n_8516));
	notech_inv i_9336(.A(cacheQ[106]), .Z(n_8517));
	notech_inv i_9337(.A(cacheQ[107]), .Z(n_8518));
	notech_inv i_9338(.A(cacheQ[108]), .Z(n_8519));
	notech_inv i_9339(.A(cacheQ[109]), .Z(n_8520));
	notech_inv i_9340(.A(cacheQ[110]), .Z(n_8521));
	notech_inv i_9341(.A(cacheQ[111]), .Z(n_8522));
	notech_inv i_9342(.A(cacheQ[112]), .Z(n_8523));
	notech_inv i_9343(.A(cacheQ[113]), .Z(n_8524));
	notech_inv i_9344(.A(cacheQ[114]), .Z(n_8525));
	notech_inv i_9345(.A(cacheQ[115]), .Z(n_8526));
	notech_inv i_9346(.A(cacheQ[116]), .Z(n_8527));
	notech_inv i_9347(.A(cacheQ[117]), .Z(n_8528));
	notech_inv i_9348(.A(cacheQ[118]), .Z(n_8529));
	notech_inv i_9349(.A(cacheQ[119]), .Z(n_8530));
	notech_inv i_9350(.A(cacheQ[120]), .Z(n_8531));
	notech_inv i_9351(.A(cacheQ[121]), .Z(n_8532));
	notech_inv i_9352(.A(cacheQ[122]), .Z(n_8533));
	notech_inv i_9353(.A(cacheQ[123]), .Z(n_8534));
	notech_inv i_9354(.A(cacheQ[124]), .Z(n_8535));
	notech_inv i_9355(.A(cacheQ[125]), .Z(n_8536));
	notech_inv i_9356(.A(cacheQ[126]), .Z(n_8537));
	notech_inv i_9357(.A(cacheQ[127]), .Z(n_8538));
	notech_inv i_9358(.A(cacheQ[128]), .Z(n_8539));
	notech_inv i_9359(.A(cacheQ[129]), .Z(n_8540));
	notech_inv i_9360(.A(cacheQ[130]), .Z(n_8541));
	notech_inv i_9361(.A(cacheQ[131]), .Z(n_8542));
	notech_inv i_9362(.A(cacheQ[132]), .Z(n_8543));
	notech_inv i_9363(.A(cacheQ[133]), .Z(n_8544));
	notech_inv i_9364(.A(cacheQ[134]), .Z(n_8545));
	notech_inv i_9365(.A(cacheQ[135]), .Z(n_8546));
	notech_inv i_9366(.A(cacheQ[136]), .Z(n_8547));
	notech_inv i_9367(.A(cacheQ[137]), .Z(n_8548));
	notech_inv i_9368(.A(cacheQ[138]), .Z(n_8549));
	notech_inv i_9369(.A(cacheQ[139]), .Z(n_8550));
	notech_inv i_9370(.A(cacheQ[140]), .Z(n_8551));
	notech_inv i_9371(.A(cacheQ[141]), .Z(n_8552));
	notech_inv i_9372(.A(cacheQ[142]), .Z(n_8553));
	notech_inv i_9373(.A(cacheQ[143]), .Z(n_8554));
	notech_inv i_9374(.A(cacheQ[144]), .Z(n_8555));
	notech_inv i_9375(.A(cacheQ[145]), .Z(n_8556));
	notech_inv i_9376(.A(cacheQ[148]), .Z(n_8557));
	notech_inv i_9377(.A(write_msk[0]), .Z(n_8558));
	notech_inv i_9378(.A(axi_AR[31]), .Z(n_8559));
	notech_inv i_9379(.A(writeio_ack), .Z(n_8560));
	notech_inv i_9380(.A(n_62719), .Z(n_8561));
	notech_inv i_9381(.A(n_21466), .Z(n_8562));
	notech_inv i_9382(.A(write_ack), .Z(n_8563));
	notech_inv i_9383(.A(code_req), .Z(n_8564));
	notech_inv i_9384(.A(read_req), .Z(n_8565));
	notech_inv i_9385(.A(code_wreq), .Z(n_8566));
	datacache datacache1(.A(cacheA), .D(cacheD), .Q(cacheQ), .M(cacheM), .WEN
		(cacheWEN), .clk(clk));
endmodule
module AWDP_INC_23(O0, fsm5_cnt);

	output [8:0] O0;
	input [8:0] fsm5_cnt;




	notech_ha2 i_8(.A(fsm5_cnt[8]), .B(n_86), .Z(O0[8]));
	notech_ha2 i_7(.A(fsm5_cnt[7]), .B(n_84), .Z(O0[7]), .CO(n_86));
	notech_ha2 i_6(.A(fsm5_cnt[6]), .B(n_82), .Z(O0[6]), .CO(n_84));
	notech_ha2 i_5(.A(fsm5_cnt[5]), .B(n_80), .Z(O0[5]), .CO(n_82));
	notech_ha2 i_4(.A(fsm5_cnt[4]), .B(n_78), .Z(O0[4]), .CO(n_80));
	notech_ha2 i_3(.A(fsm5_cnt[3]), .B(n_76), .Z(O0[3]), .CO(n_78));
	notech_ha2 i_2(.A(fsm5_cnt[2]), .B(n_74), .Z(O0[2]), .CO(n_76));
	notech_ha2 i_1(.A(fsm5_cnt[1]), .B(fsm5_cnt[0]), .Z(O0[1]), .CO(n_74));
	notech_inv i_0(.A(fsm5_cnt[0]), .Z(O0[0]));
endmodule
module cmp14_0(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_xor2 i_10(.A(inb[2]), .B(ina[2]), .Z(n_34));
	notech_xor2 i_9(.A(inb[4]), .B(ina[4]), .Z(n_33));
	notech_xor2 i_8(.A(inb[6]), .B(ina[6]), .Z(n_32));
	notech_xor2 i_6(.A(inb[3]), .B(ina[3]), .Z(n_31));
	notech_xor2 i_5(.A(inb[5]), .B(ina[5]), .Z(n_30));
	notech_xor2 i_4(.A(inb[7]), .B(ina[7]), .Z(n_29));
	notech_xor2 i_0(.A(inb[9]), .B(ina[9]), .Z(n_55));
	notech_xor2 i_1(.A(inb[8]), .B(ina[8]), .Z(n_56));
	notech_xor2 i_3(.A(inb[1]), .B(ina[1]), .Z(n_57));
	notech_xor2 i_7(.A(inb[0]), .B(ina[0]), .Z(n_58));
	notech_or4 i_38(.A(n_57), .B(n_56), .C(n_55), .D(ina[13]), .Z(n_61));
	notech_or4 i_37(.A(n_34), .B(n_31), .C(n_33), .D(n_30), .Z(n_66));
	notech_or4 i_39(.A(n_32), .B(n_29), .C(n_58), .D(n_66), .Z(n_67));
	notech_nor2 i_2(.A(n_67), .B(n_61), .Z(out));
endmodule
module cmp14_1(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_xor2 i_10(.A(inb[2]), .B(ina[2]), .Z(n_34));
	notech_xor2 i_9(.A(inb[4]), .B(ina[4]), .Z(n_33));
	notech_xor2 i_8(.A(inb[6]), .B(ina[6]), .Z(n_32));
	notech_xor2 i_6(.A(inb[3]), .B(ina[3]), .Z(n_31));
	notech_xor2 i_5(.A(inb[5]), .B(ina[5]), .Z(n_30));
	notech_xor2 i_4(.A(inb[7]), .B(ina[7]), .Z(n_29));
	notech_xor2 i_0(.A(inb[9]), .B(ina[9]), .Z(n_55));
	notech_xor2 i_1(.A(inb[8]), .B(ina[8]), .Z(n_56));
	notech_xor2 i_3(.A(inb[1]), .B(ina[1]), .Z(n_57));
	notech_xor2 i_7(.A(inb[0]), .B(ina[0]), .Z(n_58));
	notech_or4 i_38(.A(n_57), .B(n_56), .C(n_55), .D(ina[13]), .Z(n_61));
	notech_or4 i_37(.A(n_34), .B(n_31), .C(n_33), .D(n_30), .Z(n_66));
	notech_or4 i_39(.A(n_32), .B(n_29), .C(n_58), .D(n_66), .Z(n_67));
	notech_nor2 i_2(.A(n_67), .B(n_61), .Z(out));
endmodule
module cmp14_2(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_nand2 i_41(.A(ina[10]), .B(n_63), .Z(n_62));
	notech_or2 i_0(.A(ina[12]), .B(inb[12]), .Z(n_63));
	notech_nand2 i_1(.A(inb[10]), .B(n_62), .Z(n_64));
	notech_xor2 i_26(.A(inb[5]), .B(ina[5]), .Z(n_65));
	notech_xor2 i_27(.A(inb[4]), .B(ina[4]), .Z(n_66));
	notech_xor2 i_28(.A(inb[3]), .B(ina[3]), .Z(n_68));
	notech_xor2 i_29(.A(inb[2]), .B(ina[2]), .Z(n_69));
	notech_or4 i_39(.A(n_69), .B(n_68), .C(n_66), .D(n_65), .Z(n_71));
	notech_xor2 i_30(.A(inb[1]), .B(ina[1]), .Z(n_72));
	notech_xor2 i_31(.A(inb[0]), .B(ina[0]), .Z(n_73));
	notech_xor2 i_22(.A(inb[9]), .B(ina[9]), .Z(n_75));
	notech_xor2 i_23(.A(inb[8]), .B(ina[8]), .Z(n_76));
	notech_xor2 i_24(.A(inb[7]), .B(ina[7]), .Z(n_78));
	notech_xor2 i_25(.A(inb[6]), .B(ina[6]), .Z(n_79));
	notech_or4 i_38(.A(n_79), .B(n_78), .C(n_76), .D(n_75), .Z(n_81));
	notech_ao3 i_216(.A(n_64), .B(out2), .C(ina[13]), .Z(out));
	notech_or4 i_32(.A(n_73), .B(n_72), .C(n_81), .D(n_71), .Z(out2100999)
		);
	notech_inv i_9538(.A(out2100999), .Z(out2));
endmodule
module cmp14_3(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_nand2 i_41(.A(ina[10]), .B(n_63), .Z(n_62));
	notech_or2 i_0(.A(ina[12]), .B(inb[12]), .Z(n_63));
	notech_nand2 i_1(.A(inb[10]), .B(n_62), .Z(n_64));
	notech_xor2 i_26(.A(inb[5]), .B(ina[5]), .Z(n_65));
	notech_xor2 i_27(.A(inb[4]), .B(ina[4]), .Z(n_66));
	notech_xor2 i_28(.A(inb[3]), .B(ina[3]), .Z(n_68));
	notech_xor2 i_29(.A(inb[2]), .B(ina[2]), .Z(n_69));
	notech_or4 i_39(.A(n_69), .B(n_68), .C(n_66), .D(n_65), .Z(n_71));
	notech_xor2 i_30(.A(inb[1]), .B(ina[1]), .Z(n_72));
	notech_xor2 i_31(.A(inb[0]), .B(ina[0]), .Z(n_73));
	notech_xor2 i_22(.A(inb[9]), .B(ina[9]), .Z(n_75));
	notech_xor2 i_23(.A(inb[8]), .B(ina[8]), .Z(n_76));
	notech_xor2 i_24(.A(inb[7]), .B(ina[7]), .Z(n_78));
	notech_xor2 i_25(.A(inb[6]), .B(ina[6]), .Z(n_79));
	notech_or4 i_38(.A(n_79), .B(n_78), .C(n_76), .D(n_75), .Z(n_81));
	notech_ao3 i_216(.A(n_64), .B(out2), .C(ina[13]), .Z(out));
	notech_or4 i_32(.A(n_73), .B(n_72), .C(n_81), .D(n_71), .Z(out2100998)
		);
	notech_inv i_9519(.A(out2100998), .Z(out2));
endmodule
module cmp14_4(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_nand2 i_41(.A(ina[10]), .B(n_63), .Z(n_62));
	notech_or2 i_0(.A(ina[12]), .B(inb[12]), .Z(n_63));
	notech_nand2 i_1(.A(inb[10]), .B(n_62), .Z(n_64));
	notech_xor2 i_26(.A(inb[5]), .B(ina[5]), .Z(n_65));
	notech_xor2 i_27(.A(inb[4]), .B(ina[4]), .Z(n_66));
	notech_xor2 i_28(.A(inb[3]), .B(ina[3]), .Z(n_68));
	notech_xor2 i_29(.A(inb[2]), .B(ina[2]), .Z(n_69));
	notech_or4 i_39(.A(n_69), .B(n_68), .C(n_66), .D(n_65), .Z(n_71));
	notech_xor2 i_30(.A(inb[1]), .B(ina[1]), .Z(n_72));
	notech_xor2 i_31(.A(inb[0]), .B(ina[0]), .Z(n_73));
	notech_xor2 i_22(.A(inb[9]), .B(ina[9]), .Z(n_75));
	notech_xor2 i_23(.A(inb[8]), .B(ina[8]), .Z(n_76));
	notech_xor2 i_24(.A(inb[7]), .B(ina[7]), .Z(n_78));
	notech_xor2 i_25(.A(inb[6]), .B(ina[6]), .Z(n_79));
	notech_or4 i_38(.A(n_79), .B(n_78), .C(n_76), .D(n_75), .Z(n_81));
	notech_ao3 i_216(.A(n_64), .B(out2), .C(ina[13]), .Z(out));
	notech_or4 i_32(.A(n_73), .B(n_72), .C(n_81), .D(n_71), .Z(out2100997)
		);
	notech_inv i_9500(.A(out2100997), .Z(out2));
endmodule
module cmp14_5(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_nand2 i_41(.A(ina[10]), .B(n_63), .Z(n_62));
	notech_or2 i_0(.A(ina[12]), .B(inb[12]), .Z(n_63));
	notech_nand2 i_1(.A(inb[10]), .B(n_62), .Z(n_64));
	notech_xor2 i_26(.A(inb[5]), .B(ina[5]), .Z(n_65));
	notech_xor2 i_27(.A(inb[4]), .B(ina[4]), .Z(n_66));
	notech_xor2 i_28(.A(inb[3]), .B(ina[3]), .Z(n_68));
	notech_xor2 i_29(.A(inb[2]), .B(ina[2]), .Z(n_69));
	notech_or4 i_39(.A(n_69), .B(n_68), .C(n_66), .D(n_65), .Z(n_71));
	notech_xor2 i_30(.A(inb[1]), .B(ina[1]), .Z(n_72));
	notech_xor2 i_31(.A(inb[0]), .B(ina[0]), .Z(n_73));
	notech_xor2 i_22(.A(inb[9]), .B(ina[9]), .Z(n_75));
	notech_xor2 i_23(.A(inb[8]), .B(ina[8]), .Z(n_76));
	notech_xor2 i_24(.A(inb[7]), .B(ina[7]), .Z(n_78));
	notech_xor2 i_25(.A(inb[6]), .B(ina[6]), .Z(n_79));
	notech_or4 i_38(.A(n_79), .B(n_78), .C(n_76), .D(n_75), .Z(n_81));
	notech_ao3 i_216(.A(n_64), .B(out2), .C(ina[13]), .Z(out));
	notech_or4 i_32(.A(n_73), .B(n_72), .C(n_81), .D(n_71), .Z(out2100996)
		);
	notech_inv i_9481(.A(out2100996), .Z(out2));
endmodule
module cmp14_6(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_nand2 i_41(.A(ina[10]), .B(n_63), .Z(n_62));
	notech_or2 i_0(.A(ina[12]), .B(inb[12]), .Z(n_63));
	notech_nand2 i_1(.A(inb[10]), .B(n_62), .Z(n_64));
	notech_xor2 i_26(.A(inb[5]), .B(ina[5]), .Z(n_65));
	notech_xor2 i_27(.A(inb[4]), .B(ina[4]), .Z(n_66));
	notech_xor2 i_28(.A(inb[3]), .B(ina[3]), .Z(n_68));
	notech_xor2 i_29(.A(inb[2]), .B(ina[2]), .Z(n_69));
	notech_or4 i_39(.A(n_69), .B(n_68), .C(n_66), .D(n_65), .Z(n_71));
	notech_xor2 i_30(.A(inb[1]), .B(ina[1]), .Z(n_72));
	notech_xor2 i_31(.A(inb[0]), .B(ina[0]), .Z(n_73));
	notech_xor2 i_22(.A(inb[9]), .B(ina[9]), .Z(n_75));
	notech_xor2 i_23(.A(inb[8]), .B(ina[8]), .Z(n_76));
	notech_xor2 i_24(.A(inb[7]), .B(ina[7]), .Z(n_78));
	notech_xor2 i_25(.A(inb[6]), .B(ina[6]), .Z(n_79));
	notech_or4 i_38(.A(n_79), .B(n_78), .C(n_76), .D(n_75), .Z(n_81));
	notech_ao3 i_216(.A(n_64), .B(out2), .C(ina[13]), .Z(out));
	notech_or4 i_32(.A(n_73), .B(n_72), .C(n_81), .D(n_71), .Z(out2100995)
		);
	notech_inv i_9462(.A(out2100995), .Z(out2));
endmodule
module cmp14_7(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_nand2 i_41(.A(ina[10]), .B(n_63), .Z(n_62));
	notech_or2 i_0(.A(ina[12]), .B(inb[12]), .Z(n_63));
	notech_nand2 i_1(.A(inb[10]), .B(n_62), .Z(n_64));
	notech_xor2 i_26(.A(inb[5]), .B(ina[5]), .Z(n_65));
	notech_xor2 i_27(.A(inb[4]), .B(ina[4]), .Z(n_66));
	notech_xor2 i_28(.A(inb[3]), .B(ina[3]), .Z(n_68));
	notech_xor2 i_29(.A(inb[2]), .B(ina[2]), .Z(n_69));
	notech_or4 i_39(.A(n_69), .B(n_68), .C(n_66), .D(n_65), .Z(n_71));
	notech_xor2 i_30(.A(inb[1]), .B(ina[1]), .Z(n_72));
	notech_xor2 i_31(.A(inb[0]), .B(ina[0]), .Z(n_73));
	notech_xor2 i_22(.A(inb[9]), .B(ina[9]), .Z(n_75));
	notech_xor2 i_23(.A(inb[8]), .B(ina[8]), .Z(n_76));
	notech_xor2 i_24(.A(inb[7]), .B(ina[7]), .Z(n_78));
	notech_xor2 i_25(.A(inb[6]), .B(ina[6]), .Z(n_79));
	notech_or4 i_38(.A(n_79), .B(n_78), .C(n_76), .D(n_75), .Z(n_81));
	notech_ao3 i_216(.A(n_64), .B(out2), .C(ina[13]), .Z(out));
	notech_or4 i_32(.A(n_73), .B(n_72), .C(n_81), .D(n_71), .Z(out2100994)
		);
	notech_inv i_9443(.A(out2100994), .Z(out2));
endmodule
module cmp14_8(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_nand2 i_41(.A(ina[10]), .B(n_63), .Z(n_62));
	notech_or2 i_0(.A(ina[12]), .B(inb[12]), .Z(n_63));
	notech_nand2 i_1(.A(inb[10]), .B(n_62), .Z(n_64));
	notech_xor2 i_26(.A(inb[5]), .B(ina[5]), .Z(n_65));
	notech_xor2 i_27(.A(inb[4]), .B(ina[4]), .Z(n_66));
	notech_xor2 i_28(.A(inb[3]), .B(ina[3]), .Z(n_68));
	notech_xor2 i_29(.A(inb[2]), .B(ina[2]), .Z(n_69));
	notech_or4 i_39(.A(n_69), .B(n_68), .C(n_66), .D(n_65), .Z(n_71));
	notech_xor2 i_30(.A(inb[1]), .B(ina[1]), .Z(n_72));
	notech_xor2 i_31(.A(inb[0]), .B(ina[0]), .Z(n_73));
	notech_xor2 i_22(.A(inb[9]), .B(ina[9]), .Z(n_75));
	notech_xor2 i_23(.A(inb[8]), .B(ina[8]), .Z(n_76));
	notech_xor2 i_24(.A(inb[7]), .B(ina[7]), .Z(n_78));
	notech_xor2 i_25(.A(inb[6]), .B(ina[6]), .Z(n_79));
	notech_or4 i_38(.A(n_79), .B(n_78), .C(n_76), .D(n_75), .Z(n_81));
	notech_ao3 i_216(.A(n_64), .B(out2), .C(ina[13]), .Z(out));
	notech_or4 i_32(.A(n_73), .B(n_72), .C(n_81), .D(n_71), .Z(out2100993)
		);
	notech_inv i_9424(.A(out2100993), .Z(out2));
endmodule
module cmp14_9(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_nand2 i_41(.A(ina[10]), .B(n_63), .Z(n_62));
	notech_or2 i_0(.A(ina[12]), .B(inb[12]), .Z(n_63));
	notech_nand2 i_1(.A(inb[10]), .B(n_62), .Z(n_64));
	notech_xor2 i_26(.A(inb[5]), .B(ina[5]), .Z(n_65));
	notech_xor2 i_27(.A(inb[4]), .B(ina[4]), .Z(n_66));
	notech_xor2 i_28(.A(inb[3]), .B(ina[3]), .Z(n_68));
	notech_xor2 i_29(.A(inb[2]), .B(ina[2]), .Z(n_69));
	notech_or4 i_39(.A(n_69), .B(n_68), .C(n_66), .D(n_65), .Z(n_71));
	notech_xor2 i_30(.A(inb[1]), .B(ina[1]), .Z(n_72));
	notech_xor2 i_31(.A(inb[0]), .B(ina[0]), .Z(n_73));
	notech_xor2 i_22(.A(inb[9]), .B(ina[9]), .Z(n_75));
	notech_xor2 i_23(.A(inb[8]), .B(ina[8]), .Z(n_76));
	notech_xor2 i_24(.A(inb[7]), .B(ina[7]), .Z(n_78));
	notech_xor2 i_25(.A(inb[6]), .B(ina[6]), .Z(n_79));
	notech_or4 i_38(.A(n_79), .B(n_78), .C(n_76), .D(n_75), .Z(n_81));
	notech_ao3 i_216(.A(n_64), .B(out2), .C(ina[13]), .Z(out));
	notech_or4 i_32(.A(n_73), .B(n_72), .C(n_81), .D(n_71), .Z(out2100992)
		);
	notech_inv i_9405(.A(out2100992), .Z(out2));
endmodule
module Dtlb(clk, rstn, addr_phys, cr3, cr0, data_miss, iDaddr, pg_en, iwrite_data
		, owrite_data, iread_req, iread_ack, iwrite_req, iwrite_ack, iread_sz
		, oread_sz, iwrite_sz, owrite_sz, oread_req, oread_ack, owrite_req
		, owrite_ack, pg_fault, wr_fault, cr2, flush_tlb, cs, pt_fault, busy_ram
		, outstanding);

	input clk;
	input rstn;
	output [31:0] addr_phys;
	input [31:0] cr3;
	input [31:0] cr0;
	input [31:0] data_miss;
	input [31:0] iDaddr;
	input pg_en;
	input [31:0] iwrite_data;
	output [31:0] owrite_data;
	input iread_req;
	input iread_ack;
	input iwrite_req;
	input iwrite_ack;
	input [1:0] iread_sz;
	output [1:0] oread_sz;
	input [1:0] iwrite_sz;
	output [1:0] owrite_sz;
	output oread_req;
	output oread_ack;
	output owrite_req;
	output owrite_ack;
	output pg_fault;
	output wr_fault;
	output [31:0] cr2;
	input flush_tlb;
	input [31:0] cs;
	output pt_fault;
	input busy_ram;
	output outstanding;

	wire [3:0] fsm;
	wire [31:0] addr_miss;
	wire [31:0] wrA;
	wire [31:0] iDaddr_f;
	wire [31:0] wrD;
	wire [1:0] nx_dir;
	wire [8:0] fsm5_cnt_0;
	wire [8:0] fsm5_cnt;



	notech_inv i_14914(.A(n_63053), .Z(n_63080));
	notech_inv i_14913(.A(n_63053), .Z(n_63079));
	notech_inv i_14912(.A(n_63053), .Z(n_63078));
	notech_inv i_14910(.A(n_63053), .Z(n_63076));
	notech_inv i_14909(.A(n_63053), .Z(n_63075));
	notech_inv i_14908(.A(n_63053), .Z(n_63074));
	notech_inv i_14905(.A(n_63053), .Z(n_63071));
	notech_inv i_14904(.A(n_63053), .Z(n_63070));
	notech_inv i_14903(.A(n_63053), .Z(n_63069));
	notech_inv i_14901(.A(n_63053), .Z(n_63067));
	notech_inv i_14900(.A(n_63053), .Z(n_63066));
	notech_inv i_14899(.A(n_63053), .Z(n_63065));
	notech_inv i_14896(.A(n_63053), .Z(n_63062));
	notech_inv i_14895(.A(n_63053), .Z(n_63061));
	notech_inv i_14894(.A(n_63053), .Z(n_63060));
	notech_inv i_14892(.A(n_63053), .Z(n_63058));
	notech_inv i_14891(.A(n_63053), .Z(n_63057));
	notech_inv i_14890(.A(n_63053), .Z(n_63056));
	notech_inv i_14887(.A(clk), .Z(n_63053));
	notech_inv i_14886(.A(n_63025), .Z(n_63052));
	notech_inv i_14885(.A(n_63025), .Z(n_63051));
	notech_inv i_14884(.A(n_63025), .Z(n_63050));
	notech_inv i_14882(.A(n_63025), .Z(n_63048));
	notech_inv i_14881(.A(n_63025), .Z(n_63047));
	notech_inv i_14880(.A(n_63025), .Z(n_63046));
	notech_inv i_14877(.A(n_63025), .Z(n_63043));
	notech_inv i_14876(.A(n_63025), .Z(n_63042));
	notech_inv i_14875(.A(n_63025), .Z(n_63041));
	notech_inv i_14873(.A(n_63025), .Z(n_63039));
	notech_inv i_14872(.A(n_63025), .Z(n_63038));
	notech_inv i_14871(.A(n_63025), .Z(n_63037));
	notech_inv i_14868(.A(n_63025), .Z(n_63034));
	notech_inv i_14867(.A(n_63025), .Z(n_63033));
	notech_inv i_14866(.A(n_63025), .Z(n_63032));
	notech_inv i_14864(.A(n_63025), .Z(n_63030));
	notech_inv i_14863(.A(n_63025), .Z(n_63029));
	notech_inv i_14862(.A(n_63025), .Z(n_63028));
	notech_inv i_14859(.A(clk), .Z(n_63025));
	notech_inv i_14858(.A(n_62997), .Z(n_63024));
	notech_inv i_14857(.A(n_62997), .Z(n_63023));
	notech_inv i_14856(.A(n_62997), .Z(n_63022));
	notech_inv i_14854(.A(n_62997), .Z(n_63020));
	notech_inv i_14853(.A(n_62997), .Z(n_63019));
	notech_inv i_14852(.A(n_62997), .Z(n_63018));
	notech_inv i_14849(.A(n_62997), .Z(n_63015));
	notech_inv i_14848(.A(n_62997), .Z(n_63014));
	notech_inv i_14847(.A(n_62997), .Z(n_63013));
	notech_inv i_14845(.A(n_62997), .Z(n_63011));
	notech_inv i_14844(.A(n_62997), .Z(n_63010));
	notech_inv i_14843(.A(n_62997), .Z(n_63009));
	notech_inv i_14840(.A(n_62997), .Z(n_63006));
	notech_inv i_14838(.A(n_62997), .Z(n_63004));
	notech_inv i_14835(.A(n_62997), .Z(n_63001));
	notech_inv i_14834(.A(n_62997), .Z(n_63000));
	notech_inv i_14831(.A(clk), .Z(n_62997));
	notech_inv i_14736(.A(n_62892), .Z(n_62899));
	notech_inv i_14735(.A(n_62892), .Z(n_62898));
	notech_inv i_14730(.A(n_62892), .Z(n_62893));
	notech_inv i_14729(.A(pg_en), .Z(n_62892));
	notech_inv i_14188(.A(n_62319), .Z(n_62346));
	notech_inv i_14187(.A(n_62319), .Z(n_62345));
	notech_inv i_14186(.A(n_62319), .Z(n_62344));
	notech_inv i_14184(.A(n_62319), .Z(n_62342));
	notech_inv i_14183(.A(n_62319), .Z(n_62341));
	notech_inv i_14182(.A(n_62319), .Z(n_62340));
	notech_inv i_14179(.A(n_62319), .Z(n_62337));
	notech_inv i_14178(.A(n_62319), .Z(n_62336));
	notech_inv i_14177(.A(n_62319), .Z(n_62335));
	notech_inv i_14175(.A(n_62319), .Z(n_62333));
	notech_inv i_14174(.A(n_62319), .Z(n_62332));
	notech_inv i_14173(.A(n_62319), .Z(n_62331));
	notech_inv i_14170(.A(n_62319), .Z(n_62328));
	notech_inv i_14169(.A(n_62319), .Z(n_62327));
	notech_inv i_14168(.A(n_62319), .Z(n_62326));
	notech_inv i_14166(.A(n_62319), .Z(n_62324));
	notech_inv i_14165(.A(n_62319), .Z(n_62323));
	notech_inv i_14164(.A(n_62319), .Z(n_62322));
	notech_inv i_14161(.A(rstn), .Z(n_62319));
	notech_inv i_14160(.A(n_62291), .Z(n_62318));
	notech_inv i_14159(.A(n_62291), .Z(n_62317));
	notech_inv i_14158(.A(n_62291), .Z(n_62316));
	notech_inv i_14156(.A(n_62291), .Z(n_62314));
	notech_inv i_14155(.A(n_62291), .Z(n_62313));
	notech_inv i_14154(.A(n_62291), .Z(n_62312));
	notech_inv i_14151(.A(n_62291), .Z(n_62309));
	notech_inv i_14150(.A(n_62291), .Z(n_62308));
	notech_inv i_14149(.A(n_62291), .Z(n_62307));
	notech_inv i_14147(.A(n_62291), .Z(n_62305));
	notech_inv i_14146(.A(n_62291), .Z(n_62304));
	notech_inv i_14145(.A(n_62291), .Z(n_62303));
	notech_inv i_14142(.A(n_62291), .Z(n_62300));
	notech_inv i_14141(.A(n_62291), .Z(n_62299));
	notech_inv i_14140(.A(n_62291), .Z(n_62298));
	notech_inv i_14138(.A(n_62291), .Z(n_62296));
	notech_inv i_14137(.A(n_62291), .Z(n_62295));
	notech_inv i_14136(.A(n_62291), .Z(n_62294));
	notech_inv i_14133(.A(rstn), .Z(n_62291));
	notech_inv i_14132(.A(n_62263), .Z(n_62290));
	notech_inv i_14131(.A(n_62263), .Z(n_62289));
	notech_inv i_14130(.A(n_62263), .Z(n_62288));
	notech_inv i_14128(.A(n_62263), .Z(n_62286));
	notech_inv i_14127(.A(n_62263), .Z(n_62285));
	notech_inv i_14126(.A(n_62263), .Z(n_62284));
	notech_inv i_14123(.A(n_62263), .Z(n_62281));
	notech_inv i_14122(.A(n_62263), .Z(n_62280));
	notech_inv i_14121(.A(n_62263), .Z(n_62279));
	notech_inv i_14119(.A(n_62263), .Z(n_62277));
	notech_inv i_14118(.A(n_62263), .Z(n_62276));
	notech_inv i_14117(.A(n_62263), .Z(n_62275));
	notech_inv i_14114(.A(n_62263), .Z(n_62272));
	notech_inv i_14112(.A(n_62263), .Z(n_62270));
	notech_inv i_14109(.A(n_62263), .Z(n_62267));
	notech_inv i_14108(.A(n_62263), .Z(n_62266));
	notech_inv i_14105(.A(rstn), .Z(n_62263));
	notech_inv i_10763(.A(n_58742), .Z(n_58743));
	notech_inv i_10762(.A(n_948), .Z(n_58742));
	notech_inv i_10754(.A(n_58733), .Z(n_58734));
	notech_inv i_10753(.A(hit_tab21), .Z(n_58733));
	notech_inv i_10745(.A(n_58724), .Z(n_58725));
	notech_inv i_10744(.A(hit_tab11), .Z(n_58724));
	notech_inv i_8497(.A(n_56309), .Z(n_56310));
	notech_inv i_8496(.A(\nbus_14514[0] ), .Z(n_56309));
	notech_inv i_8489(.A(n_56300), .Z(n_56301));
	notech_inv i_8488(.A(n_1043), .Z(n_56300));
	notech_inv i_8479(.A(n_56289), .Z(n_56290));
	notech_inv i_8478(.A(n_1040), .Z(n_56289));
	notech_inv i_8361(.A(n_56176), .Z(n_56177));
	notech_inv i_8360(.A(\nbus_14517[0] ), .Z(n_56176));
	notech_inv i_8353(.A(n_56167), .Z(n_56168));
	notech_inv i_8352(.A(n_11870), .Z(n_56167));
	notech_inv i_8345(.A(n_56158), .Z(n_56159));
	notech_inv i_8344(.A(\nbus_14520[0] ), .Z(n_56158));
	notech_inv i_8340(.A(n_56147), .Z(n_56153));
	notech_inv i_8335(.A(n_56147), .Z(n_56148));
	notech_inv i_8334(.A(n_56825), .Z(n_56147));
	notech_inv i_8327(.A(n_56138), .Z(n_56139));
	notech_inv i_8326(.A(\nbus_14503[0] ), .Z(n_56138));
	notech_inv i_8319(.A(n_56129), .Z(n_56130));
	notech_inv i_8318(.A(\nbus_14511[0] ), .Z(n_56129));
	notech_inv i_8311(.A(n_56120), .Z(n_56121));
	notech_inv i_8310(.A(\nbus_14502[0] ), .Z(n_56120));
	notech_inv i_8301(.A(n_56109), .Z(n_56110));
	notech_inv i_8300(.A(\nbus_14516[0] ), .Z(n_56109));
	notech_inv i_8293(.A(n_56100), .Z(n_56101));
	notech_inv i_8292(.A(\nbus_14508[0] ), .Z(n_56100));
	notech_inv i_8285(.A(n_56091), .Z(n_56092));
	notech_inv i_8284(.A(\nbus_14510[0] ), .Z(n_56091));
	notech_inv i_8277(.A(n_56082), .Z(n_56083));
	notech_inv i_8276(.A(\nbus_14492[0] ), .Z(n_56082));
	notech_inv i_8269(.A(n_56073), .Z(n_56074));
	notech_inv i_8268(.A(\nbus_14489[0] ), .Z(n_56073));
	notech_inv i_7803(.A(n_55558), .Z(n_55559));
	notech_inv i_7802(.A(n_945), .Z(n_55558));
	notech_inv i_7751(.A(n_55410), .Z(n_55416));
	notech_inv i_7746(.A(n_55410), .Z(n_55411));
	notech_inv i_7745(.A(n_1042), .Z(n_55410));
	notech_inv i_7743(.A(n_1085), .Z(n_55407));
	notech_inv i_7742(.A(n_1085), .Z(n_55406));
	notech_inv i_7738(.A(n_1085), .Z(n_55402));
	notech_inv i_7730(.A(n_55392), .Z(n_55393));
	notech_inv i_7729(.A(n_1098), .Z(n_55392));
	notech_inv i_7722(.A(n_55383), .Z(n_55384));
	notech_inv i_7721(.A(n_1081), .Z(n_55383));
	notech_inv i_7719(.A(\nbus_14488[0] ), .Z(n_55307));
	notech_inv i_7717(.A(\nbus_14488[0] ), .Z(n_55305));
	notech_inv i_7714(.A(\nbus_14488[0] ), .Z(n_55302));
	notech_inv i_7712(.A(\nbus_14488[0] ), .Z(n_55300));
	notech_xor2 i_149(.A(n_11990), .B(\nnx_tab2[0] ), .Z(n_573));
	notech_or4 i_139(.A(hit_adr23), .B(hit_adr24), .C(hit_adr22), .D(hit_adr21
		), .Z(n_571));
	notech_ao4 i_148(.A(hit_adr22), .B(n_1024), .C(n_11995), .D(n_1025), .Z(n_564
		));
	notech_nor2 i_96(.A(hit_adr24), .B(\nx_tab2[0] ), .Z(n_562));
	notech_nor2 i_607(.A(hit_adr23), .B(n_562), .Z(n_561));
	notech_nor2 i_147(.A(hit_adr22), .B(n_561), .Z(n_559));
	notech_or4 i_604(.A(n_1001), .B(n_1010), .C(\nx_tab1[1] ), .D(\nx_tab1[0] 
		), .Z(n_557));
	notech_or2 i_79(.A(fsm5_cnt[2]), .B(fsm5_cnt[3]), .Z(n_556));
	notech_and3 i_603(.A(fsm5_cnt[4]), .B(fsm5_cnt[5]), .C(n_556), .Z(n_555)
		);
	notech_or2 i_153(.A(fsm5_cnt[6]), .B(n_555), .Z(n_554));
	notech_and2 i_602(.A(fsm5_cnt[7]), .B(n_554), .Z(n_553));
	notech_or4 i_601(.A(fsm5_cnt[8]), .B(n_1028), .C(n_553), .D(n_12166), .Z
		(n_552));
	notech_ao3 i_78675(.A(data_miss[5]), .B(n_960), .C(n_972), .Z(n_550));
	notech_nao3 i_596(.A(n_995), .B(n_11847), .C(n_550), .Z(n_549));
	notech_or4 i_145(.A(hit_dir2), .B(\hit_dir1[7] ), .C(n_972), .D(busy_ram
		), .Z(n_547));
	notech_ao4 i_144(.A(n_12000), .B(n_11998), .C(fsm[0]), .D(n_12001), .Z(n_546
		));
	notech_or4 i_589(.A(fsm[2]), .B(fsm[1]), .C(n_1015), .D(n_12166), .Z(n_545
		));
	notech_xor2 i_143(.A(fsm[0]), .B(iwrite_ack), .Z(n_541));
	notech_nao3 i_142(.A(n_1043), .B(n_947), .C(n_946), .Z(n_538));
	notech_ao4 i_141(.A(iwrite_req), .B(n_62899), .C(n_946), .D(n_1053), .Z(n_536
		));
	notech_nand2 i_575(.A(\dir2[29] ), .B(n_1055), .Z(n_534));
	notech_nand2 i_572(.A(\dir2[28] ), .B(n_1055), .Z(n_533));
	notech_nand2 i_569(.A(\dir2[27] ), .B(n_1055), .Z(n_532));
	notech_nand2 i_566(.A(\dir2[26] ), .B(n_1055), .Z(n_531));
	notech_nand2 i_563(.A(\dir2[25] ), .B(n_1055), .Z(n_530));
	notech_nand2 i_560(.A(\dir2[24] ), .B(n_1055), .Z(n_529));
	notech_nand2 i_557(.A(\dir2[23] ), .B(n_1055), .Z(n_528));
	notech_nand2 i_554(.A(\dir2[22] ), .B(n_1055), .Z(n_527));
	notech_nand2 i_551(.A(\dir2[21] ), .B(n_1055), .Z(n_526));
	notech_nand2 i_548(.A(\dir2[20] ), .B(n_1055), .Z(n_525));
	notech_nand2 i_545(.A(\dir2[19] ), .B(n_1055), .Z(n_524));
	notech_nand2 i_542(.A(\dir2[18] ), .B(n_1055), .Z(n_523));
	notech_nand2 i_539(.A(\dir2[17] ), .B(n_1055), .Z(n_522));
	notech_nand2 i_536(.A(\dir2[16] ), .B(n_1055), .Z(n_521));
	notech_nand2 i_533(.A(\dir2[15] ), .B(n_1055), .Z(n_520));
	notech_nand2 i_530(.A(\dir2[14] ), .B(n_1055), .Z(n_519));
	notech_nand2 i_527(.A(\dir2[13] ), .B(n_1055), .Z(n_518));
	notech_nand2 i_524(.A(\dir2[12] ), .B(n_1055), .Z(n_517));
	notech_nand2 i_520(.A(\dir2[11] ), .B(n_1055), .Z(n_516));
	notech_nand2 i_517(.A(\dir2[10] ), .B(n_1055), .Z(n_515));
	notech_nand3 i_494(.A(n_56896), .B(iread_ack), .C(n_62899), .Z(n_494));
	notech_nao3 i_491(.A(n_406), .B(n_11844), .C(req_miss), .Z(n_491));
	notech_xor2 i_140(.A(iread_req), .B(iread_ack), .Z(n_490));
	notech_nand3 i_266(.A(n_62899), .B(n_11843), .C(wrA[11]), .Z(n_487));
	notech_and2 i_18(.A(n_62899), .B(n_1080), .Z(n_486));
	notech_nand3 i_263(.A(n_62899), .B(n_11843), .C(wrA[10]), .Z(n_485));
	notech_nand3 i_260(.A(n_62899), .B(n_11843), .C(wrA[9]), .Z(n_484));
	notech_nand3 i_257(.A(n_62898), .B(n_11843), .C(wrA[8]), .Z(n_483));
	notech_nand3 i_254(.A(n_62898), .B(n_11843), .C(wrA[7]), .Z(n_482));
	notech_nand3 i_251(.A(n_62898), .B(n_11843), .C(wrA[6]), .Z(n_481));
	notech_nand3 i_248(.A(n_62898), .B(n_11843), .C(wrA[5]), .Z(n_480));
	notech_nand3 i_245(.A(n_62898), .B(n_11843), .C(wrA[4]), .Z(n_479));
	notech_nand3 i_242(.A(n_62898), .B(n_11843), .C(wrA[3]), .Z(n_478));
	notech_nand3 i_239(.A(n_62899), .B(n_11843), .C(wrA[2]), .Z(n_477));
	notech_nand3 i_236(.A(n_62899), .B(n_11843), .C(wrA[1]), .Z(n_476));
	notech_nand3 i_233(.A(n_62899), .B(wrA[0]), .C(n_11843), .Z(n_475));
	notech_and4 i_157(.A(n_995), .B(n_11847), .C(iread_ack), .D(n_62899), .Z
		(n_410));
	notech_ao3 i_156(.A(n_62899), .B(n_1030), .C(n_1028), .Z(n_409));
	notech_nand2 i_146(.A(n_1032), .B(n_12001), .Z(n_408));
	notech_nand2 i_137(.A(n_986), .B(n_62899), .Z(n_407));
	notech_nand3 i_82(.A(n_983), .B(iread_req), .C(n_11895), .Z(n_406));
	notech_or4 i_619(.A(n_1001), .B(n_1002), .C(n_11993), .D(n_11995), .Z(n_577
		));
	notech_or4 i_620(.A(n_1001), .B(n_1002), .C(n_11995), .D(\nx_tab2[0] ), 
		.Z(n_578));
	notech_or4 i_621(.A(n_1001), .B(n_1002), .C(\nx_tab2[1] ), .D(n_11993), 
		.Z(n_579));
	notech_or4 i_138(.A(hit_adr13), .B(hit_adr14), .C(hit_adr12), .D(hit_adr11
		), .Z(n_583));
	notech_xor2 i_150(.A(\nnx_tab1[1] ), .B(n_11922), .Z(n_585));
	notech_nor2 i_151(.A(hit_adr12), .B(n_592), .Z(n_590));
	notech_nor2 i_631(.A(hit_adr13), .B(n_593), .Z(n_592));
	notech_nor2 i_128(.A(hit_adr14), .B(\nx_tab1[0] ), .Z(n_593));
	notech_ao4 i_152(.A(hit_adr12), .B(n_1018), .C(n_11920), .D(n_1019), .Z(n_595
		));
	notech_or4 i_636(.A(n_1001), .B(n_1010), .C(n_11918), .D(n_11920), .Z(n_599
		));
	notech_or4 i_637(.A(n_1001), .B(n_1010), .C(n_11920), .D(\nx_tab1[0] ), 
		.Z(n_600));
	notech_or4 i_638(.A(n_1001), .B(\nx_tab1[1] ), .C(n_1010), .D(n_11918), 
		.Z(n_601));
	notech_or4 i_641(.A(n_1001), .B(n_1002), .C(\nx_tab2[1] ), .D(\nx_tab2[0] 
		), .Z(n_604));
	notech_nao3 i_642(.A(iwrite_req), .B(n_606), .C(data_miss[1]), .Z(n_605)
		);
	notech_nao3 i_92(.A(n_12138), .B(n_12139), .C(cs[0]), .Z(n_606));
	notech_or4 i_661(.A(data_miss[0]), .B(n_989), .C(n_12167), .D(n_12166), 
		.Z(n_625));
	notech_nor2 i_662(.A(n_627), .B(n_977), .Z(n_626));
	notech_nor2 i_70(.A(nx_dir[0]), .B(nx_dir[1]), .Z(n_627));
	notech_nand3 i_663(.A(flush_tlb), .B(n_62899), .C(n_11895), .Z(n_628));
	notech_nand2 i_667(.A(n_627), .B(n_12140), .Z(n_631));
	notech_and2 i_689(.A(\hit_dir1[7] ), .B(n_653), .Z(n_652));
	notech_or4 i_154(.A(hit_tab12), .B(hit_tab11), .C(hit_tab13), .D(hit_tab14
		), .Z(n_653));
	notech_and2 i_690(.A(hit_dir2), .B(n_655), .Z(n_654));
	notech_or4 i_155(.A(hit_tab22), .B(hit_tab24), .C(hit_tab21), .D(hit_tab23
		), .Z(n_655));
	notech_ao3 i_759(.A(n_974), .B(n_999), .C(data_miss[1]), .Z(n_656));
	notech_nand3 i_275(.A(n_55407), .B(\tab13[10] ), .C(n_1096), .Z(n_685)
		);
	notech_nand3 i_272(.A(hit_tab11), .B(\tab11[10] ), .C(n_55406), .Z(n_688
		));
	notech_nao3 i_269(.A(hit_tab21), .B(\tab21[10] ), .C(n_1081), .Z(n_691)
		);
	notech_nand3 i_286(.A(n_55407), .B(n_1096), .C(\tab13[11] ), .Z(n_696)
		);
	notech_nand3 i_283(.A(hit_tab11), .B(n_55407), .C(\tab11[11] ), .Z(n_699
		));
	notech_nao3 i_280(.A(hit_tab21), .B(\tab21[11] ), .C(n_1081), .Z(n_702)
		);
	notech_nand3 i_297(.A(n_55407), .B(n_1096), .C(\tab13[12] ), .Z(n_707)
		);
	notech_nand3 i_294(.A(hit_tab11), .B(n_55406), .C(\tab11[12] ), .Z(n_710
		));
	notech_nao3 i_291(.A(hit_tab21), .B(\tab21[12] ), .C(n_1081), .Z(n_713)
		);
	notech_nand3 i_308(.A(n_55406), .B(n_1096), .C(\tab13[13] ), .Z(n_718)
		);
	notech_nand3 i_305(.A(hit_tab11), .B(n_55406), .C(\tab11[13] ), .Z(n_721
		));
	notech_nao3 i_302(.A(hit_tab21), .B(\tab21[13] ), .C(n_1081), .Z(n_724)
		);
	notech_nand3 i_319(.A(n_55406), .B(n_1096), .C(\tab13[14] ), .Z(n_729)
		);
	notech_nand3 i_316(.A(hit_tab11), .B(n_55406), .C(\tab11[14] ), .Z(n_732
		));
	notech_nao3 i_313(.A(hit_tab21), .B(\tab21[14] ), .C(n_1081), .Z(n_735)
		);
	notech_nand3 i_330(.A(n_55407), .B(n_1096), .C(\tab13[15] ), .Z(n_740)
		);
	notech_nand3 i_327(.A(hit_tab11), .B(n_55407), .C(\tab11[15] ), .Z(n_743
		));
	notech_nao3 i_324(.A(hit_tab21), .B(\tab21[15] ), .C(n_1081), .Z(n_746)
		);
	notech_nand3 i_341(.A(n_55407), .B(n_1096), .C(\tab13[16] ), .Z(n_751)
		);
	notech_nand3 i_338(.A(hit_tab11), .B(n_55407), .C(\tab11[16] ), .Z(n_754
		));
	notech_nao3 i_335(.A(hit_tab21), .B(\tab21[16] ), .C(n_1081), .Z(n_757)
		);
	notech_nand3 i_352(.A(n_55407), .B(n_1096), .C(\tab13[17] ), .Z(n_762)
		);
	notech_nand3 i_349(.A(hit_tab11), .B(n_55407), .C(\tab11[17] ), .Z(n_765
		));
	notech_nao3 i_346(.A(hit_tab21), .B(\tab21[17] ), .C(n_1081), .Z(n_768)
		);
	notech_nand3 i_363(.A(n_55407), .B(n_1096), .C(\tab13[18] ), .Z(n_773)
		);
	notech_nand3 i_360(.A(hit_tab11), .B(n_55407), .C(\tab11[18] ), .Z(n_776
		));
	notech_nao3 i_357(.A(hit_tab21), .B(\tab21[18] ), .C(n_1081), .Z(n_779)
		);
	notech_nand3 i_374(.A(n_55407), .B(n_1096), .C(\tab13[19] ), .Z(n_784)
		);
	notech_nand3 i_371(.A(hit_tab11), .B(n_55407), .C(\tab11[19] ), .Z(n_787
		));
	notech_nao3 i_368(.A(hit_tab21), .B(\tab21[19] ), .C(n_1081), .Z(n_790)
		);
	notech_nand3 i_385(.A(n_55406), .B(n_1096), .C(\tab13[20] ), .Z(n_795)
		);
	notech_nand3 i_382(.A(hit_tab11), .B(n_55402), .C(\tab11[20] ), .Z(n_798
		));
	notech_nao3 i_379(.A(hit_tab21), .B(\tab21[20] ), .C(n_1081), .Z(n_801)
		);
	notech_nand3 i_396(.A(n_55402), .B(n_1096), .C(\tab13[21] ), .Z(n_806)
		);
	notech_nand3 i_393(.A(n_58725), .B(n_55402), .C(\tab11[21] ), .Z(n_809)
		);
	notech_nao3 i_390(.A(n_58734), .B(\tab21[21] ), .C(n_1081), .Z(n_812));
	notech_nand3 i_407(.A(n_55402), .B(n_1096), .C(\tab13[22] ), .Z(n_817)
		);
	notech_nand3 i_404(.A(n_58725), .B(n_55402), .C(\tab11[22] ), .Z(n_820)
		);
	notech_nao3 i_401(.A(n_58734), .B(\tab21[22] ), .C(n_55384), .Z(n_823)
		);
	notech_nand3 i_418(.A(n_55402), .B(n_1096), .C(\tab13[23] ), .Z(n_828)
		);
	notech_nand3 i_415(.A(n_58725), .B(n_55402), .C(\tab11[23] ), .Z(n_831)
		);
	notech_nao3 i_412(.A(n_58734), .B(\tab21[23] ), .C(n_55384), .Z(n_834)
		);
	notech_nand3 i_429(.A(n_55402), .B(n_1096), .C(\tab13[24] ), .Z(n_839)
		);
	notech_nand3 i_426(.A(n_58725), .B(n_55402), .C(\tab11[24] ), .Z(n_842)
		);
	notech_nao3 i_423(.A(n_58734), .B(\tab21[24] ), .C(n_55384), .Z(n_845)
		);
	notech_nand3 i_440(.A(n_55402), .B(n_1096), .C(\tab13[25] ), .Z(n_850)
		);
	notech_nand3 i_437(.A(n_58725), .B(n_55406), .C(\tab11[25] ), .Z(n_853)
		);
	notech_nao3 i_434(.A(n_58734), .B(\tab21[25] ), .C(n_55384), .Z(n_856)
		);
	notech_nand3 i_451(.A(n_55406), .B(n_1096), .C(\tab13[26] ), .Z(n_861)
		);
	notech_nand3 i_448(.A(n_58725), .B(n_55406), .C(\tab11[26] ), .Z(n_864)
		);
	notech_nao3 i_445(.A(n_58734), .B(\tab21[26] ), .C(n_55384), .Z(n_867)
		);
	notech_nand3 i_462(.A(n_55406), .B(n_1096), .C(\tab13[27] ), .Z(n_872)
		);
	notech_nand3 i_459(.A(n_58725), .B(n_55406), .C(\tab11[27] ), .Z(n_875)
		);
	notech_nao3 i_456(.A(n_58734), .B(\tab21[27] ), .C(n_55384), .Z(n_878)
		);
	notech_nand3 i_473(.A(n_55402), .B(n_1096), .C(\tab13[28] ), .Z(n_883)
		);
	notech_nand3 i_470(.A(n_58725), .B(n_55402), .C(\tab11[28] ), .Z(n_886)
		);
	notech_nao3 i_467(.A(n_58734), .B(\tab21[28] ), .C(n_55384), .Z(n_889)
		);
	notech_nand3 i_484(.A(n_55402), .B(n_1096), .C(\tab13[29] ), .Z(n_894)
		);
	notech_nand3 i_481(.A(n_58725), .B(n_55406), .C(\tab11[29] ), .Z(n_897)
		);
	notech_nao3 i_478(.A(n_58734), .B(\tab21[29] ), .C(n_55384), .Z(n_900)
		);
	notech_and2 i_982(.A(iwrite_sz[0]), .B(n_55416), .Z(n_901));
	notech_and2 i_983(.A(iwrite_sz[1]), .B(n_55416), .Z(n_902));
	notech_nao3 i_489(.A(n_62899), .B(n_1077), .C(iread_ack), .Z(n_903));
	notech_nand2 i_490(.A(n_490), .B(n_12166), .Z(n_904));
	notech_nand3 i_90(.A(iread_ack), .B(n_62899), .C(n_11996), .Z(n_945));
	notech_and3 i_84(.A(n_983), .B(iwrite_req), .C(n_11895), .Z(n_946));
	notech_nand2 i_580(.A(iwrite_req), .B(n_1053), .Z(n_947));
	notech_or4 i_91(.A(fsm[0]), .B(fsm[2]), .C(fsm[1]), .D(fsm[3]), .Z(n_948
		));
	notech_and4 i_583(.A(n_11847), .B(n_988), .C(data_miss[0]), .D(data_miss
		[5]), .Z(n_951));
	notech_or4 i_586(.A(n_954), .B(n_992), .C(n_972), .D(n_1005), .Z(n_952)
		);
	notech_or4 i_587(.A(fsm[2]), .B(fsm[1]), .C(n_12001), .D(n_12166), .Z(n_953
		));
	notech_ao4 i_67(.A(hit_dir2), .B(\hit_dir1[7] ), .C(pg_fault), .D(n_983)
		, .Z(n_954));
	notech_nao3 i_592(.A(n_547), .B(n_11847), .C(n_984), .Z(n_957));
	notech_or2 i_597(.A(iread_req), .B(data_miss[6]), .Z(n_960));
	notech_and2 i_1021(.A(iwrite_ack), .B(n_408), .Z(n_961));
	notech_and4 i_1022(.A(fsm[0]), .B(fsm5_cnt_0[0]), .C(n_12001), .D(n_995)
		, .Z(n_962));
	notech_and4 i_1024(.A(fsm[0]), .B(n_995), .C(fsm5_cnt_0[1]), .D(n_12001)
		, .Z(n_963));
	notech_and4 i_1025(.A(fsm[0]), .B(n_995), .C(fsm5_cnt_0[2]), .D(n_12001)
		, .Z(n_964));
	notech_and4 i_1026(.A(fsm[0]), .B(n_995), .C(fsm5_cnt_0[3]), .D(n_12001)
		, .Z(n_965));
	notech_and4 i_1027(.A(fsm[0]), .B(n_995), .C(fsm5_cnt_0[4]), .D(n_12001)
		, .Z(n_966));
	notech_and4 i_1028(.A(fsm[0]), .B(n_995), .C(fsm5_cnt_0[5]), .D(n_12001)
		, .Z(n_967));
	notech_and4 i_1029(.A(fsm[0]), .B(n_995), .C(fsm5_cnt_0[6]), .D(n_12001)
		, .Z(n_968));
	notech_and4 i_1030(.A(fsm[0]), .B(n_995), .C(fsm5_cnt_0[7]), .D(n_12001)
		, .Z(n_969));
	notech_and4 i_1031(.A(fsm[0]), .B(n_995), .C(fsm5_cnt_0[8]), .D(n_12001)
		, .Z(n_970));
	notech_or4 i_1053(.A(n_972), .B(n_992), .C(n_1006), .D(n_1007), .Z(n_971
		));
	notech_nor2 i_4(.A(iwrite_req), .B(iread_req), .Z(n_972));
	notech_nor2 i_1063(.A(n_996), .B(n_12156), .Z(n_973));
	notech_and3 i_136(.A(n_995), .B(iwrite_req), .C(n_11847), .Z(n_974));
	notech_and3 i_1065(.A(n_995), .B(data_miss[1]), .C(n_11847), .Z(n_975)
		);
	notech_and4 i_1066(.A(n_988), .B(data_miss[0]), .C(n_11847), .D(\dir1_0[4] 
		), .Z(n_976));
	notech_nao3 i_94(.A(data_miss[0]), .B(n_11844), .C(n_989), .Z(n_977));
	notech_and2 i_1069(.A(iwrite_ack), .B(n_407), .Z(owrite_ack));
	notech_reg nx_dir_reg_0(.CP(n_63056), .D(n_8577), .CD(n_62322), .Q(nx_dir
		[0]));
	notech_mux2 i_9572(.S(n_977), .A(n_627), .B(nx_dir[0]), .Z(n_8577));
	notech_or2 i_78692(.A(n_654), .B(n_652), .Z(n_983));
	notech_reg nx_dir_reg_1(.CP(n_63056), .D(n_8587), .CD(n_62322), .Q(nx_dir
		[1]));
	notech_nand2 i_129(.A(n_12000), .B(n_11998), .Z(n_984));
	notech_ao3 i_9584(.A(nx_dir[1]), .B(1'b1), .C(n_12140), .Z(n_8587));
	notech_reg iDaddr_f_reg_0(.CP(n_63056), .D(n_8589), .CD(n_62322), .Q(iDaddr_f
		[0]));
	notech_mux2 i_9588(.S(n_948), .A(iDaddr[0]), .B(iDaddr_f[0]), .Z(n_8589)
		);
	notech_or2 i_130(.A(fsm[0]), .B(fsm[3]), .Z(n_985));
	notech_reg iDaddr_f_reg_1(.CP(n_63056), .D(n_8595), .CD(n_62322), .Q(iDaddr_f
		[1]));
	notech_mux2 i_9596(.S(n_948), .A(iDaddr[1]), .B(iDaddr_f[1]), .Z(n_8595)
		);
	notech_nao3 i_7(.A(n_983), .B(n_11847), .C(n_984), .Z(n_986));
	notech_reg iDaddr_f_reg_2(.CP(n_63056), .D(n_8601), .CD(n_62322), .Q(iDaddr_f
		[2]));
	notech_mux2 i_9604(.S(n_948), .A(iDaddr[2]), .B(iDaddr_f[2]), .Z(n_8601)
		);
	notech_nand2 i_11(.A(iread_ack), .B(n_62899), .Z(n_987));
	notech_reg iDaddr_f_reg_3(.CP(n_63052), .D(n_8607), .CD(n_62318), .Q(iDaddr_f
		[3]));
	notech_mux2 i_9612(.S(n_948), .A(iDaddr[3]), .B(iDaddr_f[3]), .Z(n_8607)
		);
	notech_and2 i_969(.A(fsm[1]), .B(n_12000), .Z(n_988));
	notech_reg iDaddr_f_reg_4(.CP(n_63052), .D(n_8613), .CD(n_62318), .Q(iDaddr_f
		[4]));
	notech_mux2 i_9620(.S(n_948), .A(iDaddr[4]), .B(iDaddr_f[4]), .Z(n_8613)
		);
	notech_nao3 i_89(.A(n_988), .B(n_12001), .C(fsm[0]), .Z(n_989));
	notech_reg iDaddr_f_reg_5(.CP(n_63052), .D(n_8619), .CD(n_62318), .Q(iDaddr_f
		[5]));
	notech_mux2 i_9628(.S(n_948), .A(iDaddr[5]), .B(iDaddr_f[5]), .Z(n_8619)
		);
	notech_nand3 i_10(.A(n_988), .B(data_miss[0]), .C(n_11847), .Z(n_990));
	notech_reg iDaddr_f_reg_6(.CP(n_63052), .D(n_8625), .CD(n_62318), .Q(iDaddr_f
		[6]));
	notech_mux2 i_9636(.S(n_948), .A(iDaddr[6]), .B(iDaddr_f[6]), .Z(n_8625)
		);
	notech_reg iDaddr_f_reg_7(.CP(n_63057), .D(n_8631), .CD(n_62323), .Q(iDaddr_f
		[7]));
	notech_mux2 i_9644(.S(n_948), .A(iDaddr[7]), .B(iDaddr_f[7]), .Z(n_8631)
		);
	notech_or4 i_72(.A(fsm[0]), .B(n_984), .C(fsm[3]), .D(n_12166), .Z(n_992
		));
	notech_reg iDaddr_f_reg_8(.CP(n_63056), .D(n_8637), .CD(n_62322), .Q(iDaddr_f
		[8]));
	notech_mux2 i_9652(.S(n_948), .A(iDaddr[8]), .B(iDaddr_f[8]), .Z(n_8637)
		);
	notech_reg iDaddr_f_reg_9(.CP(n_63057), .D(n_8643), .CD(n_62323), .Q(iDaddr_f
		[9]));
	notech_mux2 i_9660(.S(n_948), .A(iDaddr[9]), .B(iDaddr_f[9]), .Z(n_8643)
		);
	notech_reg iDaddr_f_reg_10(.CP(n_63057), .D(n_8649), .CD(n_62323), .Q(iDaddr_f
		[10]));
	notech_mux2 i_9668(.S(n_948), .A(iDaddr[10]), .B(iDaddr_f[10]), .Z(n_8649
		));
	notech_and2 i_966(.A(fsm[2]), .B(n_11998), .Z(n_995));
	notech_reg iDaddr_f_reg_11(.CP(n_63056), .D(n_8655), .CD(n_62322), .Q(iDaddr_f
		[11]));
	notech_mux2 i_9676(.S(n_948), .A(iDaddr[11]), .B(iDaddr_f[11]), .Z(n_8655
		));
	notech_nao3 i_88(.A(n_995), .B(n_12001), .C(fsm[0]), .Z(n_996));
	notech_reg iDaddr_f_reg_12(.CP(n_63056), .D(\tab11_0[0] ), .CD(n_62322),
		 .Q(iDaddr_f[12]));
	notech_reg iDaddr_f_reg_13(.CP(n_63056), .D(\tab11_0[1] ), .CD(n_62322),
		 .Q(iDaddr_f[13]));
	notech_reg iDaddr_f_reg_14(.CP(n_63056), .D(\tab11_0[2] ), .CD(n_62322),
		 .Q(iDaddr_f[14]));
	notech_nand2 i_78736(.A(data_miss[0]), .B(n_605), .Z(n_999));
	notech_reg iDaddr_f_reg_15(.CP(n_63056), .D(\tab11_0[3] ), .CD(n_62322),
		 .Q(iDaddr_f[15]));
	notech_nand3 i_961(.A(n_995), .B(n_11847), .C(n_11845), .Z(n_1000));
	notech_reg iDaddr_f_reg_16(.CP(n_63051), .D(\tab11_0[4] ), .CD(n_62317),
		 .Q(iDaddr_f[16]));
	notech_nao3 i_17(.A(iread_ack), .B(n_62899), .C(n_1000), .Z(n_1001));
	notech_reg iDaddr_f_reg_17(.CP(n_63051), .D(\tab11_0[5] ), .CD(n_62317),
		 .Q(iDaddr_f[17]));
	notech_nand2 i_98(.A(hit_dir2), .B(n_12164), .Z(n_1002));
	notech_reg iDaddr_f_reg_18(.CP(n_63051), .D(\tab11_0[6] ), .CD(n_62317),
		 .Q(iDaddr_f[18]));
	notech_or4 i_12(.A(n_1000), .B(n_1002), .C(n_12167), .D(n_12166), .Z(n_1003
		));
	notech_reg iDaddr_f_reg_19(.CP(n_63051), .D(\tab11_0[7] ), .CD(n_62317),
		 .Q(iDaddr_f[19]));
	notech_reg iDaddr_f_reg_20(.CP(n_63051), .D(\tab11_0[8] ), .CD(n_62317),
		 .Q(iDaddr_f[20]));
	notech_or2 i_958(.A(busy_ram), .B(flush_tlb), .Z(n_1005));
	notech_reg iDaddr_f_reg_21(.CP(n_63051), .D(\tab11_0[9] ), .CD(n_62317),
		 .Q(iDaddr_f[21]));
	notech_or4 i_959(.A(pg_fault), .B(n_1005), .C(n_654), .D(n_652), .Z(n_1006
		));
	notech_reg iDaddr_f_reg_22(.CP(n_63051), .D(\dir1_0[0] ), .CD(n_62317), 
		.Q(iDaddr_f[22]));
	notech_nor2 i_6(.A(hit_dir2), .B(\hit_dir1[7] ), .Z(n_1007));
	notech_reg iDaddr_f_reg_23(.CP(n_63051), .D(\dir1_0[1] ), .CD(n_62317), 
		.Q(iDaddr_f[23]));
	notech_reg iDaddr_f_reg_24(.CP(n_63051), .D(\dir1_0[2] ), .CD(n_62317), 
		.Q(iDaddr_f[24]));
	notech_reg iDaddr_f_reg_25(.CP(n_63052), .D(\dir1_0[3] ), .CD(n_62318), 
		.Q(iDaddr_f[25]));
	notech_or2 i_97(.A(hit_dir2), .B(n_12164), .Z(n_1010));
	notech_reg iDaddr_f_reg_26(.CP(n_63052), .D(\dir1_0[4] ), .CD(n_62318), 
		.Q(iDaddr_f[26]));
	notech_or4 i_13(.A(n_1000), .B(n_1010), .C(n_12167), .D(n_12166), .Z(n_1011
		));
	notech_reg iDaddr_f_reg_27(.CP(n_63052), .D(\dir1_0[5] ), .CD(n_62318), 
		.Q(iDaddr_f[27]));
	notech_reg iDaddr_f_reg_28(.CP(n_63052), .D(\dir1_0[6] ), .CD(n_62318), 
		.Q(iDaddr_f[28]));
	notech_reg iDaddr_f_reg_29(.CP(n_63052), .D(\dir1_0[7] ), .CD(n_62318), 
		.Q(iDaddr_f[29]));
	notech_reg iDaddr_f_reg_30(.CP(n_63051), .D(\dir1_0[8] ), .CD(n_62317), 
		.Q(iDaddr_f[30]));
	notech_nand2 i_78(.A(fsm[0]), .B(n_12001), .Z(n_1015));
	notech_reg iDaddr_f_reg_31(.CP(n_63051), .D(\dir1_0[9] ), .CD(n_62317), 
		.Q(iDaddr_f[31]));
	notech_nao3 i_78790(.A(fsm[1]), .B(n_11846), .C(fsm[2]), .Z(n_1016));
	notech_reg_set dir1_reg_0(.CP(n_63052), .D(n_8781), .SD(n_62318), .Q(\dir1[0] 
		));
	notech_mux2 i_9844(.S(\nbus_14516[0] ), .A(\dir1[0] ), .B(n_59751), .Z(n_8781
		));
	notech_nao3 i_71(.A(n_988), .B(n_11846), .C(hit_adr11), .Z(n_1017));
	notech_reg_set dir1_reg_1(.CP(n_63052), .D(n_8787), .SD(n_62318), .Q(\dir1[1] 
		));
	notech_mux2 i_9852(.S(\nbus_14516[0] ), .A(\dir1[1] ), .B(n_59757), .Z(n_8787
		));
	notech_nor2 i_16(.A(hit_adr13), .B(hit_adr14), .Z(n_1018));
	notech_reg_set dir1_reg_2(.CP(n_63057), .D(n_8793), .SD(n_62323), .Q(\dir1[2] 
		));
	notech_mux2 i_9860(.S(\nbus_14516[0] ), .A(\dir1[2] ), .B(n_59763), .Z(n_8793
		));
	notech_nand2 i_131(.A(n_1018), .B(n_11894), .Z(n_1019));
	notech_reg_set dir1_reg_3(.CP(n_63060), .D(n_8799), .SD(n_62326), .Q(\dir1[3] 
		));
	notech_mux2 i_9868(.S(\nbus_14516[0] ), .A(\dir1[3] ), .B(n_59769), .Z(n_8799
		));
	notech_nand3 i_9(.A(n_988), .B(n_11846), .C(n_62899), .Z(n_1020));
	notech_reg dir1_reg_4(.CP(n_63060), .D(n_8805), .CD(n_62326), .Q(\dir1[4] 
		));
	notech_mux2 i_9876(.S(\nbus_14516[0] ), .A(\dir1[4] ), .B(n_976), .Z(n_8805
		));
	notech_reg_set dir1_reg_5(.CP(n_63060), .D(n_8811), .SD(n_62326), .Q(\dir1[5] 
		));
	notech_mux2 i_9884(.S(\nbus_14516[0] ), .A(\dir1[5] ), .B(n_59781), .Z(n_8811
		));
	notech_reg_set dir1_reg_6(.CP(n_63060), .D(n_8817), .SD(n_62326), .Q(\dir1[6] 
		));
	notech_mux2 i_9892(.S(\nbus_14516[0] ), .A(\dir1[6] ), .B(n_59787), .Z(n_8817
		));
	notech_reg_set dir1_reg_7(.CP(n_63060), .D(n_8823), .SD(n_62326), .Q(\dir1[7] 
		));
	notech_mux2 i_9900(.S(\nbus_14516[0] ), .A(\dir1[7] ), .B(n_59793), .Z(n_8823
		));
	notech_nor2 i_31(.A(hit_adr23), .B(hit_adr24), .Z(n_1024));
	notech_reg_set dir1_reg_8(.CP(n_63060), .D(n_8829), .SD(n_62326), .Q(\dir1[8] 
		));
	notech_mux2 i_9908(.S(\nbus_14516[0] ), .A(\dir1[8] ), .B(n_59799), .Z(n_8829
		));
	notech_nand2 i_132(.A(n_1024), .B(n_11946), .Z(n_1025));
	notech_reg_set dir1_reg_9(.CP(n_63060), .D(n_8835), .SD(n_62326), .Q(\dir1[9] 
		));
	notech_mux2 i_9916(.S(\nbus_14516[0] ), .A(\dir1[9] ), .B(n_59805), .Z(n_8835
		));
	notech_nao3 i_73(.A(n_988), .B(n_11846), .C(hit_adr21), .Z(n_1026));
	notech_reg_set dir1_reg_10(.CP(n_63060), .D(n_8841), .SD(n_62326), .Q(\dir1[10] 
		));
	notech_mux2 i_9924(.S(\nbus_14516[0] ), .A(\dir1[10] ), .B(n_59811), .Z(n_8841
		));
	notech_reg_set dir1_reg_11(.CP(n_63060), .D(n_8847), .SD(n_62326), .Q(\dir1[11] 
		));
	notech_mux2 i_9932(.S(\nbus_14516[0] ), .A(\dir1[11] ), .B(n_59817), .Z(n_8847
		));
	notech_nao3 i_78797(.A(fsm[2]), .B(n_11846), .C(fsm[1]), .Z(n_1028));
	notech_reg_set dir1_reg_12(.CP(n_63061), .D(n_8853), .SD(n_62327), .Q(\dir1[12] 
		));
	notech_mux2 i_9940(.S(\nbus_14516[0] ), .A(\dir1[12] ), .B(n_59823), .Z(n_8853
		));
	notech_reg_set dir1_reg_13(.CP(n_63061), .D(n_8859), .SD(n_62327), .Q(\dir1[13] 
		));
	notech_mux2 i_9948(.S(\nbus_14516[0] ), .A(\dir1[13] ), .B(n_59829), .Z(n_8859
		));
	notech_or2 i_50(.A(n_553), .B(fsm5_cnt[8]), .Z(n_1030));
	notech_reg_set dir1_reg_14(.CP(n_63061), .D(n_8865), .SD(n_62327), .Q(\dir1[14] 
		));
	notech_mux2 i_9956(.S(\nbus_14516[0] ), .A(\dir1[14] ), .B(n_59835), .Z(n_8865
		));
	notech_reg_set dir1_reg_15(.CP(n_63061), .D(n_8871), .SD(n_62327), .Q(\dir1[15] 
		));
	notech_mux2 i_9964(.S(\nbus_14516[0] ), .A(\dir1[15] ), .B(n_59841), .Z(n_8871
		));
	notech_nand2 i_69(.A(fsm[2]), .B(fsm[1]), .Z(n_1032));
	notech_reg_set dir1_reg_16(.CP(n_63061), .D(n_8877), .SD(n_62327), .Q(\dir1[16] 
		));
	notech_mux2 i_9972(.S(n_56110), .A(\dir1[16] ), .B(n_59847), .Z(n_8877)
		);
	notech_ao4 i_932(.A(n_990), .B(data_miss[5]), .C(iwrite_ack), .D(n_1032)
		, .Z(n_1033));
	notech_reg_set dir1_reg_17(.CP(n_63060), .D(n_8883), .SD(n_62326), .Q(\dir1[17] 
		));
	notech_mux2 i_9980(.S(n_56110), .A(\dir1[17] ), .B(n_59853), .Z(n_8883)
		);
	notech_reg_set dir1_reg_18(.CP(n_63060), .D(n_8889), .SD(n_62326), .Q(\dir1[18] 
		));
	notech_mux2 i_9988(.S(n_56110), .A(\dir1[18] ), .B(n_59859), .Z(n_8889)
		);
	notech_nand2 i_95(.A(n_549), .B(n_56853), .Z(n_1035));
	notech_reg_set dir1_reg_19(.CP(n_63061), .D(n_8895), .SD(n_62327), .Q(\dir1[19] 
		));
	notech_mux2 i_9996(.S(n_56110), .A(\dir1[19] ), .B(n_59865), .Z(n_8895)
		);
	notech_reg_set dir1_reg_20(.CP(n_63061), .D(n_8901), .SD(n_62327), .Q(\dir1[20] 
		));
	notech_mux2 i_10004(.S(n_56110), .A(\dir1[20] ), .B(n_59871), .Z(n_8901)
		);
	notech_reg_set dir1_reg_21(.CP(n_63057), .D(n_8907), .SD(n_62323), .Q(\dir1[21] 
		));
	notech_mux2 i_10012(.S(n_56110), .A(\dir1[21] ), .B(n_59877), .Z(n_8907)
		);
	notech_ao4 i_927(.A(n_546), .B(iwrite_ack), .C(n_550), .D(n_1000), .Z(n_1038
		));
	notech_reg_set dir1_reg_22(.CP(n_63057), .D(n_8913), .SD(n_62323), .Q(\dir1[22] 
		));
	notech_mux2 i_10020(.S(n_56110), .A(\dir1[22] ), .B(n_59883), .Z(n_8913)
		);
	notech_reg_set dir1_reg_23(.CP(n_63058), .D(n_8919), .SD(n_62324), .Q(\dir1[23] 
		));
	notech_mux2 i_10028(.S(n_56110), .A(\dir1[23] ), .B(n_59889), .Z(n_8919)
		);
	notech_nao3 i_78783(.A(fsm[0]), .B(n_12001), .C(n_984), .Z(n_1040));
	notech_reg_set dir1_reg_24(.CP(n_63058), .D(n_8925), .SD(n_62324), .Q(\dir1[24] 
		));
	notech_mux2 i_10036(.S(n_56110), .A(\dir1[24] ), .B(n_59895), .Z(n_8925)
		);
	notech_reg_set dir1_reg_25(.CP(n_63057), .D(n_8931), .SD(n_62323), .Q(\dir1[25] 
		));
	notech_mux2 i_10044(.S(n_56110), .A(\dir1[25] ), .B(n_59901), .Z(n_8931)
		);
	notech_nand3 i_81(.A(fsm[2]), .B(fsm[1]), .C(n_12001), .Z(n_1042));
	notech_reg_set dir1_reg_26(.CP(n_63057), .D(n_8937), .SD(n_62323), .Q(\dir1[26] 
		));
	notech_mux2 i_10052(.S(n_56110), .A(\dir1[26] ), .B(n_59907), .Z(n_8937)
		);
	notech_or4 i_14(.A(n_12000), .B(n_11998), .C(fsm[3]), .D(n_12166), .Z(n_1043
		));
	notech_reg_set dir1_reg_27(.CP(n_63057), .D(n_8943), .SD(n_62323), .Q(\dir1[27] 
		));
	notech_mux2 i_10060(.S(n_56110), .A(\dir1[27] ), .B(n_59913), .Z(n_8943)
		);
	notech_reg_set dir1_reg_28(.CP(n_63057), .D(n_8949), .SD(n_62323), .Q(\dir1[28] 
		));
	notech_mux2 i_10068(.S(n_56110), .A(\dir1[28] ), .B(n_59919), .Z(n_8949)
		);
	notech_reg_set dir1_reg_29(.CP(n_63057), .D(n_8955), .SD(n_62323), .Q(\dir1[29] 
		));
	notech_mux2 i_10076(.S(n_56110), .A(\dir1[29] ), .B(n_59925), .Z(n_8955)
		);
	notech_reg_set dir1_reg_33(.CP(n_63058), .D(n_8961), .SD(n_62324), .Q(\dir1[33] 
		));
	notech_mux2 i_10084(.S(n_56110), .A(\dir1[33] ), .B(n_11870), .Z(n_8961)
		);
	notech_reg_set dir2_reg_0(.CP(n_63058), .D(n_8967), .SD(n_62324), .Q(\dir2[0] 
		));
	notech_mux2 i_10092(.S(\nbus_14517[0] ), .A(\dir2[0] ), .B(n_59751), .Z(n_8967
		));
	notech_nand3 i_921(.A(n_952), .B(n_1043), .C(n_953), .Z(n_1048));
	notech_reg_set dir2_reg_1(.CP(n_63058), .D(n_8973), .SD(n_62324), .Q(\dir2[1] 
		));
	notech_mux2 i_10100(.S(\nbus_14517[0] ), .A(\dir2[1] ), .B(n_59757), .Z(n_8973
		));
	notech_reg_set dir2_reg_2(.CP(n_63058), .D(n_8979), .SD(n_62324), .Q(\dir2[2] 
		));
	notech_mux2 i_10108(.S(\nbus_14517[0] ), .A(\dir2[2] ), .B(n_59763), .Z(n_8979
		));
	notech_ao4 i_917(.A(n_1032), .B(n_1015), .C(n_541), .D(n_12001), .Z(n_1050
		));
	notech_reg_set dir2_reg_3(.CP(n_63058), .D(n_8985), .SD(n_62324), .Q(\dir2[3] 
		));
	notech_mux2 i_10116(.S(\nbus_14517[0] ), .A(\dir2[3] ), .B(n_59769), .Z(n_8985
		));
	notech_reg dir2_reg_4(.CP(n_63058), .D(n_8991), .CD(n_62324), .Q(\dir2[4] 
		));
	notech_mux2 i_10124(.S(\nbus_14517[0] ), .A(\dir2[4] ), .B(n_976), .Z(n_8991
		));
	notech_reg_set dir2_reg_5(.CP(n_63058), .D(n_8997), .SD(n_62324), .Q(\dir2[5] 
		));
	notech_mux2 i_10132(.S(\nbus_14517[0] ), .A(\dir2[5] ), .B(n_59781), .Z(n_8997
		));
	notech_nand2 i_44(.A(n_62893), .B(n_55416), .Z(n_1053));
	notech_reg_set dir2_reg_6(.CP(n_63058), .D(n_9003), .SD(n_62324), .Q(\dir2[6] 
		));
	notech_mux2 i_10140(.S(\nbus_14517[0] ), .A(\dir2[6] ), .B(n_59787), .Z(n_9003
		));
	notech_reg_set dir2_reg_7(.CP(n_63058), .D(n_9009), .SD(n_62324), .Q(\dir2[7] 
		));
	notech_mux2 i_10148(.S(\nbus_14517[0] ), .A(\dir2[7] ), .B(n_59793), .Z(n_9009
		));
	notech_ao3 i_21(.A(n_988), .B(n_11846), .C(\hit_dir1[7] ), .Z(n_1055));
	notech_reg_set dir2_reg_8(.CP(n_63050), .D(n_9015), .SD(n_62316), .Q(\dir2[8] 
		));
	notech_mux2 i_10156(.S(\nbus_14517[0] ), .A(\dir2[8] ), .B(n_59799), .Z(n_9015
		));
	notech_nand3 i_29(.A(n_988), .B(\hit_dir1[7] ), .C(n_11846), .Z(n_1056)
		);
	notech_reg_set dir2_reg_9(.CP(n_63043), .D(n_9021), .SD(n_62309), .Q(\dir2[9] 
		));
	notech_mux2 i_10164(.S(\nbus_14517[0] ), .A(\dir2[9] ), .B(n_59805), .Z(n_9021
		));
	notech_ao4 i_913(.A(n_1056), .B(n_11869), .C(n_1040), .D(n_12086), .Z(n_1057
		));
	notech_reg_set dir2_reg_10(.CP(n_63043), .D(n_9027), .SD(n_62309), .Q(\dir2[10] 
		));
	notech_mux2 i_10172(.S(\nbus_14517[0] ), .A(\dir2[10] ), .B(n_59811), .Z
		(n_9027));
	notech_ao4 i_912(.A(n_1056), .B(n_11868), .C(n_1040), .D(n_12087), .Z(n_1058
		));
	notech_reg_set dir2_reg_11(.CP(n_63043), .D(n_9033), .SD(n_62309), .Q(\dir2[11] 
		));
	notech_mux2 i_10180(.S(\nbus_14517[0] ), .A(\dir2[11] ), .B(n_59817), .Z
		(n_9033));
	notech_ao4 i_911(.A(n_1056), .B(n_11867), .C(n_1040), .D(n_12088), .Z(n_1059
		));
	notech_reg_set dir2_reg_12(.CP(n_63043), .D(n_9039), .SD(n_62309), .Q(\dir2[12] 
		));
	notech_mux2 i_10188(.S(\nbus_14517[0] ), .A(\dir2[12] ), .B(n_59823), .Z
		(n_9039));
	notech_ao4 i_910(.A(n_1056), .B(n_11865), .C(n_1040), .D(n_12089), .Z(n_1060
		));
	notech_reg_set dir2_reg_13(.CP(n_63043), .D(n_9045), .SD(n_62309), .Q(\dir2[13] 
		));
	notech_mux2 i_10196(.S(\nbus_14517[0] ), .A(\dir2[13] ), .B(n_59829), .Z
		(n_9045));
	notech_ao4 i_909(.A(n_1056), .B(n_11864), .C(n_1040), .D(n_12090), .Z(n_1061
		));
	notech_reg_set dir2_reg_14(.CP(n_63043), .D(n_9051), .SD(n_62309), .Q(\dir2[14] 
		));
	notech_mux2 i_10204(.S(\nbus_14517[0] ), .A(\dir2[14] ), .B(n_59835), .Z
		(n_9051));
	notech_ao4 i_908(.A(n_1056), .B(n_11863), .C(n_1040), .D(n_12091), .Z(n_1062
		));
	notech_reg_set dir2_reg_15(.CP(n_63042), .D(n_9057), .SD(n_62308), .Q(\dir2[15] 
		));
	notech_mux2 i_10212(.S(\nbus_14517[0] ), .A(\dir2[15] ), .B(n_59841), .Z
		(n_9057));
	notech_ao4 i_907(.A(n_1056), .B(n_11862), .C(n_1040), .D(n_12092), .Z(n_1063
		));
	notech_reg_set dir2_reg_16(.CP(n_63043), .D(n_9063), .SD(n_62309), .Q(\dir2[16] 
		));
	notech_mux2 i_10220(.S(n_56177), .A(\dir2[16] ), .B(n_59847), .Z(n_9063)
		);
	notech_ao4 i_906(.A(n_1056), .B(n_11861), .C(n_1040), .D(n_12093), .Z(n_1064
		));
	notech_reg_set dir2_reg_17(.CP(n_63043), .D(n_9069), .SD(n_62309), .Q(\dir2[17] 
		));
	notech_mux2 i_10228(.S(n_56177), .A(\dir2[17] ), .B(n_59853), .Z(n_9069)
		);
	notech_ao4 i_905(.A(n_1056), .B(n_11860), .C(n_1040), .D(n_12094), .Z(n_1065
		));
	notech_reg_set dir2_reg_18(.CP(n_63046), .D(n_9075), .SD(n_62312), .Q(\dir2[18] 
		));
	notech_mux2 i_10236(.S(n_56177), .A(\dir2[18] ), .B(n_59859), .Z(n_9075)
		);
	notech_ao4 i_904(.A(n_1056), .B(n_11859), .C(n_1040), .D(n_12095), .Z(n_1066
		));
	notech_reg_set dir2_reg_19(.CP(n_63046), .D(n_9081), .SD(n_62312), .Q(\dir2[19] 
		));
	notech_mux2 i_10244(.S(n_56177), .A(\dir2[19] ), .B(n_59865), .Z(n_9081)
		);
	notech_ao4 i_903(.A(n_1056), .B(n_11858), .C(n_1040), .D(n_12096), .Z(n_1067
		));
	notech_reg_set dir2_reg_20(.CP(n_63046), .D(n_9087), .SD(n_62312), .Q(\dir2[20] 
		));
	notech_mux2 i_10252(.S(n_56177), .A(\dir2[20] ), .B(n_59871), .Z(n_9087)
		);
	notech_ao4 i_902(.A(n_1056), .B(n_11857), .C(n_1040), .D(n_12097), .Z(n_1068
		));
	notech_reg_set dir2_reg_21(.CP(n_63046), .D(n_9093), .SD(n_62312), .Q(\dir2[21] 
		));
	notech_mux2 i_10260(.S(n_56177), .A(\dir2[21] ), .B(n_59877), .Z(n_9093)
		);
	notech_ao4 i_901(.A(n_1056), .B(n_11856), .C(n_1040), .D(n_12098), .Z(n_1069
		));
	notech_reg_set dir2_reg_22(.CP(n_63046), .D(n_9099), .SD(n_62312), .Q(\dir2[22] 
		));
	notech_mux2 i_10268(.S(n_56177), .A(\dir2[22] ), .B(n_59883), .Z(n_9099)
		);
	notech_ao4 i_900(.A(n_1056), .B(n_11855), .C(n_1040), .D(n_12099), .Z(n_1070
		));
	notech_reg_set dir2_reg_23(.CP(n_63043), .D(n_9105), .SD(n_62309), .Q(\dir2[23] 
		));
	notech_mux2 i_10276(.S(n_56177), .A(\dir2[23] ), .B(n_59889), .Z(n_9105)
		);
	notech_ao4 i_899(.A(n_1056), .B(n_11854), .C(n_1040), .D(n_12100), .Z(n_1071
		));
	notech_reg_set dir2_reg_24(.CP(n_63043), .D(n_9111), .SD(n_62309), .Q(\dir2[24] 
		));
	notech_mux2 i_10284(.S(n_56177), .A(\dir2[24] ), .B(n_59895), .Z(n_9111)
		);
	notech_ao4 i_898(.A(n_1056), .B(n_11853), .C(n_1040), .D(n_12101), .Z(n_1072
		));
	notech_reg_set dir2_reg_25(.CP(n_63046), .D(n_9117), .SD(n_62312), .Q(\dir2[25] 
		));
	notech_mux2 i_10292(.S(n_56177), .A(\dir2[25] ), .B(n_59901), .Z(n_9117)
		);
	notech_ao4 i_897(.A(n_1056), .B(n_11852), .C(n_56290), .D(n_12102), .Z(n_1073
		));
	notech_reg_set dir2_reg_26(.CP(n_63043), .D(n_9123), .SD(n_62309), .Q(\dir2[26] 
		));
	notech_mux2 i_10300(.S(n_56177), .A(\dir2[26] ), .B(n_59907), .Z(n_9123)
		);
	notech_ao4 i_896(.A(n_1056), .B(n_11851), .C(n_56290), .D(n_12103), .Z(n_1074
		));
	notech_reg_set dir2_reg_27(.CP(n_63041), .D(n_9129), .SD(n_62307), .Q(\dir2[27] 
		));
	notech_mux2 i_10308(.S(n_56177), .A(\dir2[27] ), .B(n_59913), .Z(n_9129)
		);
	notech_ao4 i_895(.A(n_1056), .B(n_11850), .C(n_56290), .D(n_12104), .Z(n_1075
		));
	notech_reg_set dir2_reg_28(.CP(n_63041), .D(n_9135), .SD(n_62307), .Q(\dir2[28] 
		));
	notech_mux2 i_10316(.S(n_56177), .A(\dir2[28] ), .B(n_59919), .Z(n_9135)
		);
	notech_ao4 i_894(.A(n_1056), .B(n_11849), .C(n_56290), .D(n_12105), .Z(n_1076
		));
	notech_reg_set dir2_reg_29(.CP(n_63042), .D(n_9141), .SD(n_62308), .Q(\dir2[29] 
		));
	notech_mux2 i_10324(.S(n_56177), .A(\dir2[29] ), .B(n_59925), .Z(n_9141)
		);
	notech_nand2 i_83(.A(n_406), .B(n_12012), .Z(n_1077));
	notech_reg_set dir2_reg_33(.CP(n_63041), .D(n_9147), .SD(n_62307), .Q(\dir2[33] 
		));
	notech_mux2 i_10332(.S(n_56177), .A(\dir2[33] ), .B(n_11870), .Z(n_9147)
		);
	notech_reg_set tab21_reg_0(.CP(n_63041), .D(n_9153), .SD(n_62307), .Q(\tab21[0] 
		));
	notech_mux2 i_10340(.S(\nbus_14511[0] ), .A(\tab21[0] ), .B(n_56627), .Z
		(n_9153));
	notech_reg_set tab21_reg_1(.CP(n_63041), .D(n_9159), .SD(n_62307), .Q(\tab21[1] 
		));
	notech_mux2 i_10348(.S(\nbus_14511[0] ), .A(\tab21[1] ), .B(n_56633), .Z
		(n_9159));
	notech_nand3 i_1(.A(n_62893), .B(n_55416), .C(n_983), .Z(n_1080));
	notech_reg_set tab21_reg_2(.CP(n_63041), .D(n_9165), .SD(n_62307), .Q(\tab21[2] 
		));
	notech_mux2 i_10356(.S(\nbus_14511[0] ), .A(\tab21[2] ), .B(n_56639), .Z
		(n_9165));
	notech_or4 i_77(.A(\hit_dir1[7] ), .B(n_12166), .C(n_11843), .D(n_11848)
		, .Z(n_1081));
	notech_reg_set tab21_reg_3(.CP(n_63041), .D(n_9171), .SD(n_62307), .Q(\tab21[3] 
		));
	notech_mux2 i_10364(.S(\nbus_14511[0] ), .A(\tab21[3] ), .B(n_56645), .Z
		(n_9171));
	notech_reg tab21_reg_4(.CP(n_63041), .D(n_9177), .CD(n_62307), .Q(\tab21[4] 
		));
	notech_mux2 i_10372(.S(\nbus_14511[0] ), .A(\tab21[4] ), .B(n_973), .Z(n_9177
		));
	notech_reg_set tab21_reg_5(.CP(n_63042), .D(n_9183), .SD(n_62308), .Q(\tab21[5] 
		));
	notech_mux2 i_10380(.S(\nbus_14511[0] ), .A(\tab21[5] ), .B(n_56657), .Z
		(n_9183));
	notech_nao3 i_27(.A(hit_tab22), .B(n_12165), .C(n_55384), .Z(n_1084));
	notech_reg_set tab21_reg_6(.CP(n_63042), .D(n_9189), .SD(n_62308), .Q(\tab21[6] 
		));
	notech_mux2 i_10388(.S(\nbus_14511[0] ), .A(\tab21[6] ), .B(n_56663), .Z
		(n_9189));
	notech_nao3 i_75(.A(\hit_dir1[7] ), .B(n_983), .C(n_1053), .Z(n_1085));
	notech_reg_set tab21_reg_7(.CP(n_63042), .D(n_9195), .SD(n_62308), .Q(\tab21[7] 
		));
	notech_mux2 i_10396(.S(\nbus_14511[0] ), .A(\tab21[7] ), .B(n_56669), .Z
		(n_9195));
	notech_or4 i_30(.A(hit_tab12), .B(n_58725), .C(hit_tab13), .D(n_1085), .Z
		(n_1086));
	notech_reg_set tab21_reg_8(.CP(n_63042), .D(n_9201), .SD(n_62308), .Q(\tab21[8] 
		));
	notech_mux2 i_10404(.S(\nbus_14511[0] ), .A(\tab21[8] ), .B(n_56675), .Z
		(n_9201));
	notech_ao4 i_883(.A(n_1086), .B(n_11916), .C(n_1084), .D(n_11945), .Z(n_1087
		));
	notech_reg_set tab21_reg_9(.CP(n_63042), .D(n_9207), .SD(n_62308), .Q(\tab21[9] 
		));
	notech_mux2 i_10412(.S(\nbus_14511[0] ), .A(\tab21[9] ), .B(n_56681), .Z
		(n_9207));
	notech_reg_set tab21_reg_10(.CP(n_63042), .D(n_9213), .SD(n_62308), .Q(\tab21[10] 
		));
	notech_mux2 i_10420(.S(\nbus_14511[0] ), .A(\tab21[10] ), .B(n_56687), .Z
		(n_9213));
	notech_reg_set tab21_reg_11(.CP(n_63042), .D(n_9219), .SD(n_62308), .Q(\tab21[11] 
		));
	notech_mux2 i_10428(.S(\nbus_14511[0] ), .A(\tab21[11] ), .B(n_56693), .Z
		(n_9219));
	notech_or4 i_24(.A(hit_tab22), .B(n_58734), .C(n_55384), .D(hit_tab23), 
		.Z(n_1090));
	notech_reg_set tab21_reg_12(.CP(n_63042), .D(n_9225), .SD(n_62308), .Q(\tab21[12] 
		));
	notech_mux2 i_10436(.S(\nbus_14511[0] ), .A(\tab21[12] ), .B(n_56699), .Z
		(n_9225));
	notech_reg_set tab21_reg_13(.CP(n_63042), .D(n_9231), .SD(n_62308), .Q(\tab21[13] 
		));
	notech_mux2 i_10444(.S(\nbus_14511[0] ), .A(\tab21[13] ), .B(n_56705), .Z
		(n_9231));
	notech_or4 i_26(.A(hit_tab22), .B(n_58734), .C(n_55384), .D(n_12163), .Z
		(n_1092));
	notech_reg_set tab21_reg_14(.CP(n_63046), .D(n_9237), .SD(n_62312), .Q(\tab21[14] 
		));
	notech_mux2 i_10452(.S(\nbus_14511[0] ), .A(\tab21[14] ), .B(n_56711), .Z
		(n_9237));
	notech_ao4 i_881(.A(n_1092), .B(n_11966), .C(n_1090), .D(n_11986), .Z(n_1093
		));
	notech_reg_set tab21_reg_15(.CP(n_63048), .D(n_9243), .SD(n_62314), .Q(\tab21[15] 
		));
	notech_mux2 i_10460(.S(\nbus_14511[0] ), .A(\tab21[15] ), .B(n_56717), .Z
		(n_9243));
	notech_reg_set tab21_reg_16(.CP(n_63048), .D(n_9249), .SD(n_62314), .Q(\tab21[16] 
		));
	notech_mux2 i_10468(.S(\nbus_14511[0] ), .A(\tab21[16] ), .B(n_56723), .Z
		(n_9249));
	notech_and4 i_885(.A(n_1093), .B(n_1087), .C(n_897), .D(n_900), .Z(n_1095
		));
	notech_reg_set tab21_reg_17(.CP(n_63050), .D(n_9255), .SD(n_62316), .Q(\tab21[17] 
		));
	notech_mux2 i_10476(.S(n_56130), .A(\tab21[17] ), .B(n_56729), .Z(n_9255
		));
	notech_ao3 i_886(.A(hit_tab13), .B(n_12162), .C(n_58725), .Z(n_1096));
	notech_reg_set tab21_reg_18(.CP(n_63048), .D(n_9261), .SD(n_62314), .Q(\tab21[18] 
		));
	notech_mux2 i_10484(.S(n_56130), .A(\tab21[18] ), .B(n_56735), .Z(n_9261
		));
	notech_reg_set tab21_reg_19(.CP(n_63048), .D(n_9267), .SD(n_62314), .Q(\tab21[19] 
		));
	notech_mux2 i_10492(.S(n_56130), .A(\tab21[19] ), .B(n_56741), .Z(n_9267
		));
	notech_or4 i_15(.A(n_654), .B(n_652), .C(n_12166), .D(n_11843), .Z(n_1098
		));
	notech_reg_set tab21_reg_20(.CP(n_63048), .D(n_9273), .SD(n_62314), .Q(\tab21[20] 
		));
	notech_mux2 i_10500(.S(n_56130), .A(\tab21[20] ), .B(n_56747), .Z(n_9273
		));
	notech_reg_set tab21_reg_21(.CP(n_63048), .D(n_9279), .SD(n_62314), .Q(\tab21[21] 
		));
	notech_mux2 i_10508(.S(n_56130), .A(\tab21[21] ), .B(n_56753), .Z(n_9279
		));
	notech_nao3 i_23(.A(hit_tab12), .B(n_55406), .C(n_58725), .Z(n_1100));
	notech_reg_set tab21_reg_22(.CP(n_63048), .D(n_9285), .SD(n_62314), .Q(\tab21[22] 
		));
	notech_mux2 i_10516(.S(n_56130), .A(\tab21[22] ), .B(n_56759), .Z(n_9285
		));
	notech_ao4 i_878(.A(n_1100), .B(n_11893), .C(n_1098), .D(n_12063), .Z(n_1101
		));
	notech_reg_set tab21_reg_23(.CP(n_63048), .D(n_9291), .SD(n_62314), .Q(\tab21[23] 
		));
	notech_mux2 i_10524(.S(n_56130), .A(\tab21[23] ), .B(n_56765), .Z(n_9291
		));
	notech_reg_set tab21_reg_24(.CP(n_63050), .D(n_9297), .SD(n_62316), .Q(\tab21[24] 
		));
	notech_mux2 i_10532(.S(n_56130), .A(\tab21[24] ), .B(n_56771), .Z(n_9297
		));
	notech_ao4 i_877(.A(n_62893), .B(n_12137), .C(n_1043), .D(n_12064), .Z(n_1103
		));
	notech_reg_set tab21_reg_25(.CP(n_63050), .D(n_9303), .SD(n_62316), .Q(\tab21[25] 
		));
	notech_mux2 i_10540(.S(n_56130), .A(\tab21[25] ), .B(n_56777), .Z(n_9303
		));
	notech_reg_set tab21_reg_26(.CP(n_63050), .D(n_9309), .SD(n_62316), .Q(\tab21[26] 
		));
	notech_mux2 i_10548(.S(n_56130), .A(\tab21[26] ), .B(n_56783), .Z(n_9309
		));
	notech_ao4 i_874(.A(n_1086), .B(n_11915), .C(n_1084), .D(n_11944), .Z(n_1105
		));
	notech_reg_set tab21_reg_27(.CP(n_63050), .D(n_9315), .SD(n_62316), .Q(\tab21[27] 
		));
	notech_mux2 i_10556(.S(\nbus_14511[0] ), .A(\tab21[27] ), .B(n_56789), .Z
		(n_9315));
	notech_reg_set tab21_reg_28(.CP(n_63050), .D(n_9321), .SD(n_62316), .Q(\tab21[28] 
		));
	notech_mux2 i_10564(.S(n_56130), .A(\tab21[28] ), .B(n_56795), .Z(n_9321
		));
	notech_ao4 i_872(.A(n_1092), .B(n_11965), .C(n_1090), .D(n_11985), .Z(n_1107
		));
	notech_reg_set tab21_reg_29(.CP(n_63050), .D(n_9327), .SD(n_62316), .Q(\tab21[29] 
		));
	notech_mux2 i_10572(.S(n_56130), .A(\tab21[29] ), .B(n_56801), .Z(n_9327
		));
	notech_reg tab21_reg_30(.CP(n_63050), .D(n_9333), .CD(n_62316), .Q(\tab21[30] 
		));
	notech_mux2 i_10580(.S(n_56130), .A(\tab21[30] ), .B(n_974), .Z(n_9333)
		);
	notech_and4 i_876(.A(n_1107), .B(n_1105), .C(n_886), .D(n_889), .Z(n_1109
		));
	notech_reg tab21_reg_32(.CP(n_63050), .D(n_9339), .CD(n_62316), .Q(\tab21[32] 
		));
	notech_mux2 i_10588(.S(n_56130), .A(\tab21[32] ), .B(n_975), .Z(n_9339)
		);
	notech_ao4 i_869(.A(n_1100), .B(n_11892), .C(n_1098), .D(n_12061), .Z(n_1110
		));
	notech_reg_set tab21_reg_33(.CP(n_63050), .D(n_9345), .SD(n_62316), .Q(\tab21[33] 
		));
	notech_mux2 i_10596(.S(n_56130), .A(\tab21[33] ), .B(n_56153), .Z(n_9345
		));
	notech_reg hit_adr11_reg(.CP(n_63047), .D(n_9351), .CD(n_62313), .Q(hit_adr11
		));
	notech_mux2 i_10604(.S(n_971), .A(hit_add11), .B(hit_adr11), .Z(n_9351)
		);
	notech_ao4 i_868(.A(n_62893), .B(n_12136), .C(n_1043), .D(n_12062), .Z(n_1112
		));
	notech_reg_set tab12_reg_0(.CP(n_63047), .D(n_9357), .SD(n_62313), .Q(\tab12[0] 
		));
	notech_mux2 i_10612(.S(\nbus_14508[0] ), .A(\tab12[0] ), .B(n_56627), .Z
		(n_9357));
	notech_reg_set tab12_reg_1(.CP(n_63047), .D(n_9363), .SD(n_62313), .Q(\tab12[1] 
		));
	notech_mux2 i_10620(.S(\nbus_14508[0] ), .A(\tab12[1] ), .B(n_56633), .Z
		(n_9363));
	notech_ao4 i_865(.A(n_1086), .B(n_11914), .C(n_1084), .D(n_11943), .Z(n_1114
		));
	notech_reg_set tab12_reg_2(.CP(n_63047), .D(n_9369), .SD(n_62313), .Q(\tab12[2] 
		));
	notech_mux2 i_10628(.S(\nbus_14508[0] ), .A(\tab12[2] ), .B(n_56639), .Z
		(n_9369));
	notech_reg_set tab12_reg_3(.CP(n_63047), .D(n_9375), .SD(n_62313), .Q(\tab12[3] 
		));
	notech_mux2 i_10636(.S(\nbus_14508[0] ), .A(\tab12[3] ), .B(n_56645), .Z
		(n_9375));
	notech_ao4 i_863(.A(n_1092), .B(n_11964), .C(n_1090), .D(n_11984), .Z(n_1116
		));
	notech_reg tab12_reg_4(.CP(n_63046), .D(n_9381), .CD(n_62312), .Q(\tab12[4] 
		));
	notech_mux2 i_10644(.S(\nbus_14508[0] ), .A(\tab12[4] ), .B(n_973), .Z(n_9381
		));
	notech_reg_set tab12_reg_5(.CP(n_63046), .D(n_9387), .SD(n_62312), .Q(\tab12[5] 
		));
	notech_mux2 i_10652(.S(\nbus_14508[0] ), .A(\tab12[5] ), .B(n_56657), .Z
		(n_9387));
	notech_and4 i_867(.A(n_1116), .B(n_1114), .C(n_875), .D(n_878), .Z(n_1118
		));
	notech_reg_set tab12_reg_6(.CP(n_63046), .D(n_9393), .SD(n_62312), .Q(\tab12[6] 
		));
	notech_mux2 i_10660(.S(\nbus_14508[0] ), .A(\tab12[6] ), .B(n_56663), .Z
		(n_9393));
	notech_ao4 i_860(.A(n_1100), .B(n_11891), .C(n_1098), .D(n_12059), .Z(n_1119
		));
	notech_reg_set tab12_reg_7(.CP(n_63046), .D(n_9399), .SD(n_62312), .Q(\tab12[7] 
		));
	notech_mux2 i_10668(.S(\nbus_14508[0] ), .A(\tab12[7] ), .B(n_56669), .Z
		(n_9399));
	notech_reg_set tab12_reg_8(.CP(n_63048), .D(n_9405), .SD(n_62314), .Q(\tab12[8] 
		));
	notech_mux2 i_10676(.S(\nbus_14508[0] ), .A(\tab12[8] ), .B(n_56675), .Z
		(n_9405));
	notech_ao4 i_859(.A(n_62893), .B(n_12135), .C(n_1043), .D(n_12060), .Z(n_1121
		));
	notech_reg_set tab12_reg_9(.CP(n_63047), .D(n_9411), .SD(n_62313), .Q(\tab12[9] 
		));
	notech_mux2 i_10684(.S(\nbus_14508[0] ), .A(\tab12[9] ), .B(n_56681), .Z
		(n_9411));
	notech_reg_set tab12_reg_10(.CP(n_63048), .D(n_9417), .SD(n_62314), .Q(\tab12[10] 
		));
	notech_mux2 i_10692(.S(\nbus_14508[0] ), .A(\tab12[10] ), .B(n_56687), .Z
		(n_9417));
	notech_ao4 i_856(.A(n_1086), .B(n_11913), .C(n_1084), .D(n_11942), .Z(n_1123
		));
	notech_reg_set tab12_reg_11(.CP(n_63048), .D(n_9423), .SD(n_62314), .Q(\tab12[11] 
		));
	notech_mux2 i_10700(.S(\nbus_14508[0] ), .A(\tab12[11] ), .B(n_56693), .Z
		(n_9423));
	notech_reg_set tab12_reg_12(.CP(n_63047), .D(n_9429), .SD(n_62313), .Q(\tab12[12] 
		));
	notech_mux2 i_10708(.S(\nbus_14508[0] ), .A(\tab12[12] ), .B(n_56699), .Z
		(n_9429));
	notech_ao4 i_854(.A(n_1092), .B(n_11963), .C(n_1090), .D(n_11983), .Z(n_1125
		));
	notech_reg_set tab12_reg_13(.CP(n_63047), .D(n_9435), .SD(n_62313), .Q(\tab12[13] 
		));
	notech_mux2 i_10716(.S(\nbus_14508[0] ), .A(\tab12[13] ), .B(n_56705), .Z
		(n_9435));
	notech_reg_set tab12_reg_14(.CP(n_63047), .D(n_9441), .SD(n_62313), .Q(\tab12[14] 
		));
	notech_mux2 i_10724(.S(\nbus_14508[0] ), .A(\tab12[14] ), .B(n_56711), .Z
		(n_9441));
	notech_and4 i_858(.A(n_1125), .B(n_1123), .C(n_864), .D(n_867), .Z(n_1127
		));
	notech_reg_set tab12_reg_15(.CP(n_63047), .D(n_9447), .SD(n_62313), .Q(\tab12[15] 
		));
	notech_mux2 i_10732(.S(\nbus_14508[0] ), .A(\tab12[15] ), .B(n_56717), .Z
		(n_9447));
	notech_ao4 i_851(.A(n_1100), .B(n_11890), .C(n_1098), .D(n_12057), .Z(n_1128
		));
	notech_reg_set tab12_reg_16(.CP(n_63047), .D(n_9453), .SD(n_62313), .Q(\tab12[16] 
		));
	notech_mux2 i_10740(.S(\nbus_14508[0] ), .A(\tab12[16] ), .B(n_56723), .Z
		(n_9453));
	notech_reg_set tab12_reg_17(.CP(n_63075), .D(n_9459), .SD(n_62341), .Q(\tab12[17] 
		));
	notech_mux2 i_10748(.S(n_56101), .A(\tab12[17] ), .B(n_56729), .Z(n_9459
		));
	notech_ao4 i_850(.A(n_62893), .B(n_12134), .C(n_1043), .D(n_12058), .Z(n_1130
		));
	notech_reg_set tab12_reg_18(.CP(n_63075), .D(n_9465), .SD(n_62341), .Q(\tab12[18] 
		));
	notech_mux2 i_10756(.S(n_56101), .A(\tab12[18] ), .B(n_56735), .Z(n_9465
		));
	notech_reg_set tab12_reg_19(.CP(n_63075), .D(n_9471), .SD(n_62341), .Q(\tab12[19] 
		));
	notech_mux2 i_10764(.S(n_56101), .A(\tab12[19] ), .B(n_56741), .Z(n_9471
		));
	notech_ao4 i_847(.A(n_1086), .B(n_11912), .C(n_1084), .D(n_11941), .Z(n_1132
		));
	notech_reg_set tab12_reg_20(.CP(n_63075), .D(n_9477), .SD(n_62341), .Q(\tab12[20] 
		));
	notech_mux2 i_10772(.S(n_56101), .A(\tab12[20] ), .B(n_56747), .Z(n_9477
		));
	notech_reg_set tab12_reg_21(.CP(n_63075), .D(n_9483), .SD(n_62341), .Q(\tab12[21] 
		));
	notech_mux2 i_10780(.S(n_56101), .A(\tab12[21] ), .B(n_56753), .Z(n_9483
		));
	notech_ao4 i_845(.A(n_1092), .B(n_11962), .C(n_1090), .D(n_11982), .Z(n_1134
		));
	notech_reg_set tab12_reg_22(.CP(n_63075), .D(n_9489), .SD(n_62341), .Q(\tab12[22] 
		));
	notech_mux2 i_10788(.S(n_56101), .A(\tab12[22] ), .B(n_56759), .Z(n_9489
		));
	notech_reg_set tab12_reg_23(.CP(n_63075), .D(n_9495), .SD(n_62341), .Q(\tab12[23] 
		));
	notech_mux2 i_10796(.S(n_56101), .A(\tab12[23] ), .B(n_56765), .Z(n_9495
		));
	notech_and4 i_849(.A(n_1134), .B(n_1132), .C(n_853), .D(n_856), .Z(n_1136
		));
	notech_reg_set tab12_reg_24(.CP(n_63075), .D(n_9501), .SD(n_62341), .Q(\tab12[24] 
		));
	notech_mux2 i_10804(.S(n_56101), .A(\tab12[24] ), .B(n_56771), .Z(n_9501
		));
	notech_ao4 i_842(.A(n_1100), .B(n_11889), .C(n_1098), .D(n_12055), .Z(n_1137
		));
	notech_reg_set tab12_reg_25(.CP(n_63075), .D(n_9507), .SD(n_62341), .Q(\tab12[25] 
		));
	notech_mux2 i_10812(.S(n_56101), .A(\tab12[25] ), .B(n_56777), .Z(n_9507
		));
	notech_reg_set tab12_reg_26(.CP(n_63076), .D(n_9513), .SD(n_62342), .Q(\tab12[26] 
		));
	notech_mux2 i_10820(.S(n_56101), .A(\tab12[26] ), .B(n_56783), .Z(n_9513
		));
	notech_ao4 i_841(.A(n_62893), .B(n_12133), .C(n_1043), .D(n_12056), .Z(n_1139
		));
	notech_reg_set tab12_reg_27(.CP(n_63076), .D(n_9519), .SD(n_62342), .Q(\tab12[27] 
		));
	notech_mux2 i_10828(.S(\nbus_14508[0] ), .A(\tab12[27] ), .B(n_56789), .Z
		(n_9519));
	notech_reg_set tab12_reg_28(.CP(n_63076), .D(n_9525), .SD(n_62342), .Q(\tab12[28] 
		));
	notech_mux2 i_10836(.S(n_56101), .A(\tab12[28] ), .B(n_56795), .Z(n_9525
		));
	notech_ao4 i_838(.A(n_1086), .B(n_11911), .C(n_1084), .D(n_11940), .Z(n_1141
		));
	notech_reg_set tab12_reg_29(.CP(n_63076), .D(n_9531), .SD(n_62342), .Q(\tab12[29] 
		));
	notech_mux2 i_10844(.S(n_56101), .A(\tab12[29] ), .B(n_56801), .Z(n_9531
		));
	notech_reg tab12_reg_30(.CP(n_63076), .D(n_9537), .CD(n_62342), .Q(\tab12[30] 
		));
	notech_mux2 i_10852(.S(n_56101), .A(\tab12[30] ), .B(n_974), .Z(n_9537)
		);
	notech_ao4 i_836(.A(n_1092), .B(n_11961), .C(n_1090), .D(n_11981), .Z(n_1143
		));
	notech_reg tab12_reg_32(.CP(n_63075), .D(n_9543), .CD(n_62341), .Q(\tab12[32] 
		));
	notech_mux2 i_10860(.S(n_56101), .A(\tab12[32] ), .B(n_975), .Z(n_9543)
		);
	notech_reg_set tab12_reg_33(.CP(n_63075), .D(n_9549), .SD(n_62341), .Q(\tab12[33] 
		));
	notech_mux2 i_10868(.S(n_56101), .A(\tab12[33] ), .B(n_56153), .Z(n_9549
		));
	notech_and4 i_840(.A(n_1143), .B(n_1141), .C(n_842), .D(n_845), .Z(n_1145
		));
	notech_reg hit_adr12_reg(.CP(n_63076), .D(n_9555), .CD(n_62342), .Q(hit_adr12
		));
	notech_mux2 i_10876(.S(n_971), .A(hit_add12), .B(hit_adr12), .Z(n_9555)
		);
	notech_ao4 i_833(.A(n_1100), .B(n_11888), .C(n_1098), .D(n_12053), .Z(n_1146
		));
	notech_reg_set tab13_reg_0(.CP(n_63076), .D(n_9561), .SD(n_62342), .Q(\tab13[0] 
		));
	notech_mux2 i_10884(.S(\nbus_14492[0] ), .A(\tab13[0] ), .B(n_56627), .Z
		(n_9561));
	notech_reg_set tab13_reg_1(.CP(n_63071), .D(n_9567), .SD(n_62337), .Q(\tab13[1] 
		));
	notech_mux2 i_10892(.S(\nbus_14492[0] ), .A(\tab13[1] ), .B(n_56633), .Z
		(n_9567));
	notech_ao4 i_832(.A(n_62893), .B(n_12132), .C(n_1043), .D(n_12054), .Z(n_1148
		));
	notech_reg_set tab13_reg_2(.CP(n_63071), .D(n_9573), .SD(n_62337), .Q(\tab13[2] 
		));
	notech_mux2 i_10900(.S(\nbus_14492[0] ), .A(\tab13[2] ), .B(n_56639), .Z
		(n_9573));
	notech_reg_set tab13_reg_3(.CP(n_63074), .D(n_9579), .SD(n_62340), .Q(\tab13[3] 
		));
	notech_mux2 i_10908(.S(\nbus_14492[0] ), .A(\tab13[3] ), .B(n_56645), .Z
		(n_9579));
	notech_ao4 i_829(.A(n_1086), .B(n_11910), .C(n_1084), .D(n_11939), .Z(n_1150
		));
	notech_reg tab13_reg_4(.CP(n_63074), .D(n_9585), .CD(n_62340), .Q(\tab13[4] 
		));
	notech_mux2 i_10916(.S(\nbus_14492[0] ), .A(\tab13[4] ), .B(n_973), .Z(n_9585
		));
	notech_reg_set tab13_reg_5(.CP(n_63071), .D(n_9591), .SD(n_62337), .Q(\tab13[5] 
		));
	notech_mux2 i_10924(.S(\nbus_14492[0] ), .A(\tab13[5] ), .B(n_56657), .Z
		(n_9591));
	notech_ao4 i_827(.A(n_1092), .B(n_11960), .C(n_1090), .D(n_11980), .Z(n_1152
		));
	notech_reg_set tab13_reg_6(.CP(n_63071), .D(n_9597), .SD(n_62337), .Q(\tab13[6] 
		));
	notech_mux2 i_10932(.S(\nbus_14492[0] ), .A(\tab13[6] ), .B(n_56663), .Z
		(n_9597));
	notech_reg_set tab13_reg_7(.CP(n_63071), .D(n_9603), .SD(n_62337), .Q(\tab13[7] 
		));
	notech_mux2 i_10940(.S(\nbus_14492[0] ), .A(\tab13[7] ), .B(n_56669), .Z
		(n_9603));
	notech_and4 i_831(.A(n_1152), .B(n_1150), .C(n_831), .D(n_834), .Z(n_1154
		));
	notech_reg_set tab13_reg_8(.CP(n_63071), .D(n_9609), .SD(n_62337), .Q(\tab13[8] 
		));
	notech_mux2 i_10948(.S(\nbus_14492[0] ), .A(\tab13[8] ), .B(n_56675), .Z
		(n_9609));
	notech_ao4 i_824(.A(n_1100), .B(n_11887), .C(n_1098), .D(n_12051), .Z(n_1155
		));
	notech_reg_set tab13_reg_9(.CP(n_63071), .D(n_9615), .SD(n_62337), .Q(\tab13[9] 
		));
	notech_mux2 i_10956(.S(\nbus_14492[0] ), .A(\tab13[9] ), .B(n_56681), .Z
		(n_9615));
	notech_reg_set tab13_reg_10(.CP(n_63074), .D(n_9621), .SD(n_62340), .Q(\tab13[10] 
		));
	notech_mux2 i_10964(.S(\nbus_14492[0] ), .A(\tab13[10] ), .B(n_56687), .Z
		(n_9621));
	notech_ao4 i_823(.A(n_62893), .B(n_12131), .C(n_1043), .D(n_12052), .Z(n_1157
		));
	notech_reg_set tab13_reg_11(.CP(n_63074), .D(n_9627), .SD(n_62340), .Q(\tab13[11] 
		));
	notech_mux2 i_10972(.S(\nbus_14492[0] ), .A(\tab13[11] ), .B(n_56693), .Z
		(n_9627));
	notech_reg_set tab13_reg_12(.CP(n_63074), .D(n_9633), .SD(n_62340), .Q(\tab13[12] 
		));
	notech_mux2 i_10980(.S(\nbus_14492[0] ), .A(\tab13[12] ), .B(n_56699), .Z
		(n_9633));
	notech_ao4 i_820(.A(n_1086), .B(n_11909), .C(n_1084), .D(n_11938), .Z(n_1159
		));
	notech_reg_set tab13_reg_13(.CP(n_63074), .D(n_9639), .SD(n_62340), .Q(\tab13[13] 
		));
	notech_mux2 i_10988(.S(\nbus_14492[0] ), .A(\tab13[13] ), .B(n_56705), .Z
		(n_9639));
	notech_reg_set tab13_reg_14(.CP(n_63074), .D(n_9645), .SD(n_62340), .Q(\tab13[14] 
		));
	notech_mux2 i_10996(.S(\nbus_14492[0] ), .A(\tab13[14] ), .B(n_56711), .Z
		(n_9645));
	notech_ao4 i_818(.A(n_1092), .B(n_11959), .C(n_1090), .D(n_11979), .Z(n_1161
		));
	notech_reg_set tab13_reg_15(.CP(n_63074), .D(n_9651), .SD(n_62340), .Q(\tab13[15] 
		));
	notech_mux2 i_11004(.S(\nbus_14492[0] ), .A(\tab13[15] ), .B(n_56717), .Z
		(n_9651));
	notech_reg_set tab13_reg_16(.CP(n_63074), .D(n_9657), .SD(n_62340), .Q(\tab13[16] 
		));
	notech_mux2 i_11012(.S(\nbus_14492[0] ), .A(\tab13[16] ), .B(n_56723), .Z
		(n_9657));
	notech_and4 i_822(.A(n_1161), .B(n_1159), .C(n_820), .D(n_823), .Z(n_1163
		));
	notech_reg_set tab13_reg_17(.CP(n_63074), .D(n_9663), .SD(n_62340), .Q(\tab13[17] 
		));
	notech_mux2 i_11020(.S(n_56083), .A(\tab13[17] ), .B(n_56729), .Z(n_9663
		));
	notech_ao4 i_815(.A(n_1100), .B(n_11886), .C(n_1098), .D(n_12049), .Z(n_1164
		));
	notech_reg_set tab13_reg_18(.CP(n_63074), .D(n_9669), .SD(n_62340), .Q(\tab13[18] 
		));
	notech_mux2 i_11028(.S(n_56083), .A(\tab13[18] ), .B(n_56735), .Z(n_9669
		));
	notech_reg_set tab13_reg_19(.CP(n_63076), .D(n_9675), .SD(n_62342), .Q(\tab13[19] 
		));
	notech_mux2 i_11036(.S(n_56083), .A(\tab13[19] ), .B(n_56741), .Z(n_9675
		));
	notech_ao4 i_814(.A(n_62893), .B(n_12130), .C(n_1043), .D(n_12050), .Z(n_1166
		));
	notech_reg_set tab13_reg_20(.CP(n_63079), .D(n_9681), .SD(n_62345), .Q(\tab13[20] 
		));
	notech_mux2 i_11044(.S(n_56083), .A(\tab13[20] ), .B(n_56747), .Z(n_9681
		));
	notech_reg_set tab13_reg_21(.CP(n_63079), .D(n_9687), .SD(n_62345), .Q(\tab13[21] 
		));
	notech_mux2 i_11052(.S(n_56083), .A(\tab13[21] ), .B(n_56753), .Z(n_9687
		));
	notech_ao4 i_811(.A(n_1086), .B(n_11908), .C(n_1084), .D(n_11937), .Z(n_1168
		));
	notech_reg_set tab13_reg_22(.CP(n_63080), .D(n_9693), .SD(n_62346), .Q(\tab13[22] 
		));
	notech_mux2 i_11060(.S(n_56083), .A(\tab13[22] ), .B(n_56759), .Z(n_9693
		));
	notech_reg_set tab13_reg_23(.CP(n_63080), .D(n_9699), .SD(n_62346), .Q(\tab13[23] 
		));
	notech_mux2 i_11068(.S(n_56083), .A(\tab13[23] ), .B(n_56765), .Z(n_9699
		));
	notech_ao4 i_809(.A(n_1092), .B(n_11958), .C(n_1090), .D(n_11978), .Z(n_1170
		));
	notech_reg_set tab13_reg_24(.CP(n_63079), .D(n_9705), .SD(n_62345), .Q(\tab13[24] 
		));
	notech_mux2 i_11076(.S(n_56083), .A(\tab13[24] ), .B(n_56771), .Z(n_9705
		));
	notech_reg_set tab13_reg_25(.CP(n_63079), .D(n_9711), .SD(n_62345), .Q(\tab13[25] 
		));
	notech_mux2 i_11084(.S(n_56083), .A(\tab13[25] ), .B(n_56777), .Z(n_9711
		));
	notech_and4 i_813(.A(n_1170), .B(n_1168), .C(n_809), .D(n_812), .Z(n_1172
		));
	notech_reg_set tab13_reg_26(.CP(n_63079), .D(n_9717), .SD(n_62345), .Q(\tab13[26] 
		));
	notech_mux2 i_11092(.S(n_56083), .A(\tab13[26] ), .B(n_56783), .Z(n_9717
		));
	notech_ao4 i_806(.A(n_1100), .B(n_11885), .C(n_1098), .D(n_12047), .Z(n_1173
		));
	notech_reg_set tab13_reg_27(.CP(n_63079), .D(n_9723), .SD(n_62345), .Q(\tab13[27] 
		));
	notech_mux2 i_11100(.S(\nbus_14492[0] ), .A(\tab13[27] ), .B(n_56789), .Z
		(n_9723));
	notech_reg_set tab13_reg_28(.CP(n_63079), .D(n_9729), .SD(n_62345), .Q(\tab13[28] 
		));
	notech_mux2 i_11108(.S(n_56083), .A(\tab13[28] ), .B(n_56795), .Z(n_9729
		));
	notech_ao4 i_805(.A(n_62893), .B(n_12129), .C(n_1043), .D(n_12048), .Z(n_1175
		));
	notech_reg_set tab13_reg_29(.CP(n_63080), .D(n_9735), .SD(n_62346), .Q(\tab13[29] 
		));
	notech_mux2 i_11116(.S(n_56083), .A(\tab13[29] ), .B(n_56801), .Z(n_9735
		));
	notech_reg tab13_reg_30(.CP(n_63080), .D(n_9741), .CD(n_62346), .Q(\tab13[30] 
		));
	notech_mux2 i_11124(.S(n_56083), .A(\tab13[30] ), .B(n_974), .Z(n_9741)
		);
	notech_ao4 i_802(.A(n_1086), .B(n_11907), .C(n_1084), .D(n_11936), .Z(n_1177
		));
	notech_reg tab13_reg_32(.CP(n_63080), .D(n_9747), .CD(n_62346), .Q(\tab13[32] 
		));
	notech_mux2 i_11132(.S(n_56083), .A(\tab13[32] ), .B(n_975), .Z(n_9747)
		);
	notech_reg_set tab13_reg_33(.CP(n_63080), .D(n_9753), .SD(n_62346), .Q(\tab13[33] 
		));
	notech_mux2 i_11140(.S(n_56083), .A(\tab13[33] ), .B(n_56153), .Z(n_9753
		));
	notech_ao4 i_800(.A(n_1092), .B(n_11957), .C(n_1090), .D(n_11977), .Z(n_1179
		));
	notech_reg hit_adr13_reg(.CP(n_63080), .D(n_9759), .CD(n_62346), .Q(hit_adr13
		));
	notech_mux2 i_11148(.S(n_971), .A(hit_add13), .B(hit_adr13), .Z(n_9759)
		);
	notech_reg_set tab14_reg_0(.CP(n_63080), .D(n_9765), .SD(n_62346), .Q(\tab14[0] 
		));
	notech_mux2 i_11156(.S(\nbus_14489[0] ), .A(\tab14[0] ), .B(n_56627), .Z
		(n_9765));
	notech_and4 i_804(.A(n_1179), .B(n_1177), .C(n_798), .D(n_801), .Z(n_1181
		));
	notech_reg_set tab14_reg_1(.CP(n_63080), .D(n_9771), .SD(n_62346), .Q(\tab14[1] 
		));
	notech_mux2 i_11164(.S(\nbus_14489[0] ), .A(\tab14[1] ), .B(n_56633), .Z
		(n_9771));
	notech_ao4 i_797(.A(n_1100), .B(n_11884), .C(n_1098), .D(n_12045), .Z(n_1182
		));
	notech_reg_set tab14_reg_2(.CP(n_63080), .D(n_9777), .SD(n_62346), .Q(\tab14[2] 
		));
	notech_mux2 i_11172(.S(\nbus_14489[0] ), .A(\tab14[2] ), .B(n_56639), .Z
		(n_9777));
	notech_reg_set tab14_reg_3(.CP(n_63080), .D(n_9783), .SD(n_62346), .Q(\tab14[3] 
		));
	notech_mux2 i_11180(.S(\nbus_14489[0] ), .A(\tab14[3] ), .B(n_56645), .Z
		(n_9783));
	notech_ao4 i_796(.A(n_62893), .B(n_12128), .C(n_56301), .D(n_12046), .Z(n_1184
		));
	notech_reg tab14_reg_4(.CP(n_63078), .D(n_9789), .CD(n_62344), .Q(\tab14[4] 
		));
	notech_mux2 i_11188(.S(\nbus_14489[0] ), .A(\tab14[4] ), .B(n_973), .Z(n_9789
		));
	notech_reg_set tab14_reg_5(.CP(n_63078), .D(n_9795), .SD(n_62344), .Q(\tab14[5] 
		));
	notech_mux2 i_11196(.S(\nbus_14489[0] ), .A(\tab14[5] ), .B(n_56657), .Z
		(n_9795));
	notech_ao4 i_793(.A(n_1086), .B(n_11906), .C(n_1084), .D(n_11935), .Z(n_1186
		));
	notech_reg_set tab14_reg_6(.CP(n_63078), .D(n_9801), .SD(n_62344), .Q(\tab14[6] 
		));
	notech_mux2 i_11204(.S(\nbus_14489[0] ), .A(\tab14[6] ), .B(n_56663), .Z
		(n_9801));
	notech_reg_set tab14_reg_7(.CP(n_63078), .D(n_9807), .SD(n_62344), .Q(\tab14[7] 
		));
	notech_mux2 i_11212(.S(\nbus_14489[0] ), .A(\tab14[7] ), .B(n_56669), .Z
		(n_9807));
	notech_ao4 i_791(.A(n_1092), .B(n_11956), .C(n_1090), .D(n_11976), .Z(n_1188
		));
	notech_reg_set tab14_reg_8(.CP(n_63078), .D(n_9813), .SD(n_62344), .Q(\tab14[8] 
		));
	notech_mux2 i_11220(.S(\nbus_14489[0] ), .A(\tab14[8] ), .B(n_56675), .Z
		(n_9813));
	notech_reg_set tab14_reg_9(.CP(n_63076), .D(n_9819), .SD(n_62342), .Q(\tab14[9] 
		));
	notech_mux2 i_11228(.S(\nbus_14489[0] ), .A(\tab14[9] ), .B(n_56681), .Z
		(n_9819));
	notech_and4 i_795(.A(n_1188), .B(n_1186), .C(n_787), .D(n_790), .Z(n_1190
		));
	notech_reg_set tab14_reg_10(.CP(n_63076), .D(n_9825), .SD(n_62342), .Q(\tab14[10] 
		));
	notech_mux2 i_11236(.S(\nbus_14489[0] ), .A(\tab14[10] ), .B(n_56687), .Z
		(n_9825));
	notech_ao4 i_788(.A(n_1100), .B(n_11883), .C(n_1098), .D(n_12043), .Z(n_1191
		));
	notech_reg_set tab14_reg_11(.CP(n_63078), .D(n_9831), .SD(n_62344), .Q(\tab14[11] 
		));
	notech_mux2 i_11244(.S(\nbus_14489[0] ), .A(\tab14[11] ), .B(n_56693), .Z
		(n_9831));
	notech_reg_set tab14_reg_12(.CP(n_63076), .D(n_9837), .SD(n_62342), .Q(\tab14[12] 
		));
	notech_mux2 i_11252(.S(\nbus_14489[0] ), .A(\tab14[12] ), .B(n_56699), .Z
		(n_9837));
	notech_ao4 i_787(.A(n_62898), .B(n_12127), .C(n_56301), .D(n_12044), .Z(n_1193
		));
	notech_reg_set tab14_reg_13(.CP(n_63079), .D(n_9843), .SD(n_62345), .Q(\tab14[13] 
		));
	notech_mux2 i_11260(.S(\nbus_14489[0] ), .A(\tab14[13] ), .B(n_56705), .Z
		(n_9843));
	notech_reg_set tab14_reg_14(.CP(n_63079), .D(n_9849), .SD(n_62345), .Q(\tab14[14] 
		));
	notech_mux2 i_11268(.S(\nbus_14489[0] ), .A(\tab14[14] ), .B(n_56711), .Z
		(n_9849));
	notech_ao4 i_784(.A(n_1086), .B(n_11905), .C(n_1084), .D(n_11934), .Z(n_1195
		));
	notech_reg_set tab14_reg_15(.CP(n_63079), .D(n_9855), .SD(n_62345), .Q(\tab14[15] 
		));
	notech_mux2 i_11276(.S(\nbus_14489[0] ), .A(\tab14[15] ), .B(n_56717), .Z
		(n_9855));
	notech_reg_set tab14_reg_16(.CP(n_63079), .D(n_9861), .SD(n_62345), .Q(\tab14[16] 
		));
	notech_mux2 i_11284(.S(\nbus_14489[0] ), .A(\tab14[16] ), .B(n_56723), .Z
		(n_9861));
	notech_ao4 i_782(.A(n_1092), .B(n_11955), .C(n_1090), .D(n_11975), .Z(n_1197
		));
	notech_reg_set tab14_reg_17(.CP(n_63078), .D(n_9867), .SD(n_62344), .Q(\tab14[17] 
		));
	notech_mux2 i_11292(.S(n_56074), .A(\tab14[17] ), .B(n_56729), .Z(n_9867
		));
	notech_reg_set tab14_reg_18(.CP(n_63078), .D(n_9873), .SD(n_62344), .Q(\tab14[18] 
		));
	notech_mux2 i_11300(.S(n_56074), .A(\tab14[18] ), .B(n_56735), .Z(n_9873
		));
	notech_and4 i_786(.A(n_1197), .B(n_1195), .C(n_776), .D(n_779), .Z(n_1199
		));
	notech_reg_set tab14_reg_19(.CP(n_63078), .D(n_9879), .SD(n_62344), .Q(\tab14[19] 
		));
	notech_mux2 i_11308(.S(n_56074), .A(\tab14[19] ), .B(n_56741), .Z(n_9879
		));
	notech_ao4 i_779(.A(n_1100), .B(n_11882), .C(n_1098), .D(n_12041), .Z(n_1200
		));
	notech_reg_set tab14_reg_20(.CP(n_63078), .D(n_9885), .SD(n_62344), .Q(\tab14[20] 
		));
	notech_mux2 i_11316(.S(n_56074), .A(\tab14[20] ), .B(n_56747), .Z(n_9885
		));
	notech_reg_set tab14_reg_21(.CP(n_63078), .D(n_9891), .SD(n_62344), .Q(\tab14[21] 
		));
	notech_mux2 i_11324(.S(n_56074), .A(\tab14[21] ), .B(n_56753), .Z(n_9891
		));
	notech_ao4 i_778(.A(n_62898), .B(n_12126), .C(n_56301), .D(n_12042), .Z(n_1202
		));
	notech_reg_set tab14_reg_22(.CP(n_63071), .D(n_9897), .SD(n_62337), .Q(\tab14[22] 
		));
	notech_mux2 i_11332(.S(n_56074), .A(\tab14[22] ), .B(n_56759), .Z(n_9897
		));
	notech_reg_set tab14_reg_23(.CP(n_63065), .D(n_9903), .SD(n_62331), .Q(\tab14[23] 
		));
	notech_mux2 i_11340(.S(n_56074), .A(\tab14[23] ), .B(n_56765), .Z(n_9903
		));
	notech_ao4 i_775(.A(n_1086), .B(n_11904), .C(n_1084), .D(n_11933), .Z(n_1204
		));
	notech_reg_set tab14_reg_24(.CP(n_63065), .D(n_9909), .SD(n_62331), .Q(\tab14[24] 
		));
	notech_mux2 i_11348(.S(n_56074), .A(\tab14[24] ), .B(n_56771), .Z(n_9909
		));
	notech_reg_set tab14_reg_25(.CP(n_63066), .D(n_9915), .SD(n_62332), .Q(\tab14[25] 
		));
	notech_mux2 i_11356(.S(n_56074), .A(\tab14[25] ), .B(n_56777), .Z(n_9915
		));
	notech_ao4 i_773(.A(n_1092), .B(n_11954), .C(n_1090), .D(n_11974), .Z(n_1206
		));
	notech_reg_set tab14_reg_26(.CP(n_63065), .D(n_9921), .SD(n_62331), .Q(\tab14[26] 
		));
	notech_mux2 i_11364(.S(n_56074), .A(\tab14[26] ), .B(n_56783), .Z(n_9921
		));
	notech_reg_set tab14_reg_27(.CP(n_63065), .D(n_9927), .SD(n_62331), .Q(\tab14[27] 
		));
	notech_mux2 i_11372(.S(\nbus_14489[0] ), .A(\tab14[27] ), .B(n_56789), .Z
		(n_9927));
	notech_and4 i_777(.A(n_1206), .B(n_1204), .C(n_765), .D(n_768), .Z(n_1208
		));
	notech_reg_set tab14_reg_28(.CP(n_63065), .D(n_9933), .SD(n_62331), .Q(\tab14[28] 
		));
	notech_mux2 i_11380(.S(n_56074), .A(\tab14[28] ), .B(n_56795), .Z(n_9933
		));
	notech_ao4 i_770(.A(n_1100), .B(n_11880), .C(n_1098), .D(n_12039), .Z(n_1209
		));
	notech_reg_set tab14_reg_29(.CP(n_63065), .D(n_9939), .SD(n_62331), .Q(\tab14[29] 
		));
	notech_mux2 i_11388(.S(n_56074), .A(\tab14[29] ), .B(n_56801), .Z(n_9939
		));
	notech_reg tab14_reg_30(.CP(n_63065), .D(n_9945), .CD(n_62331), .Q(\tab14[30] 
		));
	notech_mux2 i_11396(.S(n_56074), .A(\tab14[30] ), .B(n_974), .Z(n_9945)
		);
	notech_ao4 i_769(.A(n_62898), .B(n_12125), .C(n_56301), .D(n_12040), .Z(n_1211
		));
	notech_reg tab14_reg_32(.CP(n_63065), .D(n_9951), .CD(n_62331), .Q(\tab14[32] 
		));
	notech_mux2 i_11404(.S(n_56074), .A(\tab14[32] ), .B(n_975), .Z(n_9951)
		);
	notech_reg_set tab14_reg_33(.CP(n_63066), .D(n_9957), .SD(n_62332), .Q(\tab14[33] 
		));
	notech_mux2 i_11412(.S(n_56074), .A(\tab14[33] ), .B(n_56153), .Z(n_9957
		));
	notech_ao4 i_766(.A(n_1086), .B(n_11903), .C(n_1084), .D(n_11932), .Z(n_1213
		));
	notech_reg hit_adr14_reg(.CP(n_63066), .D(n_9963), .CD(n_62332), .Q(hit_adr14
		));
	notech_mux2 i_11420(.S(n_971), .A(hit_add14), .B(hit_adr14), .Z(n_9963)
		);
	notech_reg nx_tab1_reg_0(.CP(n_63066), .D(n_9969), .CD(n_62332), .Q(\nx_tab1[0] 
		));
	notech_mux2 i_11428(.S(\nbus_14512[0] ), .A(\nx_tab1[0] ), .B(n_11917), 
		.Z(n_9969));
	notech_ao4 i_764(.A(n_1092), .B(n_11953), .C(n_1090), .D(n_11973), .Z(n_1215
		));
	notech_reg nx_tab1_reg_1(.CP(n_63066), .D(n_9975), .CD(n_62332), .Q(\nx_tab1[1] 
		));
	notech_mux2 i_11436(.S(\nbus_14512[0] ), .A(\nx_tab1[1] ), .B(n_11919), 
		.Z(n_9975));
	notech_reg_set nnx_tab1_reg_0(.CP(n_63066), .D(n_9981), .SD(n_62332), .Q
		(\nnx_tab1[0] ));
	notech_mux2 i_11444(.S(n_11925), .A(\nnx_tab1[0] ), .B(n_11921), .Z(n_9981
		));
	notech_and4 i_768(.A(n_1215), .B(n_1213), .C(n_754), .D(n_757), .Z(n_1217
		));
	notech_reg nnx_tab1_reg_1(.CP(n_63066), .D(n_9987), .CD(n_62332), .Q(\nnx_tab1[1] 
		));
	notech_mux2 i_11452(.S(n_11925), .A(\nnx_tab1[1] ), .B(n_11923), .Z(n_9987
		));
	notech_ao4 i_761(.A(n_1100), .B(n_11879), .C(n_1098), .D(n_12037), .Z(n_1218
		));
	notech_reg hit_adr21_reg(.CP(n_63066), .D(n_9993), .CD(n_62332), .Q(hit_adr21
		));
	notech_mux2 i_11460(.S(n_971), .A(hit_add21), .B(hit_adr21), .Z(n_9993)
		);
	notech_reg_set tab22_reg_0(.CP(n_63066), .D(n_9999), .SD(n_62332), .Q(\tab22[0] 
		));
	notech_mux2 i_11468(.S(\nbus_14520[0] ), .A(\tab22[0] ), .B(n_56627), .Z
		(n_9999));
	notech_ao4 i_760(.A(n_62898), .B(n_12124), .C(n_56301), .D(n_12038), .Z(n_1220
		));
	notech_reg_set tab22_reg_1(.CP(n_63066), .D(n_10005), .SD(n_62332), .Q(\tab22[1] 
		));
	notech_mux2 i_11476(.S(\nbus_14520[0] ), .A(\tab22[1] ), .B(n_56633), .Z
		(n_10005));
	notech_reg_set tab22_reg_2(.CP(n_63062), .D(n_10011), .SD(n_62328), .Q(\tab22[2] 
		));
	notech_mux2 i_11484(.S(\nbus_14520[0] ), .A(\tab22[2] ), .B(n_56639), .Z
		(n_10011));
	notech_ao4 i_756(.A(n_1086), .B(n_11902), .C(n_1084), .D(n_11931), .Z(n_1222
		));
	notech_reg_set tab22_reg_3(.CP(n_63062), .D(n_10017), .SD(n_62328), .Q(\tab22[3] 
		));
	notech_mux2 i_11492(.S(\nbus_14520[0] ), .A(\tab22[3] ), .B(n_56645), .Z
		(n_10017));
	notech_reg tab22_reg_4(.CP(n_63062), .D(n_10023), .CD(n_62328), .Q(\tab22[4] 
		));
	notech_mux2 i_11500(.S(\nbus_14520[0] ), .A(\tab22[4] ), .B(n_973), .Z(n_10023
		));
	notech_ao4 i_754(.A(n_1092), .B(n_11952), .C(n_1090), .D(n_11972), .Z(n_1224
		));
	notech_reg_set tab22_reg_5(.CP(n_63062), .D(n_10029), .SD(n_62328), .Q(\tab22[5] 
		));
	notech_mux2 i_11508(.S(\nbus_14520[0] ), .A(\tab22[5] ), .B(n_56657), .Z
		(n_10029));
	notech_reg_set tab22_reg_6(.CP(n_63062), .D(n_10035), .SD(n_62328), .Q(\tab22[6] 
		));
	notech_mux2 i_11516(.S(\nbus_14520[0] ), .A(\tab22[6] ), .B(n_56663), .Z
		(n_10035));
	notech_and4 i_758(.A(n_1224), .B(n_1222), .C(n_743), .D(n_746), .Z(n_1226
		));
	notech_reg_set tab22_reg_7(.CP(n_63061), .D(n_10041), .SD(n_62327), .Q(\tab22[7] 
		));
	notech_mux2 i_11524(.S(\nbus_14520[0] ), .A(\tab22[7] ), .B(n_56669), .Z
		(n_10041));
	notech_ao4 i_751(.A(n_1100), .B(n_11878), .C(n_1098), .D(n_12035), .Z(n_1227
		));
	notech_reg_set tab22_reg_8(.CP(n_63061), .D(n_10047), .SD(n_62327), .Q(\tab22[8] 
		));
	notech_mux2 i_11532(.S(\nbus_14520[0] ), .A(\tab22[8] ), .B(n_56675), .Z
		(n_10047));
	notech_reg_set tab22_reg_9(.CP(n_63061), .D(n_10053), .SD(n_62327), .Q(\tab22[9] 
		));
	notech_mux2 i_11540(.S(\nbus_14520[0] ), .A(\tab22[9] ), .B(n_56681), .Z
		(n_10053));
	notech_ao4 i_750(.A(n_62898), .B(n_12123), .C(n_56301), .D(n_12036), .Z(n_1229
		));
	notech_reg_set tab22_reg_10(.CP(n_63061), .D(n_10059), .SD(n_62327), .Q(\tab22[10] 
		));
	notech_mux2 i_11548(.S(\nbus_14520[0] ), .A(\tab22[10] ), .B(n_56687), .Z
		(n_10059));
	notech_reg_set tab22_reg_11(.CP(n_63065), .D(n_10065), .SD(n_62331), .Q(\tab22[11] 
		));
	notech_mux2 i_11556(.S(\nbus_14520[0] ), .A(\tab22[11] ), .B(n_56693), .Z
		(n_10065));
	notech_ao4 i_747(.A(n_1086), .B(n_11901), .C(n_1084), .D(n_11930), .Z(n_1231
		));
	notech_reg_set tab22_reg_12(.CP(n_63062), .D(n_10071), .SD(n_62328), .Q(\tab22[12] 
		));
	notech_mux2 i_11564(.S(\nbus_14520[0] ), .A(\tab22[12] ), .B(n_56699), .Z
		(n_10071));
	notech_reg_set tab22_reg_13(.CP(n_63065), .D(n_10077), .SD(n_62331), .Q(\tab22[13] 
		));
	notech_mux2 i_11572(.S(\nbus_14520[0] ), .A(\tab22[13] ), .B(n_56705), .Z
		(n_10077));
	notech_ao4 i_745(.A(n_1092), .B(n_11951), .C(n_1090), .D(n_11971), .Z(n_1233
		));
	notech_reg_set tab22_reg_14(.CP(n_63065), .D(n_10083), .SD(n_62331), .Q(\tab22[14] 
		));
	notech_mux2 i_11580(.S(\nbus_14520[0] ), .A(\tab22[14] ), .B(n_56711), .Z
		(n_10083));
	notech_reg_set tab22_reg_15(.CP(n_63062), .D(n_10089), .SD(n_62328), .Q(\tab22[15] 
		));
	notech_mux2 i_11588(.S(\nbus_14520[0] ), .A(\tab22[15] ), .B(n_56717), .Z
		(n_10089));
	notech_and4 i_749(.A(n_1233), .B(n_1231), .C(n_732), .D(n_735), .Z(n_1235
		));
	notech_reg_set tab22_reg_16(.CP(n_63062), .D(n_10095), .SD(n_62328), .Q(\tab22[16] 
		));
	notech_mux2 i_11596(.S(\nbus_14520[0] ), .A(\tab22[16] ), .B(n_56723), .Z
		(n_10095));
	notech_ao4 i_742(.A(n_1100), .B(n_11877), .C(n_1098), .D(n_12033), .Z(n_1236
		));
	notech_reg_set tab22_reg_17(.CP(n_63062), .D(n_10101), .SD(n_62328), .Q(\tab22[17] 
		));
	notech_mux2 i_11604(.S(n_56159), .A(\tab22[17] ), .B(n_56729), .Z(n_10101
		));
	notech_reg_set tab22_reg_18(.CP(n_63062), .D(n_10107), .SD(n_62328), .Q(\tab22[18] 
		));
	notech_mux2 i_11612(.S(n_56159), .A(\tab22[18] ), .B(n_56735), .Z(n_10107
		));
	notech_ao4 i_741(.A(n_62898), .B(n_12122), .C(n_56301), .D(n_12034), .Z(n_1238
		));
	notech_reg_set tab22_reg_19(.CP(n_63062), .D(n_10113), .SD(n_62328), .Q(\tab22[19] 
		));
	notech_mux2 i_11620(.S(n_56159), .A(\tab22[19] ), .B(n_56741), .Z(n_10113
		));
	notech_reg_set tab22_reg_20(.CP(n_63066), .D(n_10119), .SD(n_62332), .Q(\tab22[20] 
		));
	notech_mux2 i_11628(.S(n_56159), .A(\tab22[20] ), .B(n_56747), .Z(n_10119
		));
	notech_ao4 i_738(.A(n_1086), .B(n_11900), .C(n_1084), .D(n_11929), .Z(n_1240
		));
	notech_reg_set tab22_reg_21(.CP(n_63070), .D(n_10125), .SD(n_62336), .Q(\tab22[21] 
		));
	notech_mux2 i_11636(.S(n_56159), .A(\tab22[21] ), .B(n_56753), .Z(n_10125
		));
	notech_reg_set tab22_reg_22(.CP(n_63070), .D(n_10131), .SD(n_62336), .Q(\tab22[22] 
		));
	notech_mux2 i_11644(.S(n_56159), .A(\tab22[22] ), .B(n_56759), .Z(n_10131
		));
	notech_ao4 i_736(.A(n_1092), .B(n_11950), .C(n_1090), .D(n_11970), .Z(n_1242
		));
	notech_reg_set tab22_reg_23(.CP(n_63070), .D(n_10137), .SD(n_62336), .Q(\tab22[23] 
		));
	notech_mux2 i_11652(.S(n_56159), .A(\tab22[23] ), .B(n_56765), .Z(n_10137
		));
	notech_reg_set tab22_reg_24(.CP(n_63070), .D(n_10143), .SD(n_62336), .Q(\tab22[24] 
		));
	notech_mux2 i_11660(.S(n_56159), .A(\tab22[24] ), .B(n_56771), .Z(n_10143
		));
	notech_and4 i_740(.A(n_1242), .B(n_1240), .C(n_721), .D(n_724), .Z(n_1244
		));
	notech_reg_set tab22_reg_25(.CP(n_63070), .D(n_10149), .SD(n_62336), .Q(\tab22[25] 
		));
	notech_mux2 i_11668(.S(n_56159), .A(\tab22[25] ), .B(n_56777), .Z(n_10149
		));
	notech_ao4 i_733(.A(n_1100), .B(n_11876), .C(n_55393), .D(n_12031), .Z(n_1245
		));
	notech_reg_set tab22_reg_26(.CP(n_63069), .D(n_10155), .SD(n_62335), .Q(\tab22[26] 
		));
	notech_mux2 i_11676(.S(n_56159), .A(\tab22[26] ), .B(n_56783), .Z(n_10155
		));
	notech_reg_set tab22_reg_27(.CP(n_63069), .D(n_10161), .SD(n_62335), .Q(\tab22[27] 
		));
	notech_mux2 i_11684(.S(\nbus_14520[0] ), .A(\tab22[27] ), .B(n_56789), .Z
		(n_10161));
	notech_ao4 i_732(.A(n_62898), .B(n_12121), .C(n_1043), .D(n_12032), .Z(n_1247
		));
	notech_reg_set tab22_reg_28(.CP(n_63069), .D(n_10167), .SD(n_62335), .Q(\tab22[28] 
		));
	notech_mux2 i_11692(.S(n_56159), .A(\tab22[28] ), .B(n_56795), .Z(n_10167
		));
	notech_reg_set tab22_reg_29(.CP(n_63069), .D(n_10173), .SD(n_62335), .Q(\tab22[29] 
		));
	notech_mux2 i_11700(.S(n_56159), .A(\tab22[29] ), .B(n_56801), .Z(n_10173
		));
	notech_ao4 i_729(.A(n_1086), .B(n_11899), .C(n_1084), .D(n_11928), .Z(n_1249
		));
	notech_reg tab22_reg_30(.CP(n_63071), .D(n_10179), .CD(n_62337), .Q(\tab22[30] 
		));
	notech_mux2 i_11708(.S(n_56159), .A(\tab22[30] ), .B(n_974), .Z(n_10179)
		);
	notech_reg tab22_reg_32(.CP(n_63070), .D(n_10185), .CD(n_62336), .Q(\tab22[32] 
		));
	notech_mux2 i_11716(.S(n_56159), .A(\tab22[32] ), .B(n_975), .Z(n_10185)
		);
	notech_ao4 i_727(.A(n_1092), .B(n_11949), .C(n_1090), .D(n_11969), .Z(n_1251
		));
	notech_reg_set tab22_reg_33(.CP(n_63071), .D(n_10191), .SD(n_62337), .Q(\tab22[33] 
		));
	notech_mux2 i_11724(.S(n_56159), .A(\tab22[33] ), .B(n_56153), .Z(n_10191
		));
	notech_reg hit_adr22_reg(.CP(n_63071), .D(n_10197), .CD(n_62337), .Q(hit_adr22
		));
	notech_mux2 i_11732(.S(n_971), .A(hit_add22), .B(hit_adr22), .Z(n_10197)
		);
	notech_and4 i_731(.A(n_1251), .B(n_1249), .C(n_710), .D(n_713), .Z(n_1253
		));
	notech_reg_set tab23_reg_0(.CP(n_63070), .D(n_10203), .SD(n_62336), .Q(\tab23[0] 
		));
	notech_mux2 i_11740(.S(\nbus_14502[0] ), .A(\tab23[0] ), .B(n_56627), .Z
		(n_10203));
	notech_ao4 i_724(.A(n_1100), .B(n_11875), .C(n_55393), .D(n_12029), .Z(n_1254
		));
	notech_reg_set tab23_reg_1(.CP(n_63070), .D(n_10209), .SD(n_62336), .Q(\tab23[1] 
		));
	notech_mux2 i_11748(.S(\nbus_14502[0] ), .A(\tab23[1] ), .B(n_56633), .Z
		(n_10209));
	notech_reg_set tab23_reg_2(.CP(n_63070), .D(n_10215), .SD(n_62336), .Q(\tab23[2] 
		));
	notech_mux2 i_11756(.S(\nbus_14502[0] ), .A(\tab23[2] ), .B(n_56639), .Z
		(n_10215));
	notech_ao4 i_723(.A(n_62898), .B(n_12120), .C(n_56301), .D(n_12030), .Z(n_1256
		));
	notech_reg_set tab23_reg_3(.CP(n_63070), .D(n_10221), .SD(n_62336), .Q(\tab23[3] 
		));
	notech_mux2 i_11764(.S(\nbus_14502[0] ), .A(\tab23[3] ), .B(n_56645), .Z
		(n_10221));
	notech_reg tab23_reg_4(.CP(n_63070), .D(n_10227), .CD(n_62336), .Q(\tab23[4] 
		));
	notech_mux2 i_11772(.S(\nbus_14502[0] ), .A(\tab23[4] ), .B(n_973), .Z(n_10227
		));
	notech_ao4 i_720(.A(n_1086), .B(n_11898), .C(n_1084), .D(n_11927), .Z(n_1258
		));
	notech_reg_set tab23_reg_5(.CP(n_63067), .D(n_10233), .SD(n_62333), .Q(\tab23[5] 
		));
	notech_mux2 i_11780(.S(\nbus_14502[0] ), .A(\tab23[5] ), .B(n_56657), .Z
		(n_10233));
	notech_reg_set tab23_reg_6(.CP(n_63067), .D(n_10239), .SD(n_62333), .Q(\tab23[6] 
		));
	notech_mux2 i_11788(.S(\nbus_14502[0] ), .A(\tab23[6] ), .B(n_56663), .Z
		(n_10239));
	notech_ao4 i_718(.A(n_1092), .B(n_11948), .C(n_1090), .D(n_11968), .Z(n_1260
		));
	notech_reg_set tab23_reg_7(.CP(n_63067), .D(n_10245), .SD(n_62333), .Q(\tab23[7] 
		));
	notech_mux2 i_11796(.S(\nbus_14502[0] ), .A(\tab23[7] ), .B(n_56669), .Z
		(n_10245));
	notech_reg_set tab23_reg_8(.CP(n_63067), .D(n_10251), .SD(n_62333), .Q(\tab23[8] 
		));
	notech_mux2 i_11804(.S(\nbus_14502[0] ), .A(\tab23[8] ), .B(n_56675), .Z
		(n_10251));
	notech_and4 i_722(.A(n_1260), .B(n_1258), .C(n_699), .D(n_702), .Z(n_1262
		));
	notech_reg_set tab23_reg_9(.CP(n_63067), .D(n_10257), .SD(n_62333), .Q(\tab23[9] 
		));
	notech_mux2 i_11812(.S(\nbus_14502[0] ), .A(\tab23[9] ), .B(n_56681), .Z
		(n_10257));
	notech_ao4 i_715(.A(n_1100), .B(n_11874), .C(n_55393), .D(n_12027), .Z(n_1263
		));
	notech_reg_set tab23_reg_10(.CP(n_63067), .D(n_10263), .SD(n_62333), .Q(\tab23[10] 
		));
	notech_mux2 i_11820(.S(\nbus_14502[0] ), .A(\tab23[10] ), .B(n_56687), .Z
		(n_10263));
	notech_reg_set tab23_reg_11(.CP(n_63067), .D(n_10269), .SD(n_62333), .Q(\tab23[11] 
		));
	notech_mux2 i_11828(.S(\nbus_14502[0] ), .A(\tab23[11] ), .B(n_56693), .Z
		(n_10269));
	notech_ao4 i_714(.A(n_62898), .B(n_12119), .C(n_56301), .D(n_12028), .Z(n_1265
		));
	notech_reg_set tab23_reg_12(.CP(n_63067), .D(n_10275), .SD(n_62333), .Q(\tab23[12] 
		));
	notech_mux2 i_11836(.S(\nbus_14502[0] ), .A(\tab23[12] ), .B(n_56699), .Z
		(n_10275));
	notech_reg_set tab23_reg_13(.CP(n_63067), .D(n_10281), .SD(n_62333), .Q(\tab23[13] 
		));
	notech_mux2 i_11844(.S(\nbus_14502[0] ), .A(\tab23[13] ), .B(n_56705), .Z
		(n_10281));
	notech_ao4 i_711(.A(n_1086), .B(n_11897), .C(n_1084), .D(n_11926), .Z(n_1267
		));
	notech_reg_set tab23_reg_14(.CP(n_63069), .D(n_10287), .SD(n_62335), .Q(\tab23[14] 
		));
	notech_mux2 i_11852(.S(\nbus_14502[0] ), .A(\tab23[14] ), .B(n_56711), .Z
		(n_10287));
	notech_reg_set tab23_reg_15(.CP(n_63069), .D(n_10293), .SD(n_62335), .Q(\tab23[15] 
		));
	notech_mux2 i_11860(.S(\nbus_14502[0] ), .A(\tab23[15] ), .B(n_56717), .Z
		(n_10293));
	notech_ao4 i_709(.A(n_1092), .B(n_11947), .C(n_1090), .D(n_11967), .Z(n_1269
		));
	notech_reg_set tab23_reg_16(.CP(n_63069), .D(n_10299), .SD(n_62335), .Q(\tab23[16] 
		));
	notech_mux2 i_11868(.S(\nbus_14502[0] ), .A(\tab23[16] ), .B(n_56723), .Z
		(n_10299));
	notech_reg_set tab23_reg_17(.CP(n_63069), .D(n_10305), .SD(n_62335), .Q(\tab23[17] 
		));
	notech_mux2 i_11876(.S(n_56121), .A(\tab23[17] ), .B(n_56729), .Z(n_10305
		));
	notech_and4 i_713(.A(n_1269), .B(n_1267), .C(n_691), .D(n_688), .Z(n_1271
		));
	notech_reg_set tab23_reg_18(.CP(n_63069), .D(n_10311), .SD(n_62335), .Q(\tab23[18] 
		));
	notech_mux2 i_11884(.S(n_56121), .A(\tab23[18] ), .B(n_56735), .Z(n_10311
		));
	notech_ao4 i_706(.A(n_1100), .B(n_11873), .C(n_55393), .D(n_12025), .Z(n_1272
		));
	notech_reg_set tab23_reg_19(.CP(n_63067), .D(n_10317), .SD(n_62333), .Q(\tab23[19] 
		));
	notech_mux2 i_11892(.S(n_56121), .A(\tab23[19] ), .B(n_56741), .Z(n_10317
		));
	notech_reg_set tab23_reg_20(.CP(n_63067), .D(n_10323), .SD(n_62333), .Q(\tab23[20] 
		));
	notech_mux2 i_11900(.S(n_56121), .A(\tab23[20] ), .B(n_56747), .Z(n_10323
		));
	notech_ao4 i_705(.A(n_62898), .B(n_12118), .C(n_56301), .D(n_12026), .Z(n_1274
		));
	notech_reg_set tab23_reg_21(.CP(n_63069), .D(n_10329), .SD(n_62335), .Q(\tab23[21] 
		));
	notech_mux2 i_11908(.S(n_56121), .A(\tab23[21] ), .B(n_56753), .Z(n_10329
		));
	notech_reg_set tab23_reg_22(.CP(n_63069), .D(n_10335), .SD(n_62335), .Q(\tab23[22] 
		));
	notech_mux2 i_11916(.S(n_56121), .A(\tab23[22] ), .B(n_56759), .Z(n_10335
		));
	notech_ao4 i_704(.A(n_55393), .B(n_12024), .C(n_486), .D(n_12117), .Z(n_1276
		));
	notech_reg_set tab23_reg_23(.CP(n_63041), .D(n_10341), .SD(n_62307), .Q(\tab23[23] 
		));
	notech_mux2 i_11924(.S(n_56121), .A(\tab23[23] ), .B(n_56765), .Z(n_10341
		));
	notech_ao4 i_703(.A(n_55393), .B(n_12023), .C(n_486), .D(n_12116), .Z(n_1277
		));
	notech_reg_set tab23_reg_24(.CP(n_63013), .D(n_10347), .SD(n_62279), .Q(\tab23[24] 
		));
	notech_mux2 i_11932(.S(n_56121), .A(\tab23[24] ), .B(n_56771), .Z(n_10347
		));
	notech_ao4 i_702(.A(n_55393), .B(n_12022), .C(n_486), .D(n_12115), .Z(n_1278
		));
	notech_reg_set tab23_reg_25(.CP(n_63013), .D(n_10353), .SD(n_62279), .Q(\tab23[25] 
		));
	notech_mux2 i_11940(.S(n_56121), .A(\tab23[25] ), .B(n_56777), .Z(n_10353
		));
	notech_ao4 i_701(.A(n_55393), .B(n_12021), .C(n_486), .D(n_12114), .Z(n_1279
		));
	notech_reg_set tab23_reg_26(.CP(n_63013), .D(n_10359), .SD(n_62279), .Q(\tab23[26] 
		));
	notech_mux2 i_11948(.S(n_56121), .A(\tab23[26] ), .B(n_56783), .Z(n_10359
		));
	notech_ao4 i_700(.A(n_55393), .B(n_12020), .C(n_486), .D(n_12113), .Z(n_1280
		));
	notech_reg_set tab23_reg_27(.CP(n_63013), .D(n_10365), .SD(n_62279), .Q(\tab23[27] 
		));
	notech_mux2 i_11956(.S(\nbus_14502[0] ), .A(\tab23[27] ), .B(n_56789), .Z
		(n_10365));
	notech_ao4 i_699(.A(n_55393), .B(n_12019), .C(n_486), .D(n_12112), .Z(n_1281
		));
	notech_reg_set tab23_reg_28(.CP(n_63013), .D(n_10371), .SD(n_62279), .Q(\tab23[28] 
		));
	notech_mux2 i_11964(.S(n_56121), .A(\tab23[28] ), .B(n_56795), .Z(n_10371
		));
	notech_ao4 i_698(.A(n_1098), .B(n_12018), .C(n_486), .D(n_12111), .Z(n_1282
		));
	notech_reg_set tab23_reg_29(.CP(n_63011), .D(n_10377), .SD(n_62277), .Q(\tab23[29] 
		));
	notech_mux2 i_11972(.S(n_56121), .A(\tab23[29] ), .B(n_56801), .Z(n_10377
		));
	notech_ao4 i_697(.A(n_55393), .B(n_12017), .C(n_486), .D(n_12110), .Z(n_1283
		));
	notech_reg tab23_reg_30(.CP(n_63011), .D(n_10383), .CD(n_62277), .Q(\tab23[30] 
		));
	notech_mux2 i_11980(.S(n_56121), .A(\tab23[30] ), .B(n_974), .Z(n_10383)
		);
	notech_ao4 i_696(.A(n_55393), .B(n_12016), .C(n_486), .D(n_12109), .Z(n_1284
		));
	notech_reg tab23_reg_32(.CP(n_63013), .D(n_10389), .CD(n_62279), .Q(\tab23[32] 
		));
	notech_mux2 i_11988(.S(n_56121), .A(\tab23[32] ), .B(n_975), .Z(n_10389)
		);
	notech_ao4 i_695(.A(n_55393), .B(n_12015), .C(n_486), .D(n_12108), .Z(n_1285
		));
	notech_reg_set tab23_reg_33(.CP(n_63013), .D(n_10395), .SD(n_62279), .Q(\tab23[33] 
		));
	notech_mux2 i_11996(.S(n_56121), .A(\tab23[33] ), .B(n_56153), .Z(n_10395
		));
	notech_ao4 i_694(.A(n_55393), .B(n_12014), .C(n_486), .D(n_12107), .Z(n_1286
		));
	notech_reg hit_adr23_reg(.CP(n_63014), .D(n_10401), .CD(n_62280), .Q(hit_adr23
		));
	notech_mux2 i_12004(.S(n_971), .A(hit_add23), .B(hit_adr23), .Z(n_10401)
		);
	notech_ao4 i_693(.A(n_55393), .B(n_12013), .C(n_486), .D(n_12106), .Z(n_1287
		));
	notech_reg_set tab24_reg_0(.CP(n_63014), .D(n_10407), .SD(n_62280), .Q(\tab24[0] 
		));
	notech_mux2 i_12012(.S(\nbus_14503[0] ), .A(\tab24[0] ), .B(n_56627), .Z
		(n_10407));
	notech_reg_set tab24_reg_1(.CP(n_63014), .D(n_10413), .SD(n_62280), .Q(\tab24[1] 
		));
	notech_mux2 i_12020(.S(\nbus_14503[0] ), .A(\tab24[1] ), .B(n_56633), .Z
		(n_10413));
	notech_ao4 i_79327(.A(n_62898), .B(n_12167), .C(n_986), .D(n_987), .Z(oread_ack101000
		));
	notech_reg_set tab24_reg_2(.CP(n_63014), .D(n_10419), .SD(n_62280), .Q(\tab24[2] 
		));
	notech_mux2 i_12028(.S(\nbus_14503[0] ), .A(\tab24[2] ), .B(n_56639), .Z
		(n_10419));
	notech_nand3 i_81704(.A(n_631), .B(n_628), .C(n_625), .Z(\nbus_14516[0] 
		));
	notech_reg_set tab24_reg_3(.CP(n_63014), .D(n_10425), .SD(n_62280), .Q(\tab24[3] 
		));
	notech_mux2 i_12036(.S(\nbus_14503[0] ), .A(\tab24[3] ), .B(n_56645), .Z
		(n_10425));
	notech_nao3 i_81813(.A(n_628), .B(n_625), .C(n_626), .Z(\nbus_14517[0] )
		);
	notech_reg tab24_reg_4(.CP(n_63013), .D(n_10431), .CD(n_62279), .Q(\tab24[4] 
		));
	notech_mux2 i_12044(.S(\nbus_14503[0] ), .A(\tab24[4] ), .B(n_973), .Z(n_10431
		));
	notech_nao3 i_81242(.A(n_628), .B(n_604), .C(n_626), .Z(\nbus_14511[0] )
		);
	notech_reg_set tab24_reg_5(.CP(n_63013), .D(n_10437), .SD(n_62279), .Q(\tab24[5] 
		));
	notech_mux2 i_12052(.S(\nbus_14503[0] ), .A(\tab24[5] ), .B(n_56657), .Z
		(n_10437));
	notech_nand3 i_80979(.A(n_631), .B(n_628), .C(n_601), .Z(\nbus_14508[0] 
		));
	notech_reg_set tab24_reg_6(.CP(n_63013), .D(n_10443), .SD(n_62279), .Q(\tab24[6] 
		));
	notech_mux2 i_12060(.S(\nbus_14503[0] ), .A(\tab24[6] ), .B(n_56663), .Z
		(n_10443));
	notech_nand3 i_80264(.A(n_631), .B(n_628), .C(n_600), .Z(\nbus_14492[0] 
		));
	notech_reg_set tab24_reg_7(.CP(n_63013), .D(n_10449), .SD(n_62279), .Q(\tab24[7] 
		));
	notech_mux2 i_12068(.S(\nbus_14503[0] ), .A(\tab24[7] ), .B(n_56669), .Z
		(n_10449));
	notech_nand3 i_79986(.A(n_631), .B(n_628), .C(n_599), .Z(\nbus_14489[0] 
		));
	notech_reg_set tab24_reg_8(.CP(n_63010), .D(n_10455), .SD(n_62276), .Q(\tab24[8] 
		));
	notech_mux2 i_12076(.S(\nbus_14503[0] ), .A(\tab24[8] ), .B(n_56675), .Z
		(n_10455));
	notech_nand2 i_81352(.A(n_1020), .B(n_1011), .Z(\nbus_14512[0] ));
	notech_reg_set tab24_reg_9(.CP(n_63010), .D(n_10461), .SD(n_62276), .Q(\tab24[9] 
		));
	notech_mux2 i_12084(.S(\nbus_14503[0] ), .A(\tab24[9] ), .B(n_56681), .Z
		(n_10461));
	notech_ao4 i_80960(.A(n_1001), .B(n_1010), .C(n_1020), .D(n_11881), .Z(\nbus_14507[0] 
		));
	notech_reg_set tab24_reg_10(.CP(n_63010), .D(n_10467), .SD(n_62276), .Q(\tab24[10] 
		));
	notech_mux2 i_12092(.S(\nbus_14503[0] ), .A(\tab24[10] ), .B(n_56687), .Z
		(n_10467));
	notech_nao3 i_81932(.A(n_628), .B(n_579), .C(n_626), .Z(\nbus_14520[0] )
		);
	notech_reg_set tab24_reg_11(.CP(n_63010), .D(n_10473), .SD(n_62276), .Q(\tab24[11] 
		));
	notech_mux2 i_12100(.S(\nbus_14503[0] ), .A(\tab24[11] ), .B(n_56693), .Z
		(n_10473));
	notech_nao3 i_80481(.A(n_628), .B(n_578), .C(n_626), .Z(\nbus_14502[0] )
		);
	notech_reg_set tab24_reg_12(.CP(n_63010), .D(n_10479), .SD(n_62276), .Q(\tab24[12] 
		));
	notech_mux2 i_12108(.S(\nbus_14503[0] ), .A(\tab24[12] ), .B(n_56699), .Z
		(n_10479));
	notech_nao3 i_80657(.A(n_628), .B(n_577), .C(n_626), .Z(\nbus_14503[0] )
		);
	notech_reg_set tab24_reg_13(.CP(n_63010), .D(n_10485), .SD(n_62276), .Q(\tab24[13] 
		));
	notech_mux2 i_12116(.S(\nbus_14503[0] ), .A(\tab24[13] ), .B(n_56705), .Z
		(n_10485));
	notech_ao4 i_80936(.A(n_1002), .B(n_1001), .C(n_1020), .D(n_11872), .Z(\nbus_14506[0] 
		));
	notech_reg_set tab24_reg_14(.CP(n_63010), .D(n_10491), .SD(n_62276), .Q(\tab24[14] 
		));
	notech_mux2 i_12124(.S(\nbus_14503[0] ), .A(\tab24[14] ), .B(n_56711), .Z
		(n_10491));
	notech_nand2 i_81672(.A(n_1020), .B(n_1003), .Z(\nbus_14515[0] ));
	notech_reg_set tab24_reg_15(.CP(n_63010), .D(n_10497), .SD(n_62276), .Q(\tab24[15] 
		));
	notech_mux2 i_12132(.S(\nbus_14503[0] ), .A(\tab24[15] ), .B(n_56717), .Z
		(n_10497));
	notech_nand3 i_81130(.A(n_631), .B(n_628), .C(n_557), .Z(\nbus_14510[0] 
		));
	notech_reg_set tab24_reg_16(.CP(n_63010), .D(n_10503), .SD(n_62276), .Q(\tab24[16] 
		));
	notech_mux2 i_12140(.S(\nbus_14503[0] ), .A(\tab24[16] ), .B(n_56723), .Z
		(n_10503));
	notech_nand2 i_80886(.A(n_992), .B(n_552), .Z(\nbus_14505[0] ));
	notech_reg_set tab24_reg_17(.CP(n_63011), .D(n_10509), .SD(n_62277), .Q(\tab24[17] 
		));
	notech_mux2 i_12148(.S(n_56139), .A(\tab24[17] ), .B(n_56729), .Z(n_10509
		));
	notech_or2 i_85(.A(n_409), .B(n_11866), .Z(n_56850));
	notech_reg_set tab24_reg_18(.CP(n_63011), .D(n_10515), .SD(n_62277), .Q(\tab24[18] 
		));
	notech_mux2 i_12156(.S(n_56139), .A(\tab24[18] ), .B(n_56735), .Z(n_10515
		));
	notech_or4 i_81101(.A(n_409), .B(\nbus_14514[0] ), .C(n_1048), .D(n_11866
		), .Z(\nbus_14509[0] ));
	notech_reg_set tab24_reg_19(.CP(n_63011), .D(n_10521), .SD(n_62277), .Q(\tab24[19] 
		));
	notech_mux2 i_12164(.S(n_56139), .A(\tab24[19] ), .B(n_56741), .Z(n_10521
		));
	notech_ao4 i_68(.A(data_miss[0]), .B(n_989), .C(n_996), .D(n_11845), .Z(n_56853
		));
	notech_reg_set tab24_reg_20(.CP(n_63011), .D(n_10527), .SD(n_62277), .Q(\tab24[20] 
		));
	notech_mux2 i_12172(.S(n_56139), .A(\tab24[20] ), .B(n_56747), .Z(n_10527
		));
	notech_nand2 i_87(.A(n_1020), .B(n_545), .Z(\nbus_14514[0] ));
	notech_reg_set tab24_reg_21(.CP(n_63011), .D(n_10533), .SD(n_62277), .Q(\tab24[21] 
		));
	notech_mux2 i_12180(.S(n_56139), .A(\tab24[21] ), .B(n_56753), .Z(n_10533
		));
	notech_reg_set tab24_reg_22(.CP(n_63011), .D(n_10539), .SD(n_62277), .Q(\tab24[22] 
		));
	notech_mux2 i_12188(.S(n_56139), .A(\tab24[22] ), .B(n_56759), .Z(n_10539
		));
	notech_ao4 i_86(.A(n_1001), .B(n_550), .C(data_miss[5]), .D(n_977), .Z(\nbus_14488[0] 
		));
	notech_reg_set tab24_reg_23(.CP(n_63011), .D(n_10545), .SD(n_62277), .Q(\tab24[23] 
		));
	notech_mux2 i_12196(.S(n_56139), .A(\tab24[23] ), .B(n_56765), .Z(n_10545
		));
	notech_or2 i_80092(.A(n_409), .B(n_410), .Z(n_56836));
	notech_reg_set tab24_reg_24(.CP(n_63011), .D(n_10551), .SD(n_62277), .Q(\tab24[24] 
		));
	notech_mux2 i_12204(.S(n_56139), .A(\tab24[24] ), .B(n_56771), .Z(n_10551
		));
	notech_mux2 i_122908(.S(n_948), .A(iDaddr[12]), .B(iDaddr_f[12]), .Z(\tab11_0[0] 
		));
	notech_reg_set tab24_reg_25(.CP(n_63011), .D(n_10557), .SD(n_62277), .Q(\tab24[25] 
		));
	notech_mux2 i_12212(.S(n_56139), .A(\tab24[25] ), .B(n_56777), .Z(n_10557
		));
	notech_mux2 i_222909(.S(n_948), .A(iDaddr[13]), .B(iDaddr_f[13]), .Z(\tab11_0[1] 
		));
	notech_reg_set tab24_reg_26(.CP(n_63014), .D(n_10563), .SD(n_62280), .Q(\tab24[26] 
		));
	notech_mux2 i_12220(.S(n_56139), .A(\tab24[26] ), .B(n_56783), .Z(n_10563
		));
	notech_mux2 i_322910(.S(n_948), .A(iDaddr[14]), .B(iDaddr_f[14]), .Z(\tab11_0[2] 
		));
	notech_reg_set tab24_reg_27(.CP(n_63018), .D(n_10569), .SD(n_62284), .Q(\tab24[27] 
		));
	notech_mux2 i_12228(.S(\nbus_14503[0] ), .A(\tab24[27] ), .B(n_56789), .Z
		(n_10569));
	notech_mux2 i_422911(.S(n_948), .A(iDaddr[15]), .B(iDaddr_f[15]), .Z(\tab11_0[3] 
		));
	notech_reg_set tab24_reg_28(.CP(n_63018), .D(n_10575), .SD(n_62284), .Q(\tab24[28] 
		));
	notech_mux2 i_12236(.S(n_56139), .A(\tab24[28] ), .B(n_56795), .Z(n_10575
		));
	notech_mux2 i_522912(.S(n_948), .A(iDaddr[16]), .B(iDaddr_f[16]), .Z(\tab11_0[4] 
		));
	notech_reg_set tab24_reg_29(.CP(n_63018), .D(n_10581), .SD(n_62284), .Q(\tab24[29] 
		));
	notech_mux2 i_12244(.S(n_56139), .A(\tab24[29] ), .B(n_56801), .Z(n_10581
		));
	notech_mux2 i_622913(.S(n_58743), .A(iDaddr[17]), .B(iDaddr_f[17]), .Z(\tab11_0[5] 
		));
	notech_reg tab24_reg_30(.CP(n_63018), .D(n_10587), .CD(n_62284), .Q(\tab24[30] 
		));
	notech_mux2 i_12252(.S(n_56139), .A(\tab24[30] ), .B(n_974), .Z(n_10587)
		);
	notech_mux2 i_722914(.S(n_58743), .A(iDaddr[18]), .B(iDaddr_f[18]), .Z(\tab11_0[6] 
		));
	notech_reg tab24_reg_32(.CP(n_63018), .D(n_10593), .CD(n_62284), .Q(\tab24[32] 
		));
	notech_mux2 i_12260(.S(n_56139), .A(\tab24[32] ), .B(n_975), .Z(n_10593)
		);
	notech_mux2 i_822915(.S(n_58743), .A(iDaddr[19]), .B(iDaddr_f[19]), .Z(\tab11_0[7] 
		));
	notech_reg_set tab24_reg_33(.CP(n_63018), .D(n_10599), .SD(n_62284), .Q(\tab24[33] 
		));
	notech_mux2 i_12268(.S(n_56139), .A(\tab24[33] ), .B(n_56153), .Z(n_10599
		));
	notech_mux2 i_922916(.S(n_58743), .A(iDaddr[20]), .B(iDaddr_f[20]), .Z(\tab11_0[8] 
		));
	notech_reg hit_adr24_reg(.CP(n_63018), .D(n_10605), .CD(n_62284), .Q(hit_adr24
		));
	notech_mux2 i_12276(.S(n_971), .A(hit_add24), .B(hit_adr24), .Z(n_10605)
		);
	notech_mux2 i_1022917(.S(n_58743), .A(iDaddr[21]), .B(iDaddr_f[21]), .Z(\tab11_0[9] 
		));
	notech_reg_set nnx_tab2_reg_0(.CP(n_63018), .D(n_10611), .SD(n_62284), .Q
		(\nnx_tab2[0] ));
	notech_mux2 i_12284(.S(n_11991), .A(\nnx_tab2[0] ), .B(n_11987), .Z(n_10611
		));
	notech_mux2 i_1122918(.S(n_58743), .A(iDaddr[22]), .B(iDaddr_f[22]), .Z(\dir1_0[0] 
		));
	notech_reg nnx_tab2_reg_1(.CP(n_63018), .D(n_10617), .CD(n_62284), .Q(\nnx_tab2[1] 
		));
	notech_mux2 i_12292(.S(n_11991), .A(\nnx_tab2[1] ), .B(n_11989), .Z(n_10617
		));
	notech_mux2 i_1222919(.S(n_58743), .A(iDaddr[23]), .B(iDaddr_f[23]), .Z(\dir1_0[1] 
		));
	notech_reg nx_tab2_reg_0(.CP(n_63019), .D(n_10623), .CD(n_62285), .Q(\nx_tab2[0] 
		));
	notech_mux2 i_12300(.S(\nbus_14515[0] ), .A(\nx_tab2[0] ), .B(n_11992), 
		.Z(n_10623));
	notech_mux2 i_1322920(.S(n_58743), .A(iDaddr[24]), .B(iDaddr_f[24]), .Z(\dir1_0[2] 
		));
	notech_reg nx_tab2_reg_1(.CP(n_63019), .D(n_10629), .CD(n_62285), .Q(\nx_tab2[1] 
		));
	notech_mux2 i_12308(.S(\nbus_14515[0] ), .A(\nx_tab2[1] ), .B(n_11994), 
		.Z(n_10629));
	notech_mux2 i_1422921(.S(n_58743), .A(iDaddr[25]), .B(iDaddr_f[25]), .Z(\dir1_0[3] 
		));
	notech_reg_set tab11_reg_0(.CP(n_63019), .D(n_10635), .SD(n_62285), .Q(\tab11[0] 
		));
	notech_mux2 i_12316(.S(\nbus_14510[0] ), .A(\tab11[0] ), .B(n_56627), .Z
		(n_10635));
	notech_mux2 i_1522922(.S(n_58743), .A(iDaddr[26]), .B(iDaddr_f[26]), .Z(\dir1_0[4] 
		));
	notech_reg_set tab11_reg_1(.CP(n_63019), .D(n_10641), .SD(n_62285), .Q(\tab11[1] 
		));
	notech_mux2 i_12324(.S(\nbus_14510[0] ), .A(\tab11[1] ), .B(n_56633), .Z
		(n_10641));
	notech_mux2 i_1622923(.S(n_58743), .A(iDaddr[27]), .B(iDaddr_f[27]), .Z(\dir1_0[5] 
		));
	notech_reg_set tab11_reg_2(.CP(n_63019), .D(n_10647), .SD(n_62285), .Q(\tab11[2] 
		));
	notech_mux2 i_12332(.S(\nbus_14510[0] ), .A(\tab11[2] ), .B(n_56639), .Z
		(n_10647));
	notech_mux2 i_1722924(.S(n_948), .A(iDaddr[28]), .B(iDaddr_f[28]), .Z(\dir1_0[6] 
		));
	notech_reg_set tab11_reg_3(.CP(n_63019), .D(n_10653), .SD(n_62285), .Q(\tab11[3] 
		));
	notech_mux2 i_12340(.S(\nbus_14510[0] ), .A(\tab11[3] ), .B(n_56645), .Z
		(n_10653));
	notech_mux2 i_1822925(.S(n_58743), .A(iDaddr[29]), .B(iDaddr_f[29]), .Z(\dir1_0[7] 
		));
	notech_reg tab11_reg_4(.CP(n_63019), .D(n_10659), .CD(n_62285), .Q(\tab11[4] 
		));
	notech_mux2 i_12348(.S(\nbus_14510[0] ), .A(\tab11[4] ), .B(n_973), .Z(n_10659
		));
	notech_mux2 i_1922926(.S(n_58743), .A(iDaddr[30]), .B(iDaddr_f[30]), .Z(\dir1_0[8] 
		));
	notech_reg_set tab11_reg_5(.CP(n_63019), .D(n_10665), .SD(n_62285), .Q(\tab11[5] 
		));
	notech_mux2 i_12356(.S(\nbus_14510[0] ), .A(\tab11[5] ), .B(n_56657), .Z
		(n_10665));
	notech_mux2 i_2022927(.S(n_58743), .A(iDaddr[31]), .B(iDaddr_f[31]), .Z(\dir1_0[9] 
		));
	notech_reg_set tab11_reg_6(.CP(n_63019), .D(n_10671), .SD(n_62285), .Q(\tab11[6] 
		));
	notech_mux2 i_12364(.S(\nbus_14510[0] ), .A(\tab11[6] ), .B(n_56663), .Z
		(n_10671));
	notech_mux2 i_122429(.S(n_55416), .A(wrD[0]), .B(iwrite_data[0]), .Z(n_57299
		));
	notech_reg_set tab11_reg_7(.CP(n_63015), .D(n_10677), .SD(n_62281), .Q(\tab11[7] 
		));
	notech_mux2 i_12372(.S(\nbus_14510[0] ), .A(\tab11[7] ), .B(n_56669), .Z
		(n_10677));
	notech_mux2 i_222430(.S(n_55416), .A(wrD[1]), .B(iwrite_data[1]), .Z(n_57306
		));
	notech_reg_set tab11_reg_8(.CP(n_63015), .D(n_10683), .SD(n_62281), .Q(\tab11[8] 
		));
	notech_mux2 i_12380(.S(\nbus_14510[0] ), .A(\tab11[8] ), .B(n_56675), .Z
		(n_10683));
	notech_mux2 i_322431(.S(n_55416), .A(wrD[2]), .B(iwrite_data[2]), .Z(n_57313
		));
	notech_reg_set tab11_reg_9(.CP(n_63015), .D(n_10689), .SD(n_62281), .Q(\tab11[9] 
		));
	notech_mux2 i_12388(.S(\nbus_14510[0] ), .A(\tab11[9] ), .B(n_56681), .Z
		(n_10689));
	notech_mux2 i_422432(.S(n_55416), .A(wrD[3]), .B(iwrite_data[3]), .Z(n_57320
		));
	notech_reg_set tab11_reg_10(.CP(n_63015), .D(n_10695), .SD(n_62281), .Q(\tab11[10] 
		));
	notech_mux2 i_12396(.S(\nbus_14510[0] ), .A(\tab11[10] ), .B(n_56687), .Z
		(n_10695));
	notech_mux2 i_522433(.S(n_55416), .A(wrD[4]), .B(iwrite_data[4]), .Z(n_57327
		));
	notech_reg_set tab11_reg_11(.CP(n_63014), .D(n_10701), .SD(n_62280), .Q(\tab11[11] 
		));
	notech_mux2 i_12404(.S(\nbus_14510[0] ), .A(\tab11[11] ), .B(n_56693), .Z
		(n_10701));
	notech_mux2 i_622434(.S(n_55416), .A(wrD[5]), .B(iwrite_data[5]), .Z(n_57334
		));
	notech_reg_set tab11_reg_12(.CP(n_63014), .D(n_10707), .SD(n_62280), .Q(\tab11[12] 
		));
	notech_mux2 i_12412(.S(\nbus_14510[0] ), .A(\tab11[12] ), .B(n_56699), .Z
		(n_10707));
	notech_mux2 i_722435(.S(n_55416), .A(wrD[6]), .B(iwrite_data[6]), .Z(n_57341
		));
	notech_reg_set tab11_reg_13(.CP(n_63014), .D(n_10713), .SD(n_62280), .Q(\tab11[13] 
		));
	notech_mux2 i_12420(.S(\nbus_14510[0] ), .A(\tab11[13] ), .B(n_56705), .Z
		(n_10713));
	notech_mux2 i_822436(.S(n_55416), .A(wrD[7]), .B(iwrite_data[7]), .Z(n_57348
		));
	notech_reg_set tab11_reg_14(.CP(n_63014), .D(n_10719), .SD(n_62280), .Q(\tab11[14] 
		));
	notech_mux2 i_12428(.S(\nbus_14510[0] ), .A(\tab11[14] ), .B(n_56711), .Z
		(n_10719));
	notech_mux2 i_922437(.S(n_55416), .A(wrD[8]), .B(iwrite_data[8]), .Z(n_57355
		));
	notech_reg_set tab11_reg_15(.CP(n_63014), .D(n_10725), .SD(n_62280), .Q(\tab11[15] 
		));
	notech_mux2 i_12436(.S(\nbus_14510[0] ), .A(\tab11[15] ), .B(n_56717), .Z
		(n_10725));
	notech_mux2 i_1022438(.S(n_55416), .A(wrD[9]), .B(iwrite_data[9]), .Z(n_57362
		));
	notech_reg_set tab11_reg_16(.CP(n_63015), .D(n_10731), .SD(n_62281), .Q(\tab11[16] 
		));
	notech_mux2 i_12444(.S(\nbus_14510[0] ), .A(\tab11[16] ), .B(n_56723), .Z
		(n_10731));
	notech_mux2 i_1122439(.S(n_55416), .A(wrD[10]), .B(iwrite_data[10]), .Z(n_57369
		));
	notech_reg_set tab11_reg_17(.CP(n_63015), .D(n_10737), .SD(n_62281), .Q(\tab11[17] 
		));
	notech_mux2 i_12452(.S(n_56092), .A(\tab11[17] ), .B(n_56729), .Z(n_10737
		));
	notech_mux2 i_1222440(.S(n_55416), .A(wrD[11]), .B(iwrite_data[11]), .Z(n_57376
		));
	notech_reg_set tab11_reg_18(.CP(n_63018), .D(n_10743), .SD(n_62284), .Q(\tab11[18] 
		));
	notech_mux2 i_12460(.S(n_56092), .A(\tab11[18] ), .B(n_56735), .Z(n_10743
		));
	notech_mux2 i_1322441(.S(n_55416), .A(wrD[12]), .B(iwrite_data[12]), .Z(n_57383
		));
	notech_reg_set tab11_reg_19(.CP(n_63018), .D(n_10749), .SD(n_62284), .Q(\tab11[19] 
		));
	notech_mux2 i_12468(.S(n_56092), .A(\tab11[19] ), .B(n_56741), .Z(n_10749
		));
	notech_mux2 i_1422442(.S(n_55416), .A(wrD[13]), .B(iwrite_data[13]), .Z(n_57390
		));
	notech_reg_set tab11_reg_20(.CP(n_63015), .D(n_10755), .SD(n_62281), .Q(\tab11[20] 
		));
	notech_mux2 i_12476(.S(n_56092), .A(\tab11[20] ), .B(n_56747), .Z(n_10755
		));
	notech_mux2 i_1522443(.S(n_55416), .A(wrD[14]), .B(iwrite_data[14]), .Z(n_57397
		));
	notech_reg_set tab11_reg_21(.CP(n_63015), .D(n_10761), .SD(n_62281), .Q(\tab11[21] 
		));
	notech_mux2 i_12484(.S(n_56092), .A(\tab11[21] ), .B(n_56753), .Z(n_10761
		));
	notech_mux2 i_1622444(.S(n_55411), .A(wrD[15]), .B(iwrite_data[15]), .Z(n_57404
		));
	notech_reg_set tab11_reg_22(.CP(n_63015), .D(n_10767), .SD(n_62281), .Q(\tab11[22] 
		));
	notech_mux2 i_12492(.S(n_56092), .A(\tab11[22] ), .B(n_56759), .Z(n_10767
		));
	notech_mux2 i_1722445(.S(n_55411), .A(wrD[16]), .B(iwrite_data[16]), .Z(n_57411
		));
	notech_reg_set tab11_reg_23(.CP(n_63015), .D(n_10773), .SD(n_62281), .Q(\tab11[23] 
		));
	notech_mux2 i_12500(.S(n_56092), .A(\tab11[23] ), .B(n_56765), .Z(n_10773
		));
	notech_mux2 i_1822446(.S(n_55411), .A(wrD[17]), .B(iwrite_data[17]), .Z(n_57418
		));
	notech_reg_set tab11_reg_24(.CP(n_63015), .D(n_10779), .SD(n_62281), .Q(\tab11[24] 
		));
	notech_mux2 i_12508(.S(n_56092), .A(\tab11[24] ), .B(n_56771), .Z(n_10779
		));
	notech_mux2 i_1922447(.S(n_55411), .A(wrD[18]), .B(iwrite_data[18]), .Z(n_57425
		));
	notech_reg_set tab11_reg_25(.CP(n_63010), .D(n_10785), .SD(n_62276), .Q(\tab11[25] 
		));
	notech_mux2 i_12516(.S(n_56092), .A(\tab11[25] ), .B(n_56777), .Z(n_10785
		));
	notech_mux2 i_2022448(.S(n_55411), .A(wrD[19]), .B(iwrite_data[19]), .Z(n_57432
		));
	notech_reg_set tab11_reg_26(.CP(n_63001), .D(n_10791), .SD(n_62267), .Q(\tab11[26] 
		));
	notech_mux2 i_12524(.S(n_56092), .A(\tab11[26] ), .B(n_56783), .Z(n_10791
		));
	notech_mux2 i_2122449(.S(n_55411), .A(wrD[20]), .B(iwrite_data[20]), .Z(n_57439
		));
	notech_reg_set tab11_reg_27(.CP(n_63001), .D(n_10797), .SD(n_62267), .Q(\tab11[27] 
		));
	notech_mux2 i_12532(.S(\nbus_14510[0] ), .A(\tab11[27] ), .B(n_56789), .Z
		(n_10797));
	notech_mux2 i_2222450(.S(n_55411), .A(wrD[21]), .B(iwrite_data[21]), .Z(n_57446
		));
	notech_reg_set tab11_reg_28(.CP(n_63001), .D(n_10803), .SD(n_62267), .Q(\tab11[28] 
		));
	notech_mux2 i_12540(.S(n_56092), .A(\tab11[28] ), .B(n_56795), .Z(n_10803
		));
	notech_mux2 i_2322451(.S(n_55411), .A(wrD[22]), .B(iwrite_data[22]), .Z(n_57453
		));
	notech_reg_set tab11_reg_29(.CP(n_63001), .D(n_10809), .SD(n_62267), .Q(\tab11[29] 
		));
	notech_mux2 i_12548(.S(n_56092), .A(\tab11[29] ), .B(n_56801), .Z(n_10809
		));
	notech_mux2 i_2422452(.S(n_55411), .A(wrD[23]), .B(iwrite_data[23]), .Z(n_57460
		));
	notech_reg tab11_reg_30(.CP(n_63001), .D(n_10815), .CD(n_62267), .Q(\tab11[30] 
		));
	notech_mux2 i_12556(.S(n_56092), .A(\tab11[30] ), .B(n_974), .Z(n_10815)
		);
	notech_mux2 i_2522453(.S(n_55411), .A(wrD[24]), .B(iwrite_data[24]), .Z(n_57467
		));
	notech_reg tab11_reg_32(.CP(n_63001), .D(n_10821), .CD(n_62267), .Q(\tab11[32] 
		));
	notech_mux2 i_12564(.S(n_56092), .A(\tab11[32] ), .B(n_975), .Z(n_10821)
		);
	notech_mux2 i_2622454(.S(n_55411), .A(wrD[25]), .B(iwrite_data[25]), .Z(n_57474
		));
	notech_reg_set tab11_reg_33(.CP(n_63001), .D(n_10827), .SD(n_62267), .Q(\tab11[33] 
		));
	notech_mux2 i_12572(.S(n_56092), .A(\tab11[33] ), .B(n_56153), .Z(n_10827
		));
	notech_mux2 i_2722455(.S(n_55416), .A(wrD[26]), .B(iwrite_data[26]), .Z(n_57481
		));
	notech_reg fsm5_cnt_reg_0(.CP(n_63001), .D(n_10833), .CD(n_62267), .Q(fsm5_cnt
		[0]));
	notech_mux2 i_12580(.S(\nbus_14505[0] ), .A(fsm5_cnt[0]), .B(n_962), .Z(n_10833
		));
	notech_mux2 i_2822456(.S(n_55411), .A(wrD[27]), .B(iwrite_data[27]), .Z(n_57488
		));
	notech_reg fsm5_cnt_reg_1(.CP(n_63001), .D(n_10839), .CD(n_62267), .Q(fsm5_cnt
		[1]));
	notech_mux2 i_12588(.S(\nbus_14505[0] ), .A(fsm5_cnt[1]), .B(n_963), .Z(n_10839
		));
	notech_mux2 i_2922457(.S(n_55411), .A(wrD[28]), .B(iwrite_data[28]), .Z(n_57495
		));
	notech_reg fsm5_cnt_reg_2(.CP(n_63004), .D(n_10845), .CD(n_62270), .Q(fsm5_cnt
		[2]));
	notech_mux2 i_12596(.S(\nbus_14505[0] ), .A(fsm5_cnt[2]), .B(n_964), .Z(n_10845
		));
	notech_mux2 i_3022458(.S(n_55411), .A(wrD[29]), .B(iwrite_data[29]), .Z(n_57502
		));
	notech_reg fsm5_cnt_reg_3(.CP(n_63004), .D(n_10851), .CD(n_62270), .Q(fsm5_cnt
		[3]));
	notech_mux2 i_12604(.S(\nbus_14505[0] ), .A(fsm5_cnt[3]), .B(n_965), .Z(n_10851
		));
	notech_mux2 i_3122459(.S(n_55411), .A(wrD[30]), .B(iwrite_data[30]), .Z(n_57509
		));
	notech_reg fsm5_cnt_reg_4(.CP(n_63004), .D(n_10857), .CD(n_62270), .Q(fsm5_cnt
		[4]));
	notech_mux2 i_12612(.S(\nbus_14505[0] ), .A(fsm5_cnt[4]), .B(n_966), .Z(n_10857
		));
	notech_mux2 i_3222460(.S(n_55411), .A(wrD[31]), .B(iwrite_data[31]), .Z(n_57516
		));
	notech_reg fsm5_cnt_reg_5(.CP(n_63004), .D(n_10863), .CD(n_62270), .Q(fsm5_cnt
		[5]));
	notech_mux2 i_12620(.S(\nbus_14505[0] ), .A(fsm5_cnt[5]), .B(n_967), .Z(n_10863
		));
	notech_nand2 i_8(.A(n_996), .B(n_989), .Z(n_56896));
	notech_reg fsm5_cnt_reg_6(.CP(n_63004), .D(n_10869), .CD(n_62270), .Q(fsm5_cnt
		[6]));
	notech_mux2 i_12628(.S(\nbus_14505[0] ), .A(fsm5_cnt[6]), .B(n_968), .Z(n_10869
		));
	notech_or2 i_79240(.A(n_974), .B(data_miss[6]), .Z(n_56902));
	notech_reg fsm5_cnt_reg_7(.CP(n_63001), .D(n_10875), .CD(n_62267), .Q(fsm5_cnt
		[7]));
	notech_mux2 i_12636(.S(\nbus_14505[0] ), .A(fsm5_cnt[7]), .B(n_969), .Z(n_10875
		));
	notech_nand2 i_122397(.A(n_1287), .B(n_475), .Z(n_57966));
	notech_reg fsm5_cnt_reg_8(.CP(n_63001), .D(n_10881), .CD(n_62267), .Q(fsm5_cnt
		[8]));
	notech_mux2 i_12644(.S(\nbus_14505[0] ), .A(fsm5_cnt[8]), .B(n_970), .Z(n_10881
		));
	notech_nand2 i_222398(.A(n_1286), .B(n_476), .Z(n_57973));
	notech_reg pg_fault_reg(.CP(n_63004), .D(n_10887), .CD(n_62270), .Q(pg_fault
		));
	notech_mux2 i_12652(.S(n_56850), .A(pg_fault), .B(n_11996), .Z(n_10887)
		);
	notech_nand2 i_322399(.A(n_1285), .B(n_477), .Z(n_57980));
	notech_reg fsm_reg_0(.CP(n_63001), .D(n_10893), .CD(n_62267), .Q(fsm[0])
		);
	notech_mux2 i_12660(.S(\nbus_14509[0] ), .A(fsm[0]), .B(n_58606), .Z(n_10893
		));
	notech_nand2 i_422400(.A(n_1284), .B(n_478), .Z(n_57987));
	notech_reg fsm_reg_1(.CP(n_63000), .D(n_10899), .CD(n_62266), .Q(fsm[1])
		);
	notech_mux2 i_12668(.S(\nbus_14509[0] ), .A(fsm[1]), .B(n_11997), .Z(n_10899
		));
	notech_nand2 i_522401(.A(n_1283), .B(n_479), .Z(n_57994));
	notech_reg fsm_reg_2(.CP(n_63000), .D(n_10905), .CD(n_62266), .Q(fsm[2])
		);
	notech_mux2 i_12676(.S(\nbus_14509[0] ), .A(fsm[2]), .B(n_11999), .Z(n_10905
		));
	notech_nand2 i_622402(.A(n_1282), .B(n_480), .Z(n_58001));
	notech_reg fsm_reg_3(.CP(n_63000), .D(n_10911), .CD(n_62266), .Q(fsm[3])
		);
	notech_mux2 i_12684(.S(\nbus_14509[0] ), .A(fsm[3]), .B(n_961), .Z(n_10911
		));
	notech_nand2 i_722403(.A(n_1281), .B(n_481), .Z(n_58008));
	notech_reg owrite_req_reg(.CP(n_63000), .D(n_60392), .CD(n_62266), .Q(owrite_req
		));
	notech_reg pt_fault_reg(.CP(n_63000), .D(n_10919), .CD(n_62266), .Q(pt_fault
		));
	notech_mux2 i_12696(.S(n_945), .A(data_miss[0]), .B(pt_fault), .Z(n_10919
		));
	notech_nand2 i_822404(.A(n_1280), .B(n_482), .Z(n_58015));
	notech_reg addr_miss_reg_0(.CP(n_63000), .D(n_10928), .CD(n_62266), .Q(addr_miss
		[0]));
	notech_and3 i_12706(.A(n_1020), .B(n_545), .C(addr_miss[0]), .Z(n_10928)
		);
	notech_nand2 i_922405(.A(n_1279), .B(n_483), .Z(n_58022));
	notech_reg addr_miss_reg_1(.CP(n_63000), .D(n_10934), .CD(n_62266), .Q(addr_miss
		[1]));
	notech_and3 i_12714(.A(n_1020), .B(n_545), .C(addr_miss[1]), .Z(n_10934)
		);
	notech_nand2 i_1022406(.A(n_1278), .B(n_484), .Z(n_58029));
	notech_reg addr_miss_reg_2(.CP(n_63000), .D(n_10937), .CD(n_62266), .Q(addr_miss
		[2]));
	notech_mux2 i_12720(.S(\nbus_14514[0] ), .A(addr_miss[2]), .B(n_12002), 
		.Z(n_10937));
	notech_nand2 i_1122407(.A(n_1277), .B(n_485), .Z(n_58036));
	notech_reg addr_miss_reg_3(.CP(n_63000), .D(n_10943), .CD(n_62266), .Q(addr_miss
		[3]));
	notech_mux2 i_12728(.S(\nbus_14514[0] ), .A(addr_miss[3]), .B(n_12003), 
		.Z(n_10943));
	notech_nand2 i_1222408(.A(n_1276), .B(n_487), .Z(n_58043));
	notech_reg addr_miss_reg_4(.CP(n_63001), .D(n_10949), .CD(n_62267), .Q(addr_miss
		[4]));
	notech_mux2 i_12736(.S(\nbus_14514[0] ), .A(addr_miss[4]), .B(n_12004), 
		.Z(n_10949));
	notech_and4 i_1322409(.A(n_1272), .B(n_1274), .C(n_1271), .D(n_685), .Z(n_58050
		));
	notech_reg addr_miss_reg_5(.CP(n_63001), .D(n_10955), .CD(n_62267), .Q(addr_miss
		[5]));
	notech_mux2 i_12744(.S(\nbus_14514[0] ), .A(addr_miss[5]), .B(n_12005), 
		.Z(n_10955));
	notech_and4 i_1422410(.A(n_1263), .B(n_1265), .C(n_1262), .D(n_696), .Z(n_58057
		));
	notech_reg addr_miss_reg_6(.CP(n_63001), .D(n_10961), .CD(n_62267), .Q(addr_miss
		[6]));
	notech_mux2 i_12752(.S(\nbus_14514[0] ), .A(addr_miss[6]), .B(n_12006), 
		.Z(n_10961));
	notech_and4 i_1522411(.A(n_1254), .B(n_1256), .C(n_1253), .D(n_707), .Z(n_58064
		));
	notech_reg addr_miss_reg_7(.CP(n_63001), .D(n_10967), .CD(n_62267), .Q(addr_miss
		[7]));
	notech_mux2 i_12760(.S(\nbus_14514[0] ), .A(addr_miss[7]), .B(n_12007), 
		.Z(n_10967));
	notech_and4 i_1622412(.A(n_1245), .B(n_1247), .C(n_1244), .D(n_718), .Z(n_58071
		));
	notech_reg addr_miss_reg_8(.CP(n_63001), .D(n_10973), .CD(n_62267), .Q(addr_miss
		[8]));
	notech_mux2 i_12768(.S(\nbus_14514[0] ), .A(addr_miss[8]), .B(n_12008), 
		.Z(n_10973));
	notech_and4 i_1722413(.A(n_1236), .B(n_1238), .C(n_1235), .D(n_729), .Z(n_58078
		));
	notech_reg addr_miss_reg_9(.CP(n_63001), .D(n_10979), .CD(n_62267), .Q(addr_miss
		[9]));
	notech_mux2 i_12776(.S(\nbus_14514[0] ), .A(addr_miss[9]), .B(n_12009), 
		.Z(n_10979));
	notech_and4 i_1822414(.A(n_1227), .B(n_1229), .C(n_1226), .D(n_740), .Z(n_58085
		));
	notech_reg addr_miss_reg_10(.CP(n_63000), .D(n_10985), .CD(n_62266), .Q(addr_miss
		[10]));
	notech_mux2 i_12784(.S(\nbus_14514[0] ), .A(addr_miss[10]), .B(n_12010),
		 .Z(n_10985));
	notech_and4 i_1922415(.A(n_1218), .B(n_1220), .C(n_1217), .D(n_751), .Z(n_58092
		));
	notech_reg addr_miss_reg_11(.CP(n_63001), .D(n_10991), .CD(n_62267), .Q(addr_miss
		[11]));
	notech_mux2 i_12792(.S(\nbus_14514[0] ), .A(addr_miss[11]), .B(n_12011),
		 .Z(n_10991));
	notech_and4 i_2022416(.A(n_1209), .B(n_1211), .C(n_1208), .D(n_762), .Z(n_58099
		));
	notech_reg addr_miss_reg_12(.CP(n_63001), .D(n_10997), .CD(n_62267), .Q(addr_miss
		[12]));
	notech_mux2 i_12800(.S(\nbus_14514[0] ), .A(addr_miss[12]), .B(n_59578),
		 .Z(n_10997));
	notech_and4 i_2122417(.A(n_1200), .B(n_1202), .C(n_1199), .D(n_773), .Z(n_58106
		));
	notech_reg addr_miss_reg_13(.CP(n_63004), .D(n_11003), .CD(n_62270), .Q(addr_miss
		[13]));
	notech_mux2 i_12808(.S(\nbus_14514[0] ), .A(addr_miss[13]), .B(n_59584),
		 .Z(n_11003));
	notech_and4 i_2222418(.A(n_1191), .B(n_1193), .C(n_1190), .D(n_784), .Z(n_58113
		));
	notech_reg addr_miss_reg_14(.CP(n_63009), .D(n_11009), .CD(n_62275), .Q(addr_miss
		[14]));
	notech_mux2 i_12816(.S(\nbus_14514[0] ), .A(addr_miss[14]), .B(n_59590),
		 .Z(n_11009));
	notech_and4 i_2322419(.A(n_1182), .B(n_1184), .C(n_1181), .D(n_795), .Z(n_58120
		));
	notech_reg addr_miss_reg_15(.CP(n_63006), .D(n_11015), .CD(n_62272), .Q(addr_miss
		[15]));
	notech_mux2 i_12824(.S(\nbus_14514[0] ), .A(addr_miss[15]), .B(n_59596),
		 .Z(n_11015));
	notech_and4 i_2422420(.A(n_1173), .B(n_1175), .C(n_1172), .D(n_806), .Z(n_58127
		));
	notech_reg addr_miss_reg_16(.CP(n_63009), .D(n_11021), .CD(n_62275), .Q(addr_miss
		[16]));
	notech_mux2 i_12832(.S(\nbus_14514[0] ), .A(addr_miss[16]), .B(n_59602),
		 .Z(n_11021));
	notech_and4 i_2522421(.A(n_1164), .B(n_1166), .C(n_1163), .D(n_817), .Z(n_58134
		));
	notech_reg addr_miss_reg_17(.CP(n_63009), .D(n_11027), .CD(n_62275), .Q(addr_miss
		[17]));
	notech_mux2 i_12840(.S(n_56310), .A(addr_miss[17]), .B(n_59608), .Z(n_11027
		));
	notech_and4 i_2622422(.A(n_1155), .B(n_1157), .C(n_1154), .D(n_828), .Z(n_58141
		));
	notech_reg addr_miss_reg_18(.CP(n_63006), .D(n_11033), .CD(n_62272), .Q(addr_miss
		[18]));
	notech_mux2 i_12848(.S(n_56310), .A(addr_miss[18]), .B(n_59614), .Z(n_11033
		));
	notech_and4 i_2722423(.A(n_1146), .B(n_1148), .C(n_1145), .D(n_839), .Z(n_58148
		));
	notech_reg addr_miss_reg_19(.CP(n_63006), .D(n_11039), .CD(n_62272), .Q(addr_miss
		[19]));
	notech_mux2 i_12856(.S(n_56310), .A(addr_miss[19]), .B(n_59620), .Z(n_11039
		));
	notech_and4 i_2822424(.A(n_1137), .B(n_1139), .C(n_1136), .D(n_850), .Z(n_58155
		));
	notech_reg addr_miss_reg_20(.CP(n_63006), .D(n_11045), .CD(n_62272), .Q(addr_miss
		[20]));
	notech_mux2 i_12864(.S(n_56310), .A(addr_miss[20]), .B(n_59626), .Z(n_11045
		));
	notech_and4 i_2922425(.A(n_1128), .B(n_1130), .C(n_1127), .D(n_861), .Z(n_58162
		));
	notech_reg addr_miss_reg_21(.CP(n_63006), .D(n_11051), .CD(n_62272), .Q(addr_miss
		[21]));
	notech_mux2 i_12872(.S(n_56310), .A(addr_miss[21]), .B(n_59632), .Z(n_11051
		));
	notech_and4 i_3022426(.A(n_1119), .B(n_1121), .C(n_1118), .D(n_872), .Z(n_58169
		));
	notech_reg addr_miss_reg_22(.CP(n_63006), .D(n_11057), .CD(n_62272), .Q(addr_miss
		[22]));
	notech_mux2 i_12880(.S(n_56310), .A(addr_miss[22]), .B(n_59638), .Z(n_11057
		));
	notech_and4 i_3122427(.A(n_1110), .B(n_1112), .C(n_1109), .D(n_883), .Z(n_58176
		));
	notech_reg addr_miss_reg_23(.CP(n_63009), .D(n_11063), .CD(n_62275), .Q(addr_miss
		[23]));
	notech_mux2 i_12888(.S(n_56310), .A(addr_miss[23]), .B(n_59644), .Z(n_11063
		));
	notech_and4 i_3222428(.A(n_1101), .B(n_1103), .C(n_1095), .D(n_894), .Z(n_58183
		));
	notech_reg addr_miss_reg_24(.CP(n_63009), .D(n_11069), .CD(n_62275), .Q(addr_miss
		[24]));
	notech_mux2 i_12896(.S(n_56310), .A(addr_miss[24]), .B(n_59650), .Z(n_11069
		));
	notech_nand3 i_79189(.A(n_904), .B(n_903), .C(n_491), .Z(n_58584));
	notech_reg addr_miss_reg_25(.CP(n_63010), .D(n_11075), .CD(n_62276), .Q(addr_miss
		[25]));
	notech_mux2 i_12904(.S(n_56310), .A(addr_miss[25]), .B(n_59656), .Z(n_11075
		));
	notech_reg addr_miss_reg_26(.CP(n_63009), .D(n_11081), .CD(n_62275), .Q(addr_miss
		[26]));
	notech_mux2 i_12912(.S(n_56310), .A(addr_miss[26]), .B(n_59662), .Z(n_11081
		));
	notech_ao4 i_79089(.A(n_56290), .B(n_12150), .C(n_1016), .D(n_12160), .Z
		(n_59518));
	notech_reg addr_miss_reg_27(.CP(n_63009), .D(n_11087), .CD(n_62275), .Q(addr_miss
		[27]));
	notech_mux2 i_12920(.S(n_56310), .A(addr_miss[27]), .B(n_59668), .Z(n_11087
		));
	notech_ao4 i_79092(.A(n_56290), .B(n_12149), .C(n_1016), .D(n_12159), .Z
		(n_59524));
	notech_reg addr_miss_reg_28(.CP(n_63009), .D(n_11093), .CD(n_62275), .Q(addr_miss
		[28]));
	notech_mux2 i_12928(.S(n_56310), .A(addr_miss[28]), .B(n_59674), .Z(n_11093
		));
	notech_ao4 i_79095(.A(n_56290), .B(n_12148), .C(n_1016), .D(n_12158), .Z
		(n_59530));
	notech_reg addr_miss_reg_29(.CP(n_63009), .D(n_11099), .CD(n_62275), .Q(addr_miss
		[29]));
	notech_mux2 i_12936(.S(n_56310), .A(addr_miss[29]), .B(n_59680), .Z(n_11099
		));
	notech_ao4 i_79098(.A(n_56290), .B(n_12147), .C(n_1016), .D(n_12157), .Z
		(n_59536));
	notech_reg addr_miss_reg_30(.CP(n_63009), .D(n_11105), .CD(n_62275), .Q(addr_miss
		[30]));
	notech_mux2 i_12944(.S(n_56310), .A(addr_miss[30]), .B(n_59686), .Z(n_11105
		));
	notech_ao4 i_79101(.A(n_56290), .B(n_12146), .C(n_1016), .D(n_12156), .Z
		(n_59542));
	notech_reg addr_miss_reg_31(.CP(n_63009), .D(n_11111), .CD(n_62275), .Q(addr_miss
		[31]));
	notech_mux2 i_12952(.S(n_56310), .A(addr_miss[31]), .B(n_59692), .Z(n_11111
		));
	notech_ao4 i_79104(.A(n_56290), .B(n_12145), .C(n_1016), .D(n_12155), .Z
		(n_59548));
	notech_reg cr2_reg_0(.CP(n_63004), .D(n_11117), .CD(n_62270), .Q(cr2[0])
		);
	notech_mux2 i_12960(.S(n_945), .A(iDaddr_f[0]), .B(cr2[0]), .Z(n_11117)
		);
	notech_ao4 i_79107(.A(n_56290), .B(n_12144), .C(n_1016), .D(n_12154), .Z
		(n_59554));
	notech_reg cr2_reg_1(.CP(n_63004), .D(n_11123), .CD(n_62270), .Q(cr2[1])
		);
	notech_mux2 i_12968(.S(n_945), .A(iDaddr_f[1]), .B(cr2[1]), .Z(n_11123)
		);
	notech_ao4 i_79110(.A(n_56290), .B(n_12143), .C(n_1016), .D(n_12153), .Z
		(n_59560));
	notech_reg cr2_reg_2(.CP(n_63004), .D(n_11129), .CD(n_62270), .Q(cr2[2])
		);
	notech_mux2 i_12976(.S(n_945), .A(iDaddr_f[2]), .B(cr2[2]), .Z(n_11129)
		);
	notech_ao4 i_79113(.A(n_56290), .B(n_12142), .C(n_1016), .D(n_12152), .Z
		(n_59566));
	notech_reg cr2_reg_3(.CP(n_63004), .D(n_11135), .CD(n_62270), .Q(cr2[3])
		);
	notech_mux2 i_12984(.S(n_945), .A(iDaddr_f[3]), .B(cr2[3]), .Z(n_11135)
		);
	notech_ao4 i_79116(.A(n_56290), .B(n_12141), .C(n_1016), .D(n_12151), .Z
		(n_59572));
	notech_reg cr2_reg_4(.CP(n_63004), .D(n_11141), .CD(n_62270), .Q(cr2[4])
		);
	notech_mux2 i_12992(.S(n_945), .A(iDaddr_f[4]), .B(cr2[4]), .Z(n_11141)
		);
	notech_nand2 i_79119(.A(n_1076), .B(n_515), .Z(n_59578));
	notech_reg cr2_reg_5(.CP(n_63004), .D(n_11147), .CD(n_62270), .Q(cr2[5])
		);
	notech_mux2 i_13000(.S(n_945), .A(iDaddr_f[5]), .B(cr2[5]), .Z(n_11147)
		);
	notech_nand2 i_79122(.A(n_1075), .B(n_516), .Z(n_59584));
	notech_reg cr2_reg_6(.CP(n_63004), .D(n_11153), .CD(n_62270), .Q(cr2[6])
		);
	notech_mux2 i_13008(.S(n_945), .A(iDaddr_f[6]), .B(cr2[6]), .Z(n_11153)
		);
	notech_nand2 i_79125(.A(n_1074), .B(n_517), .Z(n_59590));
	notech_reg cr2_reg_7(.CP(n_63004), .D(n_11159), .CD(n_62270), .Q(cr2[7])
		);
	notech_mux2 i_13016(.S(n_945), .A(iDaddr_f[7]), .B(cr2[7]), .Z(n_11159)
		);
	notech_nand2 i_79128(.A(n_1073), .B(n_518), .Z(n_59596));
	notech_reg cr2_reg_8(.CP(n_63004), .D(n_11165), .CD(n_62270), .Q(cr2[8])
		);
	notech_mux2 i_13024(.S(n_945), .A(iDaddr_f[8]), .B(cr2[8]), .Z(n_11165)
		);
	notech_nand2 i_79131(.A(n_1072), .B(n_519), .Z(n_59602));
	notech_reg cr2_reg_9(.CP(n_63006), .D(n_11171), .CD(n_62272), .Q(cr2[9])
		);
	notech_mux2 i_13032(.S(n_945), .A(iDaddr_f[9]), .B(cr2[9]), .Z(n_11171)
		);
	notech_nand2 i_79134(.A(n_1071), .B(n_520), .Z(n_59608));
	notech_reg cr2_reg_10(.CP(n_63006), .D(n_11177), .CD(n_62272), .Q(cr2[10
		]));
	notech_mux2 i_13040(.S(n_945), .A(iDaddr_f[10]), .B(cr2[10]), .Z(n_11177
		));
	notech_nand2 i_79137(.A(n_1070), .B(n_521), .Z(n_59614));
	notech_reg cr2_reg_11(.CP(n_63006), .D(n_11183), .CD(n_62272), .Q(cr2[11
		]));
	notech_mux2 i_13048(.S(n_945), .A(iDaddr_f[11]), .B(cr2[11]), .Z(n_11183
		));
	notech_nand2 i_79140(.A(n_1069), .B(n_522), .Z(n_59620));
	notech_reg cr2_reg_12(.CP(n_63006), .D(n_11189), .CD(n_62272), .Q(cr2[12
		]));
	notech_mux2 i_13056(.S(n_945), .A(iDaddr_f[12]), .B(cr2[12]), .Z(n_11189
		));
	notech_nand2 i_79143(.A(n_1068), .B(n_523), .Z(n_59626));
	notech_reg cr2_reg_13(.CP(n_63006), .D(n_11195), .CD(n_62272), .Q(cr2[13
		]));
	notech_mux2 i_13064(.S(n_945), .A(iDaddr_f[13]), .B(cr2[13]), .Z(n_11195
		));
	notech_nand2 i_79146(.A(n_1067), .B(n_524), .Z(n_59632));
	notech_reg cr2_reg_14(.CP(n_63004), .D(n_11201), .CD(n_62270), .Q(cr2[14
		]));
	notech_mux2 i_13072(.S(n_945), .A(iDaddr_f[14]), .B(cr2[14]), .Z(n_11201
		));
	notech_nand2 i_79149(.A(n_1066), .B(n_525), .Z(n_59638));
	notech_reg cr2_reg_15(.CP(n_63004), .D(n_11207), .CD(n_62270), .Q(cr2[15
		]));
	notech_mux2 i_13080(.S(n_945), .A(iDaddr_f[15]), .B(cr2[15]), .Z(n_11207
		));
	notech_nand2 i_79152(.A(n_1065), .B(n_526), .Z(n_59644));
	notech_reg cr2_reg_16(.CP(n_63004), .D(n_11213), .CD(n_62270), .Q(cr2[16
		]));
	notech_mux2 i_13088(.S(n_55559), .A(iDaddr_f[16]), .B(cr2[16]), .Z(n_11213
		));
	notech_nand2 i_79155(.A(n_1064), .B(n_527), .Z(n_59650));
	notech_reg cr2_reg_17(.CP(n_63004), .D(n_11219), .CD(n_62270), .Q(cr2[17
		]));
	notech_mux2 i_13096(.S(n_55559), .A(iDaddr_f[17]), .B(cr2[17]), .Z(n_11219
		));
	notech_nand2 i_79158(.A(n_1063), .B(n_528), .Z(n_59656));
	notech_reg cr2_reg_18(.CP(n_63033), .D(n_11225), .CD(n_62299), .Q(cr2[18
		]));
	notech_mux2 i_13104(.S(n_55559), .A(iDaddr_f[18]), .B(cr2[18]), .Z(n_11225
		));
	notech_nand2 i_79161(.A(n_1062), .B(n_529), .Z(n_59662));
	notech_reg cr2_reg_19(.CP(n_63033), .D(n_11231), .CD(n_62299), .Q(cr2[19
		]));
	notech_mux2 i_13112(.S(n_55559), .A(iDaddr_f[19]), .B(cr2[19]), .Z(n_11231
		));
	notech_nand2 i_79164(.A(n_1061), .B(n_530), .Z(n_59668));
	notech_reg cr2_reg_20(.CP(n_63033), .D(n_11237), .CD(n_62299), .Q(cr2[20
		]));
	notech_mux2 i_13120(.S(n_55559), .A(iDaddr_f[20]), .B(cr2[20]), .Z(n_11237
		));
	notech_nand2 i_79167(.A(n_1060), .B(n_531), .Z(n_59674));
	notech_reg cr2_reg_21(.CP(n_63033), .D(n_11243), .CD(n_62299), .Q(cr2[21
		]));
	notech_mux2 i_13128(.S(n_55559), .A(iDaddr_f[21]), .B(cr2[21]), .Z(n_11243
		));
	notech_nand2 i_79170(.A(n_1059), .B(n_532), .Z(n_59680));
	notech_reg cr2_reg_22(.CP(n_63033), .D(n_11249), .CD(n_62299), .Q(cr2[22
		]));
	notech_mux2 i_13136(.S(n_55559), .A(iDaddr_f[22]), .B(cr2[22]), .Z(n_11249
		));
	notech_nand2 i_79173(.A(n_1058), .B(n_533), .Z(n_59686));
	notech_reg cr2_reg_23(.CP(n_63033), .D(n_11255), .CD(n_62299), .Q(cr2[23
		]));
	notech_mux2 i_13144(.S(n_55559), .A(iDaddr_f[23]), .B(cr2[23]), .Z(n_11255
		));
	notech_nand2 i_79176(.A(n_1057), .B(n_534), .Z(n_59692));
	notech_reg cr2_reg_24(.CP(n_63033), .D(n_11261), .CD(n_62299), .Q(cr2[24
		]));
	notech_mux2 i_13152(.S(n_55559), .A(iDaddr_f[24]), .B(cr2[24]), .Z(n_11261
		));
	notech_mux2 i_79080(.S(iwrite_ack), .A(n_538), .B(n_11871), .Z(n_60392)
		);
	notech_reg cr2_reg_25(.CP(n_63033), .D(n_11267), .CD(n_62299), .Q(cr2[25
		]));
	notech_mux2 i_13160(.S(n_55559), .A(iDaddr_f[25]), .B(cr2[25]), .Z(n_11267
		));
	notech_or4 i_41(.A(n_951), .B(n_1035), .C(n_11895), .D(n_11840), .Z(n_58606
		));
	notech_reg cr2_reg_26(.CP(n_63033), .D(n_11273), .CD(n_62299), .Q(cr2[26
		]));
	notech_mux2 i_13168(.S(n_945), .A(iDaddr_f[26]), .B(cr2[26]), .Z(n_11273
		));
	notech_and4 i_42(.A(n_56290), .B(n_1038), .C(n_990), .D(n_957), .Z(n_58612
		));
	notech_reg cr2_reg_27(.CP(n_63034), .D(n_11279), .CD(n_62300), .Q(cr2[27
		]));
	notech_mux2 i_13176(.S(n_55559), .A(iDaddr_f[27]), .B(cr2[27]), .Z(n_11279
		));
	notech_and4 i_43(.A(n_1016), .B(n_1033), .C(n_549), .D(n_56853), .Z(n_58618
		));
	notech_reg cr2_reg_28(.CP(n_63034), .D(n_11285), .CD(n_62300), .Q(cr2[28
		]));
	notech_mux2 i_13184(.S(n_55559), .A(iDaddr_f[28]), .B(cr2[28]), .Z(n_11285
		));
	notech_or2 i_32(.A(n_56153), .B(\tab11_0[0] ), .Z(n_56627));
	notech_reg cr2_reg_29(.CP(n_63034), .D(n_11291), .CD(n_62300), .Q(cr2[29
		]));
	notech_mux2 i_13192(.S(n_55559), .A(iDaddr_f[29]), .B(cr2[29]), .Z(n_11291
		));
	notech_or2 i_33(.A(n_56153), .B(\tab11_0[1] ), .Z(n_56633));
	notech_reg cr2_reg_30(.CP(n_63034), .D(n_11297), .CD(n_62300), .Q(cr2[30
		]));
	notech_mux2 i_13200(.S(n_55559), .A(iDaddr_f[30]), .B(cr2[30]), .Z(n_11297
		));
	notech_or2 i_34(.A(n_56153), .B(\tab11_0[2] ), .Z(n_56639));
	notech_reg cr2_reg_31(.CP(n_63034), .D(n_11303), .CD(n_62300), .Q(cr2[31
		]));
	notech_mux2 i_13208(.S(n_55559), .A(iDaddr_f[31]), .B(cr2[31]), .Z(n_11303
		));
	notech_or2 i_35(.A(n_56153), .B(\tab11_0[3] ), .Z(n_56645));
	notech_reg req_miss_reg(.CP(n_63034), .D(n_11309), .CD(n_62300), .Q(req_miss
		));
	notech_or2 i_13216(.A(n_11311), .B(n_11312), .Z(n_11309));
	notech_ao4 i_13217(.A(n_11841), .B(n_11842), .C(n_56310), .D(n_11866), .Z
		(n_11311));
	notech_and4 i_13218(.A(req_miss), .B(n_1020), .C(n_545), .D(n_494), .Z(n_11312
		));
	notech_or2 i_36(.A(n_56153), .B(\tab11_0[5] ), .Z(n_56657));
	notech_reg oread_req_reg(.CP(n_63034), .D(n_58584), .CD(n_62300), .Q(oread_req
		));
	notech_reg owrite_sz_reg_0(.CP(n_63034), .D(n_901), .CD(n_62300), .Q(owrite_sz
		[0]));
	notech_reg owrite_sz_reg_1(.CP(n_63034), .D(n_902), .CD(n_62300), .Q(owrite_sz
		[1]));
	notech_reg wrA_reg_0(.CP(n_63032), .D(n_11321), .CD(n_62298), .Q(wrA[0])
		);
	notech_mux2 i_13236(.S(n_55305), .A(wrA[0]), .B(addr_miss[0]), .Z(n_11321
		));
	notech_or2 i_37(.A(n_56153), .B(\tab11_0[6] ), .Z(n_56663));
	notech_reg wrA_reg_1(.CP(n_63032), .D(n_11327), .CD(n_62298), .Q(wrA[1])
		);
	notech_mux2 i_13244(.S(n_55305), .A(wrA[1]), .B(addr_miss[1]), .Z(n_11327
		));
	notech_or2 i_38(.A(n_56153), .B(\tab11_0[7] ), .Z(n_56669));
	notech_reg wrA_reg_2(.CP(n_63032), .D(n_11333), .CD(n_62298), .Q(wrA[2])
		);
	notech_mux2 i_13252(.S(n_55305), .A(wrA[2]), .B(addr_miss[2]), .Z(n_11333
		));
	notech_or2 i_39(.A(n_56153), .B(\tab11_0[8] ), .Z(n_56675));
	notech_reg wrA_reg_3(.CP(n_63032), .D(n_11339), .CD(n_62298), .Q(wrA[3])
		);
	notech_mux2 i_13260(.S(n_55305), .A(wrA[3]), .B(addr_miss[3]), .Z(n_11339
		));
	notech_or2 i_40(.A(n_56153), .B(\tab11_0[9] ), .Z(n_56681));
	notech_reg wrA_reg_4(.CP(n_63030), .D(n_11345), .CD(n_62296), .Q(wrA[4])
		);
	notech_mux2 i_13268(.S(n_55305), .A(wrA[4]), .B(addr_miss[4]), .Z(n_11345
		));
	notech_or2 i_45(.A(data_miss[12]), .B(n_56153), .Z(n_56687));
	notech_reg wrA_reg_5(.CP(n_63030), .D(n_11351), .CD(n_62296), .Q(wrA[5])
		);
	notech_mux2 i_13276(.S(n_55305), .A(wrA[5]), .B(addr_miss[5]), .Z(n_11351
		));
	notech_or2 i_47(.A(data_miss[13]), .B(n_56153), .Z(n_56693));
	notech_reg wrA_reg_6(.CP(n_63030), .D(n_11357), .CD(n_62296), .Q(wrA[6])
		);
	notech_mux2 i_13284(.S(n_55305), .A(wrA[6]), .B(addr_miss[6]), .Z(n_11357
		));
	notech_or2 i_48(.A(data_miss[14]), .B(n_56148), .Z(n_56699));
	notech_reg wrA_reg_7(.CP(n_63030), .D(n_11363), .CD(n_62296), .Q(wrA[7])
		);
	notech_mux2 i_13292(.S(n_55305), .A(wrA[7]), .B(addr_miss[7]), .Z(n_11363
		));
	notech_or2 i_49(.A(data_miss[15]), .B(n_56148), .Z(n_56705));
	notech_reg wrA_reg_8(.CP(n_63030), .D(n_11369), .CD(n_62296), .Q(wrA[8])
		);
	notech_mux2 i_13300(.S(n_55305), .A(wrA[8]), .B(addr_miss[8]), .Z(n_11369
		));
	notech_or2 i_51(.A(data_miss[16]), .B(n_56148), .Z(n_56711));
	notech_reg wrA_reg_9(.CP(n_63032), .D(n_11375), .CD(n_62298), .Q(wrA[9])
		);
	notech_mux2 i_13308(.S(n_55305), .A(wrA[9]), .B(addr_miss[9]), .Z(n_11375
		));
	notech_or2 i_52(.A(data_miss[17]), .B(n_56148), .Z(n_56717));
	notech_reg wrA_reg_10(.CP(n_63032), .D(n_11381), .CD(n_62298), .Q(wrA[10
		]));
	notech_mux2 i_13316(.S(n_55305), .A(wrA[10]), .B(addr_miss[10]), .Z(n_11381
		));
	notech_or2 i_53(.A(data_miss[18]), .B(n_56148), .Z(n_56723));
	notech_reg wrA_reg_11(.CP(n_63033), .D(n_11387), .CD(n_62299), .Q(wrA[11
		]));
	notech_mux2 i_13324(.S(n_55305), .A(wrA[11]), .B(addr_miss[11]), .Z(n_11387
		));
	notech_or2 i_54(.A(data_miss[19]), .B(n_56148), .Z(n_56729));
	notech_reg wrA_reg_12(.CP(n_63033), .D(n_11393), .CD(n_62299), .Q(wrA[12
		]));
	notech_mux2 i_13332(.S(n_55305), .A(wrA[12]), .B(addr_miss[12]), .Z(n_11393
		));
	notech_or2 i_55(.A(data_miss[20]), .B(n_56148), .Z(n_56735));
	notech_reg wrA_reg_13(.CP(n_63032), .D(n_11399), .CD(n_62298), .Q(wrA[13
		]));
	notech_mux2 i_13340(.S(n_55305), .A(wrA[13]), .B(addr_miss[13]), .Z(n_11399
		));
	notech_or2 i_56(.A(data_miss[21]), .B(n_56148), .Z(n_56741));
	notech_reg wrA_reg_14(.CP(n_63032), .D(n_11405), .CD(n_62298), .Q(wrA[14
		]));
	notech_mux2 i_13348(.S(n_55305), .A(wrA[14]), .B(addr_miss[14]), .Z(n_11405
		));
	notech_or2 i_57(.A(data_miss[22]), .B(n_56148), .Z(n_56747));
	notech_reg wrA_reg_15(.CP(n_63032), .D(n_11411), .CD(n_62298), .Q(wrA[15
		]));
	notech_mux2 i_13356(.S(n_55305), .A(wrA[15]), .B(addr_miss[15]), .Z(n_11411
		));
	notech_or2 i_58(.A(data_miss[23]), .B(n_56148), .Z(n_56753));
	notech_reg wrA_reg_16(.CP(n_63032), .D(n_11417), .CD(n_62298), .Q(wrA[16
		]));
	notech_mux2 i_13364(.S(n_55307), .A(wrA[16]), .B(addr_miss[16]), .Z(n_11417
		));
	notech_or2 i_59(.A(data_miss[24]), .B(n_56148), .Z(n_56759));
	notech_reg wrA_reg_17(.CP(n_63032), .D(n_11423), .CD(n_62298), .Q(wrA[17
		]));
	notech_mux2 i_13372(.S(n_55307), .A(wrA[17]), .B(addr_miss[17]), .Z(n_11423
		));
	notech_or2 i_60(.A(data_miss[25]), .B(n_56153), .Z(n_56765));
	notech_reg wrA_reg_18(.CP(n_63034), .D(n_11429), .CD(n_62300), .Q(wrA[18
		]));
	notech_mux2 i_13380(.S(n_55307), .A(wrA[18]), .B(addr_miss[18]), .Z(n_11429
		));
	notech_or2 i_61(.A(data_miss[26]), .B(n_56148), .Z(n_56771));
	notech_reg wrA_reg_19(.CP(n_63039), .D(n_11435), .CD(n_62305), .Q(wrA[19
		]));
	notech_mux2 i_13388(.S(n_55307), .A(wrA[19]), .B(addr_miss[19]), .Z(n_11435
		));
	notech_or2 i_62(.A(data_miss[27]), .B(n_56148), .Z(n_56777));
	notech_reg wrA_reg_20(.CP(n_63039), .D(n_11441), .CD(n_62305), .Q(wrA[20
		]));
	notech_mux2 i_13396(.S(n_55307), .A(wrA[20]), .B(addr_miss[20]), .Z(n_11441
		));
	notech_or2 i_63(.A(data_miss[28]), .B(n_56148), .Z(n_56783));
	notech_reg wrA_reg_21(.CP(n_63039), .D(n_11447), .CD(n_62305), .Q(wrA[21
		]));
	notech_mux2 i_13404(.S(n_55307), .A(wrA[21]), .B(addr_miss[21]), .Z(n_11447
		));
	notech_or2 i_64(.A(data_miss[29]), .B(n_56148), .Z(n_56789));
	notech_reg wrA_reg_22(.CP(n_63039), .D(n_11453), .CD(n_62305), .Q(wrA[22
		]));
	notech_mux2 i_13412(.S(n_55307), .A(wrA[22]), .B(addr_miss[22]), .Z(n_11453
		));
	notech_or2 i_65(.A(data_miss[30]), .B(n_56148), .Z(n_56795));
	notech_reg wrA_reg_23(.CP(n_63038), .D(n_11459), .CD(n_62304), .Q(wrA[23
		]));
	notech_mux2 i_13420(.S(n_55307), .A(wrA[23]), .B(addr_miss[23]), .Z(n_11459
		));
	notech_or2 i_66(.A(data_miss[31]), .B(n_56148), .Z(n_56801));
	notech_reg wrA_reg_24(.CP(n_63038), .D(n_11465), .CD(n_62304), .Q(wrA[24
		]));
	notech_mux2 i_13428(.S(n_55307), .A(wrA[24]), .B(addr_miss[24]), .Z(n_11465
		));
	notech_nand2 i_031231(.A(n_989), .B(n_58743), .Z(n_56825));
	notech_reg wrA_reg_25(.CP(n_63038), .D(n_11471), .CD(n_62304), .Q(wrA[25
		]));
	notech_mux2 i_13436(.S(n_55307), .A(wrA[25]), .B(addr_miss[25]), .Z(n_11471
		));
	notech_ao4 i_79836(.A(n_996), .B(n_11988), .C(n_559), .D(n_1026), .Z(n_59705
		));
	notech_reg wrA_reg_26(.CP(n_63038), .D(n_11477), .CD(n_62304), .Q(wrA[26
		]));
	notech_mux2 i_13444(.S(n_55307), .A(wrA[26]), .B(addr_miss[26]), .Z(n_11477
		));
	notech_ao4 i_79839(.A(n_996), .B(n_11990), .C(n_564), .D(n_1026), .Z(n_59711
		));
	notech_reg wrA_reg_27(.CP(n_63038), .D(n_11483), .CD(n_62304), .Q(wrA[27
		]));
	notech_mux2 i_13452(.S(n_55307), .A(wrA[27]), .B(addr_miss[27]), .Z(n_11483
		));
	notech_ao4 i_79826(.A(n_1016), .B(n_11993), .C(n_996), .D(\nnx_tab2[0] )
		, .Z(n_58317));
	notech_reg wrA_reg_28(.CP(n_63039), .D(n_11489), .CD(n_62305), .Q(wrA[28
		]));
	notech_mux2 i_13460(.S(n_55307), .A(wrA[28]), .B(addr_miss[28]), .Z(n_11489
		));
	notech_ao4 i_79829(.A(n_1016), .B(n_11995), .C(n_996), .D(n_573), .Z(n_58323
		));
	notech_reg wrA_reg_29(.CP(n_63039), .D(n_11495), .CD(n_62305), .Q(wrA[29
		]));
	notech_mux2 i_13468(.S(n_55307), .A(wrA[29]), .B(addr_miss[29]), .Z(n_11495
		));
	notech_ao4 i_79607(.A(n_1016), .B(n_11918), .C(n_996), .D(\nnx_tab1[0] )
		, .Z(n_58352));
	notech_reg wrA_reg_30(.CP(n_63041), .D(n_11501), .CD(n_62307), .Q(wrA[30
		]));
	notech_mux2 i_13476(.S(n_55307), .A(wrA[30]), .B(addr_miss[30]), .Z(n_11501
		));
	notech_ao4 i_79610(.A(n_1016), .B(n_11920), .C(n_996), .D(n_585), .Z(n_58358
		));
	notech_reg wrA_reg_31(.CP(n_63041), .D(n_11507), .CD(n_62307), .Q(wrA[31
		]));
	notech_mux2 i_13484(.S(n_55307), .A(wrA[31]), .B(addr_miss[31]), .Z(n_11507
		));
	notech_ao4 i_79856(.A(n_996), .B(n_11922), .C(n_590), .D(n_1017), .Z(n_59073
		));
	notech_reg addr_phys_reg_0(.CP(n_63039), .D(n_57966), .CD(n_62305), .Q(addr_phys
		[0]));
	notech_reg addr_phys_reg_1(.CP(n_63039), .D(n_57973), .CD(n_62305), .Q(addr_phys
		[1]));
	notech_reg addr_phys_reg_2(.CP(n_63039), .D(n_57980), .CD(n_62305), .Q(addr_phys
		[2]));
	notech_reg addr_phys_reg_3(.CP(n_63039), .D(n_57987), .CD(n_62305), .Q(addr_phys
		[3]));
	notech_reg addr_phys_reg_4(.CP(n_63039), .D(n_57994), .CD(n_62305), .Q(addr_phys
		[4]));
	notech_reg addr_phys_reg_5(.CP(n_63037), .D(n_58001), .CD(n_62303), .Q(addr_phys
		[5]));
	notech_reg addr_phys_reg_6(.CP(n_63037), .D(n_58008), .CD(n_62303), .Q(addr_phys
		[6]));
	notech_reg addr_phys_reg_7(.CP(n_63037), .D(n_58015), .CD(n_62303), .Q(addr_phys
		[7]));
	notech_reg addr_phys_reg_8(.CP(n_63037), .D(n_58022), .CD(n_62303), .Q(addr_phys
		[8]));
	notech_reg addr_phys_reg_9(.CP(n_63037), .D(n_58029), .CD(n_62303), .Q(addr_phys
		[9]));
	notech_reg addr_phys_reg_10(.CP(n_63037), .D(n_58036), .CD(n_62303), .Q(addr_phys
		[10]));
	notech_reg addr_phys_reg_11(.CP(n_63034), .D(n_58043), .CD(n_62300), .Q(addr_phys
		[11]));
	notech_reg addr_phys_reg_12(.CP(n_63037), .D(n_12065), .CD(n_62303), .Q(addr_phys
		[12]));
	notech_reg addr_phys_reg_13(.CP(n_63037), .D(n_12066), .CD(n_62303), .Q(addr_phys
		[13]));
	notech_reg addr_phys_reg_14(.CP(n_63038), .D(n_12067), .CD(n_62304), .Q(addr_phys
		[14]));
	notech_reg addr_phys_reg_15(.CP(n_63038), .D(n_12068), .CD(n_62304), .Q(addr_phys
		[15]));
	notech_reg addr_phys_reg_16(.CP(n_63038), .D(n_12069), .CD(n_62304), .Q(addr_phys
		[16]));
	notech_reg addr_phys_reg_17(.CP(n_63038), .D(n_12070), .CD(n_62304), .Q(addr_phys
		[17]));
	notech_reg addr_phys_reg_18(.CP(n_63038), .D(n_12071), .CD(n_62304), .Q(addr_phys
		[18]));
	notech_reg addr_phys_reg_19(.CP(n_63037), .D(n_12072), .CD(n_62303), .Q(addr_phys
		[19]));
	notech_reg addr_phys_reg_20(.CP(n_63037), .D(n_12073), .CD(n_62303), .Q(addr_phys
		[20]));
	notech_reg addr_phys_reg_21(.CP(n_63038), .D(n_12074), .CD(n_62304), .Q(addr_phys
		[21]));
	notech_reg addr_phys_reg_22(.CP(n_63037), .D(n_12075), .CD(n_62303), .Q(addr_phys
		[22]));
	notech_reg addr_phys_reg_23(.CP(n_63030), .D(n_12076), .CD(n_62296), .Q(addr_phys
		[23]));
	notech_reg addr_phys_reg_24(.CP(n_63023), .D(n_12077), .CD(n_62289), .Q(addr_phys
		[24]));
	notech_reg addr_phys_reg_25(.CP(n_63022), .D(n_12078), .CD(n_62288), .Q(addr_phys
		[25]));
	notech_reg addr_phys_reg_26(.CP(n_63023), .D(n_12079), .CD(n_62289), .Q(addr_phys
		[26]));
	notech_reg addr_phys_reg_27(.CP(n_63023), .D(n_12080), .CD(n_62289), .Q(addr_phys
		[27]));
	notech_reg addr_phys_reg_28(.CP(n_63022), .D(n_12081), .CD(n_62288), .Q(addr_phys
		[28]));
	notech_reg addr_phys_reg_29(.CP(n_63022), .D(n_12082), .CD(n_62288), .Q(addr_phys
		[29]));
	notech_reg addr_phys_reg_30(.CP(n_63022), .D(n_12083), .CD(n_62288), .Q(addr_phys
		[30]));
	notech_reg addr_phys_reg_31(.CP(n_63022), .D(n_12084), .CD(n_62288), .Q(addr_phys
		[31]));
	notech_reg wrD_reg_0(.CP(n_63022), .D(n_11577), .CD(n_62288), .Q(wrD[0])
		);
	notech_or2 i_13620(.A(wrD[0]), .B(n_55300), .Z(n_11577));
	notech_ao4 i_79859(.A(n_996), .B(n_11924), .C(n_595), .D(n_1017), .Z(n_59079
		));
	notech_reg wrD_reg_1(.CP(n_63023), .D(n_11583), .CD(n_62289), .Q(wrD[1])
		);
	notech_mux2 i_13628(.S(n_55300), .A(wrD[1]), .B(data_miss[1]), .Z(n_11583
		));
	notech_nand2 i_99(.A(n_59950), .B(n_12150), .Z(n_59751));
	notech_reg wrD_reg_2(.CP(n_63023), .D(n_11589), .CD(n_62289), .Q(wrD[2])
		);
	notech_mux2 i_13636(.S(n_55300), .A(wrD[2]), .B(data_miss[2]), .Z(n_11589
		));
	notech_nand2 i_100(.A(n_59950), .B(n_12149), .Z(n_59757));
	notech_reg wrD_reg_3(.CP(n_63024), .D(n_11595), .CD(n_62290), .Q(wrD[3])
		);
	notech_mux2 i_13644(.S(n_55300), .A(wrD[3]), .B(data_miss[3]), .Z(n_11595
		));
	notech_nand2 i_101(.A(n_59950), .B(n_12148), .Z(n_59763));
	notech_reg wrD_reg_4(.CP(n_63023), .D(n_11601), .CD(n_62289), .Q(wrD[4])
		);
	notech_mux2 i_13652(.S(n_55300), .A(wrD[4]), .B(data_miss[4]), .Z(n_11601
		));
	notech_nand2 i_102(.A(n_59950), .B(n_12147), .Z(n_59769));
	notech_reg wrD_reg_5(.CP(n_63023), .D(n_11607), .CD(n_62289), .Q(wrD[5])
		);
	notech_mux2 i_13660(.S(n_55300), .A(wrD[5]), .B(n_56896), .Z(n_11607));
	notech_nand2 i_103(.A(n_59950), .B(n_12145), .Z(n_59781));
	notech_reg wrD_reg_6(.CP(n_63023), .D(n_11613), .CD(n_62289), .Q(wrD[6])
		);
	notech_mux2 i_13668(.S(n_55300), .A(wrD[6]), .B(n_56902), .Z(n_11613));
	notech_nand2 i_104(.A(n_59950), .B(n_12144), .Z(n_59787));
	notech_reg wrD_reg_7(.CP(n_63023), .D(n_11619), .CD(n_62289), .Q(wrD[7])
		);
	notech_mux2 i_13676(.S(n_55300), .A(wrD[7]), .B(data_miss[7]), .Z(n_11619
		));
	notech_nand2 i_105(.A(n_59950), .B(n_12143), .Z(n_59793));
	notech_reg wrD_reg_8(.CP(n_63023), .D(n_11625), .CD(n_62289), .Q(wrD[8])
		);
	notech_mux2 i_13684(.S(n_55300), .A(wrD[8]), .B(data_miss[8]), .Z(n_11625
		));
	notech_nand2 i_106(.A(n_59950), .B(n_12142), .Z(n_59799));
	notech_reg wrD_reg_9(.CP(n_63023), .D(n_11631), .CD(n_62289), .Q(wrD[9])
		);
	notech_mux2 i_13692(.S(n_55300), .A(wrD[9]), .B(data_miss[9]), .Z(n_11631
		));
	notech_nand2 i_107(.A(n_59950), .B(n_12141), .Z(n_59805));
	notech_reg wrD_reg_10(.CP(n_63020), .D(n_11637), .CD(n_62286), .Q(wrD[10
		]));
	notech_mux2 i_13700(.S(n_55300), .A(wrD[10]), .B(data_miss[10]), .Z(n_11637
		));
	notech_or2 i_108(.A(data_miss[12]), .B(n_11870), .Z(n_59811));
	notech_reg wrD_reg_11(.CP(n_63020), .D(n_11643), .CD(n_62286), .Q(wrD[11
		]));
	notech_mux2 i_13708(.S(n_55300), .A(wrD[11]), .B(data_miss[11]), .Z(n_11643
		));
	notech_or2 i_109(.A(data_miss[13]), .B(n_11870), .Z(n_59817));
	notech_reg wrD_reg_12(.CP(n_63020), .D(n_11649), .CD(n_62286), .Q(wrD[12
		]));
	notech_mux2 i_13716(.S(n_55300), .A(wrD[12]), .B(data_miss[12]), .Z(n_11649
		));
	notech_or2 i_110(.A(data_miss[14]), .B(n_11870), .Z(n_59823));
	notech_reg wrD_reg_13(.CP(n_63020), .D(n_11655), .CD(n_62286), .Q(wrD[13
		]));
	notech_mux2 i_13724(.S(n_55300), .A(wrD[13]), .B(data_miss[13]), .Z(n_11655
		));
	notech_or2 i_111(.A(data_miss[15]), .B(n_11870), .Z(n_59829));
	notech_reg wrD_reg_14(.CP(n_63020), .D(n_11661), .CD(n_62286), .Q(wrD[14
		]));
	notech_mux2 i_13732(.S(n_55300), .A(wrD[14]), .B(data_miss[14]), .Z(n_11661
		));
	notech_or2 i_112(.A(data_miss[16]), .B(n_11870), .Z(n_59835));
	notech_reg wrD_reg_15(.CP(n_63019), .D(n_11667), .CD(n_62285), .Q(wrD[15
		]));
	notech_mux2 i_13740(.S(n_55300), .A(wrD[15]), .B(data_miss[15]), .Z(n_11667
		));
	notech_or2 i_113(.A(data_miss[17]), .B(n_11870), .Z(n_59841));
	notech_reg wrD_reg_16(.CP(n_63019), .D(n_11673), .CD(n_62285), .Q(wrD[16
		]));
	notech_mux2 i_13748(.S(n_55302), .A(wrD[16]), .B(data_miss[16]), .Z(n_11673
		));
	notech_or2 i_114(.A(data_miss[18]), .B(n_11870), .Z(n_59847));
	notech_reg wrD_reg_17(.CP(n_63020), .D(n_11679), .CD(n_62286), .Q(wrD[17
		]));
	notech_mux2 i_13756(.S(n_55302), .A(wrD[17]), .B(data_miss[17]), .Z(n_11679
		));
	notech_or2 i_115(.A(data_miss[19]), .B(n_11870), .Z(n_59853));
	notech_reg wrD_reg_18(.CP(n_63020), .D(n_11685), .CD(n_62286), .Q(wrD[18
		]));
	notech_mux2 i_13764(.S(n_55302), .A(wrD[18]), .B(data_miss[18]), .Z(n_11685
		));
	notech_or2 i_116(.A(data_miss[20]), .B(n_11870), .Z(n_59859));
	notech_reg wrD_reg_19(.CP(n_63022), .D(n_11691), .CD(n_62288), .Q(wrD[19
		]));
	notech_mux2 i_13772(.S(n_55302), .A(wrD[19]), .B(data_miss[19]), .Z(n_11691
		));
	notech_or2 i_117(.A(data_miss[21]), .B(n_56168), .Z(n_59865));
	notech_reg wrD_reg_20(.CP(n_63022), .D(n_11697), .CD(n_62288), .Q(wrD[20
		]));
	notech_mux2 i_13780(.S(n_55302), .A(wrD[20]), .B(data_miss[20]), .Z(n_11697
		));
	notech_or2 i_118(.A(data_miss[22]), .B(n_56168), .Z(n_59871));
	notech_reg wrD_reg_21(.CP(n_63022), .D(n_11703), .CD(n_62288), .Q(wrD[21
		]));
	notech_mux2 i_13788(.S(n_55302), .A(wrD[21]), .B(data_miss[21]), .Z(n_11703
		));
	notech_or2 i_119(.A(data_miss[23]), .B(n_56168), .Z(n_59877));
	notech_reg wrD_reg_22(.CP(n_63022), .D(n_11709), .CD(n_62288), .Q(wrD[22
		]));
	notech_mux2 i_13796(.S(n_55302), .A(wrD[22]), .B(data_miss[22]), .Z(n_11709
		));
	notech_or2 i_120(.A(data_miss[24]), .B(n_56168), .Z(n_59883));
	notech_reg wrD_reg_23(.CP(n_63022), .D(n_11715), .CD(n_62288), .Q(wrD[23
		]));
	notech_mux2 i_13804(.S(n_55302), .A(wrD[23]), .B(data_miss[23]), .Z(n_11715
		));
	notech_or2 i_121(.A(data_miss[25]), .B(n_56168), .Z(n_59889));
	notech_reg wrD_reg_24(.CP(n_63020), .D(n_11721), .CD(n_62286), .Q(wrD[24
		]));
	notech_mux2 i_13812(.S(n_55302), .A(wrD[24]), .B(data_miss[24]), .Z(n_11721
		));
	notech_or2 i_122(.A(data_miss[26]), .B(n_56168), .Z(n_59895));
	notech_reg wrD_reg_25(.CP(n_63020), .D(n_11727), .CD(n_62286), .Q(wrD[25
		]));
	notech_mux2 i_13820(.S(n_55302), .A(wrD[25]), .B(data_miss[25]), .Z(n_11727
		));
	notech_or2 i_123(.A(data_miss[27]), .B(n_56168), .Z(n_59901));
	notech_reg wrD_reg_26(.CP(n_63020), .D(n_11733), .CD(n_62286), .Q(wrD[26
		]));
	notech_mux2 i_13828(.S(n_55302), .A(wrD[26]), .B(data_miss[26]), .Z(n_11733
		));
	notech_or2 i_124(.A(data_miss[28]), .B(n_11870), .Z(n_59907));
	notech_reg wrD_reg_27(.CP(n_63020), .D(n_11739), .CD(n_62286), .Q(wrD[27
		]));
	notech_mux2 i_13836(.S(n_55302), .A(wrD[27]), .B(data_miss[27]), .Z(n_11739
		));
	notech_or2 i_125(.A(data_miss[29]), .B(n_56168), .Z(n_59913));
	notech_reg wrD_reg_28(.CP(n_63024), .D(n_11745), .CD(n_62290), .Q(wrD[28
		]));
	notech_mux2 i_13844(.S(n_55302), .A(wrD[28]), .B(data_miss[28]), .Z(n_11745
		));
	notech_or2 i_126(.A(data_miss[30]), .B(n_56168), .Z(n_59919));
	notech_reg wrD_reg_29(.CP(n_63029), .D(n_11751), .CD(n_62295), .Q(wrD[29
		]));
	notech_mux2 i_13852(.S(n_55302), .A(wrD[29]), .B(data_miss[29]), .Z(n_11751
		));
	notech_or2 i_127(.A(data_miss[31]), .B(n_56168), .Z(n_59925));
	notech_reg wrD_reg_30(.CP(n_63029), .D(n_11757), .CD(n_62295), .Q(wrD[30
		]));
	notech_mux2 i_13860(.S(n_55302), .A(wrD[30]), .B(data_miss[30]), .Z(n_11757
		));
	notech_ao4 i_3(.A(data_miss[0]), .B(n_989), .C(n_984), .D(n_985), .Z(n_59950
		));
	notech_reg wrD_reg_31(.CP(n_63029), .D(n_11763), .CD(n_62295), .Q(wrD[31
		]));
	notech_mux2 i_13868(.S(n_55302), .A(wrD[31]), .B(data_miss[31]), .Z(n_11763
		));
	notech_reg owrite_data_reg_0(.CP(n_63029), .D(n_57299), .CD(n_62295), .Q
		(owrite_data[0]));
	notech_reg owrite_data_reg_1(.CP(n_63029), .D(n_57306), .CD(n_62295), .Q
		(owrite_data[1]));
	notech_reg owrite_data_reg_2(.CP(n_63028), .D(n_57313), .CD(n_62294), .Q
		(owrite_data[2]));
	notech_reg owrite_data_reg_3(.CP(n_63028), .D(n_57320), .CD(n_62294), .Q
		(owrite_data[3]));
	notech_reg owrite_data_reg_4(.CP(n_63029), .D(n_57327), .CD(n_62295), .Q
		(owrite_data[4]));
	notech_reg owrite_data_reg_5(.CP(n_63029), .D(n_57334), .CD(n_62295), .Q
		(owrite_data[5]));
	notech_reg owrite_data_reg_6(.CP(n_63030), .D(n_57341), .CD(n_62296), .Q
		(owrite_data[6]));
	notech_reg owrite_data_reg_7(.CP(n_63030), .D(n_57348), .CD(n_62296), .Q
		(owrite_data[7]));
	notech_reg owrite_data_reg_8(.CP(n_63030), .D(n_57355), .CD(n_62296), .Q
		(owrite_data[8]));
	notech_reg owrite_data_reg_9(.CP(n_63030), .D(n_57362), .CD(n_62296), .Q
		(owrite_data[9]));
	notech_reg owrite_data_reg_10(.CP(n_63030), .D(n_57369), .CD(n_62296), .Q
		(owrite_data[10]));
	notech_reg owrite_data_reg_11(.CP(n_63029), .D(n_57376), .CD(n_62295), .Q
		(owrite_data[11]));
	notech_reg owrite_data_reg_12(.CP(n_63029), .D(n_57383), .CD(n_62295), .Q
		(owrite_data[12]));
	notech_reg owrite_data_reg_13(.CP(n_63029), .D(n_57390), .CD(n_62295), .Q
		(owrite_data[13]));
	notech_reg owrite_data_reg_14(.CP(n_63029), .D(n_57397), .CD(n_62295), .Q
		(owrite_data[14]));
	notech_reg owrite_data_reg_15(.CP(n_63024), .D(n_57404), .CD(n_62290), .Q
		(owrite_data[15]));
	notech_reg owrite_data_reg_16(.CP(n_63024), .D(n_57411), .CD(n_62290), .Q
		(owrite_data[16]));
	notech_reg owrite_data_reg_17(.CP(n_63024), .D(n_57418), .CD(n_62290), .Q
		(owrite_data[17]));
	notech_reg owrite_data_reg_18(.CP(n_63024), .D(n_57425), .CD(n_62290), .Q
		(owrite_data[18]));
	notech_reg owrite_data_reg_19(.CP(n_63024), .D(n_57432), .CD(n_62290), .Q
		(owrite_data[19]));
	notech_reg owrite_data_reg_20(.CP(n_63024), .D(n_57439), .CD(n_62290), .Q
		(owrite_data[20]));
	notech_reg owrite_data_reg_21(.CP(n_63024), .D(n_57446), .CD(n_62290), .Q
		(owrite_data[21]));
	notech_reg owrite_data_reg_22(.CP(n_63024), .D(n_57453), .CD(n_62290), .Q
		(owrite_data[22]));
	notech_reg owrite_data_reg_23(.CP(n_63024), .D(n_57460), .CD(n_62290), .Q
		(owrite_data[23]));
	notech_reg owrite_data_reg_24(.CP(n_63028), .D(n_57467), .CD(n_62294), .Q
		(owrite_data[24]));
	notech_reg owrite_data_reg_25(.CP(n_63028), .D(n_57474), .CD(n_62294), .Q
		(owrite_data[25]));
	notech_reg owrite_data_reg_26(.CP(n_63028), .D(n_57481), .CD(n_62294), .Q
		(owrite_data[26]));
	notech_reg owrite_data_reg_27(.CP(n_63028), .D(n_57488), .CD(n_62294), .Q
		(owrite_data[27]));
	notech_reg owrite_data_reg_28(.CP(n_63028), .D(n_57495), .CD(n_62294), .Q
		(owrite_data[28]));
	notech_reg owrite_data_reg_29(.CP(n_63028), .D(n_57502), .CD(n_62294), .Q
		(owrite_data[29]));
	notech_reg owrite_data_reg_30(.CP(n_63028), .D(n_57509), .CD(n_62294), .Q
		(owrite_data[30]));
	notech_reg owrite_data_reg_31(.CP(n_63028), .D(n_57516), .CD(n_62294), .Q
		(owrite_data[31]));
	notech_reg wr_fault_reg(.CP(n_63028), .D(n_11833), .CD(n_62294), .Q(wr_fault
		));
	notech_mux2 i_14004(.S(n_56836), .A(wr_fault), .B(n_656), .Z(n_11833));
	notech_inv i_15701(.A(n_1050), .Z(n_11840));
	notech_inv i_15702(.A(n_56290), .Z(n_11841));
	notech_inv i_15703(.A(n_1016), .Z(n_11842));
	notech_inv i_15704(.A(n_55411), .Z(n_11843));
	notech_inv i_15705(.A(n_987), .Z(n_11844));
	notech_inv i_15706(.A(n_999), .Z(n_11845));
	notech_inv i_15707(.A(n_1015), .Z(n_11846));
	notech_inv i_15708(.A(n_985), .Z(n_11847));
	notech_inv i_15709(.A(n_983), .Z(n_11848));
	notech_inv i_15710(.A(\dir1[10] ), .Z(n_11849));
	notech_inv i_15711(.A(\dir1[11] ), .Z(n_11850));
	notech_inv i_15712(.A(\dir1[12] ), .Z(n_11851));
	notech_inv i_15713(.A(\dir1[13] ), .Z(n_11852));
	notech_inv i_15714(.A(\dir1[14] ), .Z(n_11853));
	notech_inv i_15715(.A(\dir1[15] ), .Z(n_11854));
	notech_inv i_15716(.A(\dir1[16] ), .Z(n_11855));
	notech_inv i_15717(.A(\dir1[17] ), .Z(n_11856));
	notech_inv i_15718(.A(\dir1[18] ), .Z(n_11857));
	notech_inv i_15719(.A(\dir1[19] ), .Z(n_11858));
	notech_inv i_15720(.A(\dir1[20] ), .Z(n_11859));
	notech_inv i_15721(.A(\dir1[21] ), .Z(n_11860));
	notech_inv i_15722(.A(\dir1[22] ), .Z(n_11861));
	notech_inv i_15723(.A(\dir1[23] ), .Z(n_11862));
	notech_inv i_15724(.A(\dir1[24] ), .Z(n_11863));
	notech_inv i_15725(.A(\dir1[25] ), .Z(n_11864));
	notech_inv i_15726(.A(\dir1[26] ), .Z(n_11865));
	notech_inv i_15727(.A(n_494), .Z(n_11866));
	notech_inv i_15728(.A(\dir1[27] ), .Z(n_11867));
	notech_inv i_15729(.A(\dir1[28] ), .Z(n_11868));
	notech_inv i_15730(.A(\dir1[29] ), .Z(n_11869));
	notech_inv i_15731(.A(n_59950), .Z(n_11870));
	notech_inv i_15732(.A(n_536), .Z(n_11871));
	notech_inv i_15733(.A(n_571), .Z(n_11872));
	notech_inv i_15734(.A(\tab12[10] ), .Z(n_11873));
	notech_inv i_15735(.A(\tab12[11] ), .Z(n_11874));
	notech_inv i_15736(.A(\tab12[12] ), .Z(n_11875));
	notech_inv i_15737(.A(\tab12[13] ), .Z(n_11876));
	notech_inv i_15738(.A(\tab12[14] ), .Z(n_11877));
	notech_inv i_15739(.A(\tab12[15] ), .Z(n_11878));
	notech_inv i_15740(.A(\tab12[16] ), .Z(n_11879));
	notech_inv i_15741(.A(\tab12[17] ), .Z(n_11880));
	notech_inv i_15742(.A(n_583), .Z(n_11881));
	notech_inv i_15743(.A(\tab12[18] ), .Z(n_11882));
	notech_inv i_15744(.A(\tab12[19] ), .Z(n_11883));
	notech_inv i_15745(.A(\tab12[20] ), .Z(n_11884));
	notech_inv i_15746(.A(\tab12[21] ), .Z(n_11885));
	notech_inv i_15747(.A(\tab12[22] ), .Z(n_11886));
	notech_inv i_15748(.A(\tab12[23] ), .Z(n_11887));
	notech_inv i_15749(.A(\tab12[24] ), .Z(n_11888));
	notech_inv i_15750(.A(\tab12[25] ), .Z(n_11889));
	notech_inv i_15751(.A(\tab12[26] ), .Z(n_11890));
	notech_inv i_15752(.A(\tab12[27] ), .Z(n_11891));
	notech_inv i_15753(.A(\tab12[28] ), .Z(n_11892));
	notech_inv i_15754(.A(\tab12[29] ), .Z(n_11893));
	notech_inv i_15755(.A(hit_adr12), .Z(n_11894));
	notech_inv i_15756(.A(n_58743), .Z(n_11895));
	notech_inv i_15757(.A(n_606), .Z(n_55446));
	notech_inv i_15758(.A(\tab14[10] ), .Z(n_11897));
	notech_inv i_15759(.A(\tab14[11] ), .Z(n_11898));
	notech_inv i_15760(.A(\tab14[12] ), .Z(n_11899));
	notech_inv i_15761(.A(\tab14[13] ), .Z(n_11900));
	notech_inv i_15762(.A(\tab14[14] ), .Z(n_11901));
	notech_inv i_15763(.A(\tab14[15] ), .Z(n_11902));
	notech_inv i_15764(.A(\tab14[16] ), .Z(n_11903));
	notech_inv i_15765(.A(\tab14[17] ), .Z(n_11904));
	notech_inv i_15766(.A(\tab14[18] ), .Z(n_11905));
	notech_inv i_15767(.A(\tab14[19] ), .Z(n_11906));
	notech_inv i_15768(.A(\tab14[20] ), .Z(n_11907));
	notech_inv i_15769(.A(\tab14[21] ), .Z(n_11908));
	notech_inv i_15770(.A(\tab14[22] ), .Z(n_11909));
	notech_inv i_15771(.A(\tab14[23] ), .Z(n_11910));
	notech_inv i_15772(.A(\tab14[24] ), .Z(n_11911));
	notech_inv i_15773(.A(\tab14[25] ), .Z(n_11912));
	notech_inv i_15774(.A(\tab14[26] ), .Z(n_11913));
	notech_inv i_15775(.A(\tab14[27] ), .Z(n_11914));
	notech_inv i_15776(.A(\tab14[28] ), .Z(n_11915));
	notech_inv i_15777(.A(\tab14[29] ), .Z(n_11916));
	notech_inv i_15778(.A(n_59073), .Z(n_11917));
	notech_inv i_15779(.A(\nx_tab1[0] ), .Z(n_11918));
	notech_inv i_15780(.A(n_59079), .Z(n_11919));
	notech_inv i_15781(.A(\nx_tab1[1] ), .Z(n_11920));
	notech_inv i_15782(.A(n_58352), .Z(n_11921));
	notech_inv i_15783(.A(\nnx_tab1[0] ), .Z(n_11922));
	notech_inv i_15784(.A(n_58358), .Z(n_11923));
	notech_inv i_15785(.A(\nnx_tab1[1] ), .Z(n_11924));
	notech_inv i_15786(.A(\nbus_14507[0] ), .Z(n_11925));
	notech_inv i_15787(.A(\tab22[10] ), .Z(n_11926));
	notech_inv i_15788(.A(\tab22[11] ), .Z(n_11927));
	notech_inv i_15789(.A(\tab22[12] ), .Z(n_11928));
	notech_inv i_15790(.A(\tab22[13] ), .Z(n_11929));
	notech_inv i_15791(.A(\tab22[14] ), .Z(n_11930));
	notech_inv i_15792(.A(\tab22[15] ), .Z(n_11931));
	notech_inv i_15793(.A(\tab22[16] ), .Z(n_11932));
	notech_inv i_15794(.A(\tab22[17] ), .Z(n_11933));
	notech_inv i_15795(.A(\tab22[18] ), .Z(n_11934));
	notech_inv i_15796(.A(\tab22[19] ), .Z(n_11935));
	notech_inv i_15797(.A(\tab22[20] ), .Z(n_11936));
	notech_inv i_15798(.A(\tab22[21] ), .Z(n_11937));
	notech_inv i_15799(.A(\tab22[22] ), .Z(n_11938));
	notech_inv i_15800(.A(\tab22[23] ), .Z(n_11939));
	notech_inv i_15801(.A(\tab22[24] ), .Z(n_11940));
	notech_inv i_15802(.A(\tab22[25] ), .Z(n_11941));
	notech_inv i_15803(.A(\tab22[26] ), .Z(n_11942));
	notech_inv i_15804(.A(\tab22[27] ), .Z(n_11943));
	notech_inv i_15805(.A(\tab22[28] ), .Z(n_11944));
	notech_inv i_15806(.A(\tab22[29] ), .Z(n_11945));
	notech_inv i_15807(.A(hit_adr22), .Z(n_11946));
	notech_inv i_15808(.A(\tab23[10] ), .Z(n_11947));
	notech_inv i_15809(.A(\tab23[11] ), .Z(n_11948));
	notech_inv i_15810(.A(\tab23[12] ), .Z(n_11949));
	notech_inv i_15811(.A(\tab23[13] ), .Z(n_11950));
	notech_inv i_15812(.A(\tab23[14] ), .Z(n_11951));
	notech_inv i_15813(.A(\tab23[15] ), .Z(n_11952));
	notech_inv i_15814(.A(\tab23[16] ), .Z(n_11953));
	notech_inv i_15815(.A(\tab23[17] ), .Z(n_11954));
	notech_inv i_15816(.A(\tab23[18] ), .Z(n_11955));
	notech_inv i_15817(.A(\tab23[19] ), .Z(n_11956));
	notech_inv i_15818(.A(\tab23[20] ), .Z(n_11957));
	notech_inv i_15819(.A(\tab23[21] ), .Z(n_11958));
	notech_inv i_15820(.A(\tab23[22] ), .Z(n_11959));
	notech_inv i_15821(.A(\tab23[23] ), .Z(n_11960));
	notech_inv i_15822(.A(\tab23[24] ), .Z(n_11961));
	notech_inv i_15823(.A(\tab23[25] ), .Z(n_11962));
	notech_inv i_15824(.A(\tab23[26] ), .Z(n_11963));
	notech_inv i_15825(.A(\tab23[27] ), .Z(n_11964));
	notech_inv i_15826(.A(\tab23[28] ), .Z(n_11965));
	notech_inv i_15827(.A(\tab23[29] ), .Z(n_11966));
	notech_inv i_15828(.A(\tab24[10] ), .Z(n_11967));
	notech_inv i_15829(.A(\tab24[11] ), .Z(n_11968));
	notech_inv i_15830(.A(\tab24[12] ), .Z(n_11969));
	notech_inv i_15831(.A(\tab24[13] ), .Z(n_11970));
	notech_inv i_15832(.A(\tab24[14] ), .Z(n_11971));
	notech_inv i_15833(.A(\tab24[15] ), .Z(n_11972));
	notech_inv i_15834(.A(\tab24[16] ), .Z(n_11973));
	notech_inv i_15835(.A(\tab24[17] ), .Z(n_11974));
	notech_inv i_15836(.A(\tab24[18] ), .Z(n_11975));
	notech_inv i_15837(.A(\tab24[19] ), .Z(n_11976));
	notech_inv i_15838(.A(\tab24[20] ), .Z(n_11977));
	notech_inv i_15839(.A(\tab24[21] ), .Z(n_11978));
	notech_inv i_15840(.A(\tab24[22] ), .Z(n_11979));
	notech_inv i_15841(.A(\tab24[23] ), .Z(n_11980));
	notech_inv i_15842(.A(\tab24[24] ), .Z(n_11981));
	notech_inv i_15843(.A(\tab24[25] ), .Z(n_11982));
	notech_inv i_15844(.A(\tab24[26] ), .Z(n_11983));
	notech_inv i_15845(.A(\tab24[27] ), .Z(n_11984));
	notech_inv i_15846(.A(\tab24[28] ), .Z(n_11985));
	notech_inv i_15847(.A(\tab24[29] ), .Z(n_11986));
	notech_inv i_15848(.A(n_58317), .Z(n_11987));
	notech_inv i_15849(.A(\nnx_tab2[0] ), .Z(n_11988));
	notech_inv i_15850(.A(n_58323), .Z(n_11989));
	notech_inv i_15851(.A(\nnx_tab2[1] ), .Z(n_11990));
	notech_inv i_15852(.A(\nbus_14506[0] ), .Z(n_11991));
	notech_inv i_15853(.A(n_59705), .Z(n_11992));
	notech_inv i_15854(.A(\nx_tab2[0] ), .Z(n_11993));
	notech_inv i_15855(.A(n_59711), .Z(n_11994));
	notech_inv i_15856(.A(\nx_tab2[1] ), .Z(n_11995));
	notech_inv i_15857(.A(n_56853), .Z(n_11996));
	notech_inv i_15858(.A(n_58612), .Z(n_11997));
	notech_inv i_15859(.A(fsm[1]), .Z(n_11998));
	notech_inv i_15860(.A(n_58618), .Z(n_11999));
	notech_inv i_15861(.A(fsm[2]), .Z(n_12000));
	notech_inv i_15862(.A(fsm[3]), .Z(n_12001));
	notech_inv i_15863(.A(n_59518), .Z(n_12002));
	notech_inv i_15864(.A(n_59524), .Z(n_12003));
	notech_inv i_15865(.A(n_59530), .Z(n_12004));
	notech_inv i_15866(.A(n_59536), .Z(n_12005));
	notech_inv i_15867(.A(n_59542), .Z(n_12006));
	notech_inv i_15868(.A(n_59548), .Z(n_12007));
	notech_inv i_15869(.A(n_59554), .Z(n_12008));
	notech_inv i_15870(.A(n_59560), .Z(n_12009));
	notech_inv i_15871(.A(n_59566), .Z(n_12010));
	notech_inv i_15872(.A(n_59572), .Z(n_12011));
	notech_inv i_15873(.A(req_miss), .Z(n_12012));
	notech_inv i_15874(.A(addr_miss[0]), .Z(n_12013));
	notech_inv i_15875(.A(addr_miss[1]), .Z(n_12014));
	notech_inv i_15876(.A(addr_miss[2]), .Z(n_12015));
	notech_inv i_15877(.A(addr_miss[3]), .Z(n_12016));
	notech_inv i_15878(.A(addr_miss[4]), .Z(n_12017));
	notech_inv i_15879(.A(addr_miss[5]), .Z(n_12018));
	notech_inv i_15880(.A(addr_miss[6]), .Z(n_12019));
	notech_inv i_15881(.A(addr_miss[7]), .Z(n_12020));
	notech_inv i_15882(.A(addr_miss[8]), .Z(n_12021));
	notech_inv i_15883(.A(addr_miss[9]), .Z(n_12022));
	notech_inv i_15884(.A(addr_miss[10]), .Z(n_12023));
	notech_inv i_15885(.A(addr_miss[11]), .Z(n_12024));
	notech_inv i_15886(.A(addr_miss[12]), .Z(n_12025));
	notech_inv i_15887(.A(wrA[12]), .Z(n_12026));
	notech_inv i_15888(.A(addr_miss[13]), .Z(n_12027));
	notech_inv i_15889(.A(wrA[13]), .Z(n_12028));
	notech_inv i_15890(.A(addr_miss[14]), .Z(n_12029));
	notech_inv i_15891(.A(wrA[14]), .Z(n_12030));
	notech_inv i_15892(.A(addr_miss[15]), .Z(n_12031));
	notech_inv i_15893(.A(wrA[15]), .Z(n_12032));
	notech_inv i_15894(.A(addr_miss[16]), .Z(n_12033));
	notech_inv i_15895(.A(wrA[16]), .Z(n_12034));
	notech_inv i_15896(.A(addr_miss[17]), .Z(n_12035));
	notech_inv i_15897(.A(wrA[17]), .Z(n_12036));
	notech_inv i_15898(.A(addr_miss[18]), .Z(n_12037));
	notech_inv i_15899(.A(wrA[18]), .Z(n_12038));
	notech_inv i_15900(.A(addr_miss[19]), .Z(n_12039));
	notech_inv i_15901(.A(wrA[19]), .Z(n_12040));
	notech_inv i_15902(.A(addr_miss[20]), .Z(n_12041));
	notech_inv i_15903(.A(wrA[20]), .Z(n_12042));
	notech_inv i_15904(.A(addr_miss[21]), .Z(n_12043));
	notech_inv i_15905(.A(wrA[21]), .Z(n_12044));
	notech_inv i_15906(.A(addr_miss[22]), .Z(n_12045));
	notech_inv i_15907(.A(wrA[22]), .Z(n_12046));
	notech_inv i_15908(.A(addr_miss[23]), .Z(n_12047));
	notech_inv i_15909(.A(wrA[23]), .Z(n_12048));
	notech_inv i_15910(.A(addr_miss[24]), .Z(n_12049));
	notech_inv i_15911(.A(wrA[24]), .Z(n_12050));
	notech_inv i_15912(.A(addr_miss[25]), .Z(n_12051));
	notech_inv i_15913(.A(wrA[25]), .Z(n_12052));
	notech_inv i_15914(.A(addr_miss[26]), .Z(n_12053));
	notech_inv i_15915(.A(wrA[26]), .Z(n_12054));
	notech_inv i_15916(.A(addr_miss[27]), .Z(n_12055));
	notech_inv i_15917(.A(wrA[27]), .Z(n_12056));
	notech_inv i_15918(.A(addr_miss[28]), .Z(n_12057));
	notech_inv i_15919(.A(wrA[28]), .Z(n_12058));
	notech_inv i_15920(.A(addr_miss[29]), .Z(n_12059));
	notech_inv i_15921(.A(wrA[29]), .Z(n_12060));
	notech_inv i_15922(.A(addr_miss[30]), .Z(n_12061));
	notech_inv i_15923(.A(wrA[30]), .Z(n_12062));
	notech_inv i_15924(.A(addr_miss[31]), .Z(n_12063));
	notech_inv i_15925(.A(wrA[31]), .Z(n_12064));
	notech_inv i_15926(.A(n_58050), .Z(n_12065));
	notech_inv i_15927(.A(n_58057), .Z(n_12066));
	notech_inv i_15928(.A(n_58064), .Z(n_12067));
	notech_inv i_15929(.A(n_58071), .Z(n_12068));
	notech_inv i_15930(.A(n_58078), .Z(n_12069));
	notech_inv i_15931(.A(n_58085), .Z(n_12070));
	notech_inv i_15932(.A(n_58092), .Z(n_12071));
	notech_inv i_15933(.A(n_58099), .Z(n_12072));
	notech_inv i_15934(.A(n_58106), .Z(n_12073));
	notech_inv i_15935(.A(n_58113), .Z(n_12074));
	notech_inv i_15936(.A(n_58120), .Z(n_12075));
	notech_inv i_15937(.A(n_58127), .Z(n_12076));
	notech_inv i_15938(.A(n_58134), .Z(n_12077));
	notech_inv i_15939(.A(n_58141), .Z(n_12078));
	notech_inv i_15940(.A(n_58148), .Z(n_12079));
	notech_inv i_15941(.A(n_58155), .Z(n_12080));
	notech_inv i_15942(.A(n_58162), .Z(n_12081));
	notech_inv i_15943(.A(n_58169), .Z(n_12082));
	notech_inv i_15944(.A(n_58176), .Z(n_12083));
	notech_inv i_15945(.A(n_58183), .Z(n_12084));
	notech_inv i_15947(.A(cr3[31]), .Z(n_12086));
	notech_inv i_15948(.A(cr3[30]), .Z(n_12087));
	notech_inv i_15949(.A(cr3[29]), .Z(n_12088));
	notech_inv i_15950(.A(cr3[28]), .Z(n_12089));
	notech_inv i_15951(.A(cr3[27]), .Z(n_12090));
	notech_inv i_15952(.A(cr3[26]), .Z(n_12091));
	notech_inv i_15953(.A(cr3[25]), .Z(n_12092));
	notech_inv i_15954(.A(cr3[24]), .Z(n_12093));
	notech_inv i_15955(.A(cr3[23]), .Z(n_12094));
	notech_inv i_15956(.A(cr3[22]), .Z(n_12095));
	notech_inv i_15957(.A(cr3[21]), .Z(n_12096));
	notech_inv i_15958(.A(cr3[20]), .Z(n_12097));
	notech_inv i_15959(.A(cr3[19]), .Z(n_12098));
	notech_inv i_15960(.A(cr3[18]), .Z(n_12099));
	notech_inv i_15961(.A(cr3[17]), .Z(n_12100));
	notech_inv i_15962(.A(cr3[16]), .Z(n_12101));
	notech_inv i_15963(.A(cr3[15]), .Z(n_12102));
	notech_inv i_15964(.A(cr3[14]), .Z(n_12103));
	notech_inv i_15965(.A(cr3[13]), .Z(n_12104));
	notech_inv i_15966(.A(cr3[12]), .Z(n_12105));
	notech_inv i_15967(.A(iDaddr[0]), .Z(n_12106));
	notech_inv i_15968(.A(iDaddr[1]), .Z(n_12107));
	notech_inv i_15969(.A(iDaddr[2]), .Z(n_12108));
	notech_inv i_15970(.A(iDaddr[3]), .Z(n_12109));
	notech_inv i_15971(.A(iDaddr[4]), .Z(n_12110));
	notech_inv i_15972(.A(iDaddr[5]), .Z(n_12111));
	notech_inv i_15973(.A(iDaddr[6]), .Z(n_12112));
	notech_inv i_15974(.A(iDaddr[7]), .Z(n_12113));
	notech_inv i_15975(.A(iDaddr[8]), .Z(n_12114));
	notech_inv i_15976(.A(iDaddr[9]), .Z(n_12115));
	notech_inv i_15977(.A(iDaddr[10]), .Z(n_12116));
	notech_inv i_15978(.A(iDaddr[11]), .Z(n_12117));
	notech_inv i_15979(.A(iDaddr[12]), .Z(n_12118));
	notech_inv i_15980(.A(iDaddr[13]), .Z(n_12119));
	notech_inv i_15981(.A(iDaddr[14]), .Z(n_12120));
	notech_inv i_15982(.A(iDaddr[15]), .Z(n_12121));
	notech_inv i_15983(.A(iDaddr[16]), .Z(n_12122));
	notech_inv i_15984(.A(iDaddr[17]), .Z(n_12123));
	notech_inv i_15985(.A(iDaddr[18]), .Z(n_12124));
	notech_inv i_15986(.A(iDaddr[19]), .Z(n_12125));
	notech_inv i_15987(.A(iDaddr[20]), .Z(n_12126));
	notech_inv i_15988(.A(iDaddr[21]), .Z(n_12127));
	notech_inv i_15989(.A(iDaddr[22]), .Z(n_12128));
	notech_inv i_15990(.A(iDaddr[23]), .Z(n_12129));
	notech_inv i_15991(.A(iDaddr[24]), .Z(n_12130));
	notech_inv i_15992(.A(iDaddr[25]), .Z(n_12131));
	notech_inv i_15993(.A(iDaddr[26]), .Z(n_12132));
	notech_inv i_15994(.A(iDaddr[27]), .Z(n_12133));
	notech_inv i_15995(.A(iDaddr[28]), .Z(n_12134));
	notech_inv i_15996(.A(iDaddr[29]), .Z(n_12135));
	notech_inv i_15997(.A(iDaddr[30]), .Z(n_12136));
	notech_inv i_15998(.A(iDaddr[31]), .Z(n_12137));
	notech_inv i_15999(.A(cs[1]), .Z(n_12138));
	notech_inv i_16000(.A(cr0[16]), .Z(n_12139));
	notech_inv i_16001(.A(n_977), .Z(n_12140));
	notech_inv i_16002(.A(\dir1_0[9] ), .Z(n_12141));
	notech_inv i_16003(.A(\dir1_0[8] ), .Z(n_12142));
	notech_inv i_16004(.A(\dir1_0[7] ), .Z(n_12143));
	notech_inv i_16005(.A(\dir1_0[6] ), .Z(n_12144));
	notech_inv i_16006(.A(\dir1_0[5] ), .Z(n_12145));
	notech_inv i_16007(.A(\dir1_0[4] ), .Z(n_12146));
	notech_inv i_16008(.A(\dir1_0[3] ), .Z(n_12147));
	notech_inv i_16009(.A(\dir1_0[2] ), .Z(n_12148));
	notech_inv i_16010(.A(\dir1_0[1] ), .Z(n_12149));
	notech_inv i_16011(.A(\dir1_0[0] ), .Z(n_12150));
	notech_inv i_16012(.A(\tab11_0[9] ), .Z(n_12151));
	notech_inv i_16013(.A(\tab11_0[8] ), .Z(n_12152));
	notech_inv i_16014(.A(\tab11_0[7] ), .Z(n_12153));
	notech_inv i_16015(.A(\tab11_0[6] ), .Z(n_12154));
	notech_inv i_16016(.A(\tab11_0[5] ), .Z(n_12155));
	notech_inv i_16017(.A(\tab11_0[4] ), .Z(n_12156));
	notech_inv i_16018(.A(\tab11_0[3] ), .Z(n_12157));
	notech_inv i_16019(.A(\tab11_0[2] ), .Z(n_12158));
	notech_inv i_16020(.A(\tab11_0[1] ), .Z(n_12159));
	notech_inv i_16021(.A(\tab11_0[0] ), .Z(n_12160));
	notech_inv i_16022(.A(oread_ack101000), .Z(oread_ack));
	notech_inv i_16023(.A(hit_tab12), .Z(n_12162));
	notech_inv i_16024(.A(hit_tab23), .Z(n_12163));
	notech_inv i_16025(.A(\hit_dir1[7] ), .Z(n_12164));
	notech_inv i_16026(.A(n_58734), .Z(n_12165));
	notech_inv i_16027(.A(n_62898), .Z(n_12166));
	notech_inv i_16028(.A(iread_ack), .Z(n_12167));
	cmp14_9 t11(.ina({\tab11[33] , \tab11[32] , UNCONNECTED_000, \tab11[30] 
		, \tab11[9] , \tab11[8] , \tab11[7] , \tab11[6] , \tab11[5] , \tab11[4] 
		, \tab11[3] , \tab11[2] , \tab11[1] , \tab11[0] }), .inb({
		UNCONNECTED_001, n_55446, UNCONNECTED_002, iwrite_req, \tab11_0[9] 
		, \tab11_0[8] , \tab11_0[7] , \tab11_0[6] , \tab11_0[5] , \tab11_0[4] 
		, \tab11_0[3] , \tab11_0[2] , \tab11_0[1] , \tab11_0[0] }), .out
		(hit_tab11), .out2(hit_add11));
	cmp14_8 t24(.ina({\tab24[33] , \tab24[32] , UNCONNECTED_003, \tab24[30] 
		, \tab24[9] , \tab24[8] , \tab24[7] , \tab24[6] , \tab24[5] , \tab24[4] 
		, \tab24[3] , \tab24[2] , \tab24[1] , \tab24[0] }), .inb({
		UNCONNECTED_004, n_55446, UNCONNECTED_005, iwrite_req, \tab11_0[9] 
		, \tab11_0[8] , \tab11_0[7] , \tab11_0[6] , \tab11_0[5] , \tab11_0[4] 
		, \tab11_0[3] , \tab11_0[2] , \tab11_0[1] , \tab11_0[0] }), .out
		(hit_tab24), .out2(hit_add24));
	cmp14_7 t23(.ina({\tab23[33] , \tab23[32] , UNCONNECTED_006, \tab23[30] 
		, \tab23[9] , \tab23[8] , \tab23[7] , \tab23[6] , \tab23[5] , \tab23[4] 
		, \tab23[3] , \tab23[2] , \tab23[1] , \tab23[0] }), .inb({
		UNCONNECTED_007, n_55446, UNCONNECTED_008, iwrite_req, \tab11_0[9] 
		, \tab11_0[8] , \tab11_0[7] , \tab11_0[6] , \tab11_0[5] , \tab11_0[4] 
		, \tab11_0[3] , \tab11_0[2] , \tab11_0[1] , \tab11_0[0] }), .out
		(hit_tab23), .out2(hit_add23));
	cmp14_6 t22(.ina({\tab22[33] , \tab22[32] , UNCONNECTED_009, \tab22[30] 
		, \tab22[9] , \tab22[8] , \tab22[7] , \tab22[6] , \tab22[5] , \tab22[4] 
		, \tab22[3] , \tab22[2] , \tab22[1] , \tab22[0] }), .inb({
		UNCONNECTED_010, n_55446, UNCONNECTED_011, iwrite_req, \tab11_0[9] 
		, \tab11_0[8] , \tab11_0[7] , \tab11_0[6] , \tab11_0[5] , \tab11_0[4] 
		, \tab11_0[3] , \tab11_0[2] , \tab11_0[1] , \tab11_0[0] }), .out
		(hit_tab22), .out2(hit_add22));
	cmp14_5 t21(.ina({\tab21[33] , \tab21[32] , UNCONNECTED_012, \tab21[30] 
		, \tab21[9] , \tab21[8] , \tab21[7] , \tab21[6] , \tab21[5] , \tab21[4] 
		, \tab21[3] , \tab21[2] , \tab21[1] , \tab21[0] }), .inb({
		UNCONNECTED_013, n_55446, UNCONNECTED_014, iwrite_req, \tab11_0[9] 
		, \tab11_0[8] , \tab11_0[7] , \tab11_0[6] , \tab11_0[5] , \tab11_0[4] 
		, \tab11_0[3] , \tab11_0[2] , \tab11_0[1] , \tab11_0[0] }), .out
		(hit_tab21), .out2(hit_add21));
	cmp14_4 t14(.ina({\tab14[33] , \tab14[32] , UNCONNECTED_015, \tab14[30] 
		, \tab14[9] , \tab14[8] , \tab14[7] , \tab14[6] , \tab14[5] , \tab14[4] 
		, \tab14[3] , \tab14[2] , \tab14[1] , \tab14[0] }), .inb({
		UNCONNECTED_016, n_55446, UNCONNECTED_017, iwrite_req, \tab11_0[9] 
		, \tab11_0[8] , \tab11_0[7] , \tab11_0[6] , \tab11_0[5] , \tab11_0[4] 
		, \tab11_0[3] , \tab11_0[2] , \tab11_0[1] , \tab11_0[0] }), .out
		(hit_tab14), .out2(hit_add14));
	cmp14_3 t13(.ina({\tab13[33] , \tab13[32] , UNCONNECTED_018, \tab13[30] 
		, \tab13[9] , \tab13[8] , \tab13[7] , \tab13[6] , \tab13[5] , \tab13[4] 
		, \tab13[3] , \tab13[2] , \tab13[1] , \tab13[0] }), .inb({
		UNCONNECTED_019, n_55446, UNCONNECTED_020, iwrite_req, \tab11_0[9] 
		, \tab11_0[8] , \tab11_0[7] , \tab11_0[6] , \tab11_0[5] , \tab11_0[4] 
		, \tab11_0[3] , \tab11_0[2] , \tab11_0[1] , \tab11_0[0] }), .out
		(hit_tab13), .out2(hit_add13));
	cmp14_2 t12(.ina({\tab12[33] , \tab12[32] , UNCONNECTED_021, \tab12[30] 
		, \tab12[9] , \tab12[8] , \tab12[7] , \tab12[6] , \tab12[5] , \tab12[4] 
		, \tab12[3] , \tab12[2] , \tab12[1] , \tab12[0] }), .inb({
		UNCONNECTED_022, n_55446, UNCONNECTED_023, iwrite_req, \tab11_0[9] 
		, \tab11_0[8] , \tab11_0[7] , \tab11_0[6] , \tab11_0[5] , \tab11_0[4] 
		, \tab11_0[3] , \tab11_0[2] , \tab11_0[1] , \tab11_0[0] }), .out
		(hit_tab12), .out2(hit_add12));
	cmp14_1 d2(.ina({\dir2[33] , UNCONNECTED_024, UNCONNECTED_025, 
		UNCONNECTED_026, \dir2[9] , \dir2[8] , \dir2[7] , \dir2[6] , \dir2[5] 
		, \dir2[4] , \dir2[3] , \dir2[2] , \dir2[1] , \dir2[0] }), .inb(
		{UNCONNECTED_027, UNCONNECTED_028, UNCONNECTED_029, 
		UNCONNECTED_030, \dir1_0[9] , \dir1_0[8] , \dir1_0[7] , \dir1_0[6] 
		, \dir1_0[5] , \dir1_0[4] , \dir1_0[3] , \dir1_0[2] , \dir1_0[1] 
		, \dir1_0[0] }), .out(hit_dir2));
	cmp14_0 d1(.ina({\dir1[33] , UNCONNECTED_031, UNCONNECTED_032, 
		UNCONNECTED_033, \dir1[9] , \dir1[8] , \dir1[7] , \dir1[6] , \dir1[5] 
		, \dir1[4] , \dir1[3] , \dir1[2] , \dir1[1] , \dir1[0] }), .inb(
		{UNCONNECTED_034, UNCONNECTED_035, UNCONNECTED_036, 
		UNCONNECTED_037, \dir1_0[9] , \dir1_0[8] , \dir1_0[7] , \dir1_0[6] 
		, \dir1_0[5] , \dir1_0[4] , \dir1_0[3] , \dir1_0[2] , \dir1_0[1] 
		, \dir1_0[0] }), .out(\hit_dir1[7] ));
	AWDP_INC_23 i_78686(.O0(fsm5_cnt_0), .fsm5_cnt(fsm5_cnt));
endmodule
module AWDP_INC_422889(O0, fsm5_cnt);

	output [8:0] O0;
	input [8:0] fsm5_cnt;




	notech_ha2 i_8(.A(fsm5_cnt[8]), .B(n_86), .Z(O0[8]));
	notech_ha2 i_7(.A(fsm5_cnt[7]), .B(n_84), .Z(O0[7]), .CO(n_86));
	notech_ha2 i_6(.A(fsm5_cnt[6]), .B(n_82), .Z(O0[6]), .CO(n_84));
	notech_ha2 i_5(.A(fsm5_cnt[5]), .B(n_80), .Z(O0[5]), .CO(n_82));
	notech_ha2 i_4(.A(fsm5_cnt[4]), .B(n_78), .Z(O0[4]), .CO(n_80));
	notech_ha2 i_3(.A(fsm5_cnt[3]), .B(n_76), .Z(O0[3]), .CO(n_78));
	notech_ha2 i_2(.A(fsm5_cnt[2]), .B(n_74), .Z(O0[2]), .CO(n_76));
	notech_ha2 i_1(.A(fsm5_cnt[1]), .B(fsm5_cnt[0]), .Z(O0[1]), .CO(n_74));
	notech_inv i_0(.A(fsm5_cnt[0]), .Z(O0[0]));
endmodule
module cmp14_10(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_xor2 i_10(.A(inb[2]), .B(ina[2]), .Z(n_34));
	notech_xor2 i_9(.A(inb[4]), .B(ina[4]), .Z(n_33));
	notech_xor2 i_8(.A(inb[6]), .B(ina[6]), .Z(n_32));
	notech_xor2 i_6(.A(inb[3]), .B(ina[3]), .Z(n_31));
	notech_xor2 i_5(.A(inb[5]), .B(ina[5]), .Z(n_30));
	notech_xor2 i_4(.A(inb[7]), .B(ina[7]), .Z(n_29));
	notech_xor2 i_0(.A(inb[9]), .B(ina[9]), .Z(n_55));
	notech_xor2 i_1(.A(inb[8]), .B(ina[8]), .Z(n_56));
	notech_xor2 i_3(.A(inb[1]), .B(ina[1]), .Z(n_57));
	notech_xor2 i_7(.A(inb[0]), .B(ina[0]), .Z(n_58));
	notech_or4 i_38(.A(n_57), .B(n_56), .C(n_55), .D(ina[13]), .Z(n_61));
	notech_or4 i_37(.A(n_34), .B(n_31), .C(n_33), .D(n_30), .Z(n_66));
	notech_or4 i_39(.A(n_32), .B(n_29), .C(n_58), .D(n_66), .Z(n_67));
	notech_nor2 i_2(.A(n_67), .B(n_61), .Z(out));
endmodule
module cmp14_11(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_xor2 i_10(.A(inb[2]), .B(ina[2]), .Z(n_34));
	notech_xor2 i_9(.A(inb[4]), .B(ina[4]), .Z(n_33));
	notech_xor2 i_8(.A(inb[6]), .B(ina[6]), .Z(n_32));
	notech_xor2 i_6(.A(inb[3]), .B(ina[3]), .Z(n_31));
	notech_xor2 i_5(.A(inb[5]), .B(ina[5]), .Z(n_30));
	notech_xor2 i_4(.A(inb[7]), .B(ina[7]), .Z(n_29));
	notech_xor2 i_0(.A(inb[9]), .B(ina[9]), .Z(n_55));
	notech_xor2 i_1(.A(inb[8]), .B(ina[8]), .Z(n_56));
	notech_xor2 i_3(.A(inb[1]), .B(ina[1]), .Z(n_57));
	notech_xor2 i_7(.A(inb[0]), .B(ina[0]), .Z(n_58));
	notech_or4 i_38(.A(n_57), .B(n_56), .C(n_55), .D(ina[13]), .Z(n_61));
	notech_or4 i_37(.A(n_34), .B(n_31), .C(n_33), .D(n_30), .Z(n_66));
	notech_or4 i_39(.A(n_32), .B(n_29), .C(n_58), .D(n_66), .Z(n_67));
	notech_nor2 i_2(.A(n_67), .B(n_61), .Z(out));
endmodule
module cmp14_12(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_xor2 i_25(.A(inb[5]), .B(ina[5]), .Z(n_59));
	notech_xor2 i_26(.A(inb[4]), .B(ina[4]), .Z(n_60));
	notech_xor2 i_27(.A(inb[3]), .B(ina[3]), .Z(n_62));
	notech_xor2 i_28(.A(inb[2]), .B(ina[2]), .Z(n_63));
	notech_or4 i_38(.A(n_63), .B(n_62), .C(n_60), .D(n_59), .Z(n_65));
	notech_xor2 i_29(.A(inb[1]), .B(ina[1]), .Z(n_66));
	notech_xor2 i_30(.A(inb[0]), .B(ina[0]), .Z(n_67));
	notech_xor2 i_21(.A(inb[9]), .B(ina[9]), .Z(n_69));
	notech_xor2 i_22(.A(inb[8]), .B(ina[8]), .Z(n_70));
	notech_xor2 i_23(.A(inb[7]), .B(ina[7]), .Z(n_72));
	notech_xor2 i_24(.A(inb[6]), .B(ina[6]), .Z(n_73));
	notech_or4 i_37(.A(n_73), .B(n_72), .C(n_70), .D(n_69), .Z(n_75));
	notech_nor2 i_2(.A(ina[13]), .B(out2101008), .Z(out));
	notech_or4 i_32(.A(n_67), .B(n_66), .C(n_75), .D(n_65), .Z(out2101008)
		);
	notech_inv i_16156(.A(out2101008), .Z(out2));
endmodule
module cmp14_13(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_xor2 i_25(.A(inb[5]), .B(ina[5]), .Z(n_59));
	notech_xor2 i_26(.A(inb[4]), .B(ina[4]), .Z(n_60));
	notech_xor2 i_27(.A(inb[3]), .B(ina[3]), .Z(n_62));
	notech_xor2 i_28(.A(inb[2]), .B(ina[2]), .Z(n_63));
	notech_or4 i_38(.A(n_63), .B(n_62), .C(n_60), .D(n_59), .Z(n_65));
	notech_xor2 i_29(.A(inb[1]), .B(ina[1]), .Z(n_66));
	notech_xor2 i_30(.A(inb[0]), .B(ina[0]), .Z(n_67));
	notech_xor2 i_21(.A(inb[9]), .B(ina[9]), .Z(n_69));
	notech_xor2 i_22(.A(inb[8]), .B(ina[8]), .Z(n_70));
	notech_xor2 i_23(.A(inb[7]), .B(ina[7]), .Z(n_72));
	notech_xor2 i_24(.A(inb[6]), .B(ina[6]), .Z(n_73));
	notech_or4 i_37(.A(n_73), .B(n_72), .C(n_70), .D(n_69), .Z(n_75));
	notech_nor2 i_2(.A(ina[13]), .B(out2101007), .Z(out));
	notech_or4 i_32(.A(n_67), .B(n_66), .C(n_75), .D(n_65), .Z(out2101007)
		);
	notech_inv i_16140(.A(out2101007), .Z(out2));
endmodule
module cmp14_14(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_xor2 i_25(.A(inb[5]), .B(ina[5]), .Z(n_59));
	notech_xor2 i_26(.A(inb[4]), .B(ina[4]), .Z(n_60));
	notech_xor2 i_27(.A(inb[3]), .B(ina[3]), .Z(n_62));
	notech_xor2 i_28(.A(inb[2]), .B(ina[2]), .Z(n_63));
	notech_or4 i_38(.A(n_63), .B(n_62), .C(n_60), .D(n_59), .Z(n_65));
	notech_xor2 i_29(.A(inb[1]), .B(ina[1]), .Z(n_66));
	notech_xor2 i_30(.A(inb[0]), .B(ina[0]), .Z(n_67));
	notech_xor2 i_21(.A(inb[9]), .B(ina[9]), .Z(n_69));
	notech_xor2 i_22(.A(inb[8]), .B(ina[8]), .Z(n_70));
	notech_xor2 i_23(.A(inb[7]), .B(ina[7]), .Z(n_72));
	notech_xor2 i_24(.A(inb[6]), .B(ina[6]), .Z(n_73));
	notech_or4 i_37(.A(n_73), .B(n_72), .C(n_70), .D(n_69), .Z(n_75));
	notech_nor2 i_2(.A(ina[13]), .B(out2101006), .Z(out));
	notech_or4 i_32(.A(n_67), .B(n_66), .C(n_75), .D(n_65), .Z(out2101006)
		);
	notech_inv i_16124(.A(out2101006), .Z(out2));
endmodule
module cmp14_15(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_xor2 i_25(.A(inb[5]), .B(ina[5]), .Z(n_59));
	notech_xor2 i_26(.A(inb[4]), .B(ina[4]), .Z(n_60));
	notech_xor2 i_27(.A(inb[3]), .B(ina[3]), .Z(n_62));
	notech_xor2 i_28(.A(inb[2]), .B(ina[2]), .Z(n_63));
	notech_or4 i_38(.A(n_63), .B(n_62), .C(n_60), .D(n_59), .Z(n_65));
	notech_xor2 i_29(.A(inb[1]), .B(ina[1]), .Z(n_66));
	notech_xor2 i_30(.A(inb[0]), .B(ina[0]), .Z(n_67));
	notech_xor2 i_21(.A(inb[9]), .B(ina[9]), .Z(n_69));
	notech_xor2 i_22(.A(inb[8]), .B(ina[8]), .Z(n_70));
	notech_xor2 i_23(.A(inb[7]), .B(ina[7]), .Z(n_72));
	notech_xor2 i_24(.A(inb[6]), .B(ina[6]), .Z(n_73));
	notech_or4 i_37(.A(n_73), .B(n_72), .C(n_70), .D(n_69), .Z(n_75));
	notech_nor2 i_2(.A(ina[13]), .B(out2101005), .Z(out));
	notech_or4 i_32(.A(n_67), .B(n_66), .C(n_75), .D(n_65), .Z(out2101005)
		);
	notech_inv i_16108(.A(out2101005), .Z(out2));
endmodule
module cmp14_16(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_xor2 i_25(.A(inb[5]), .B(ina[5]), .Z(n_59));
	notech_xor2 i_26(.A(inb[4]), .B(ina[4]), .Z(n_60));
	notech_xor2 i_27(.A(inb[3]), .B(ina[3]), .Z(n_62));
	notech_xor2 i_28(.A(inb[2]), .B(ina[2]), .Z(n_63));
	notech_or4 i_38(.A(n_63), .B(n_62), .C(n_60), .D(n_59), .Z(n_65));
	notech_xor2 i_29(.A(inb[1]), .B(ina[1]), .Z(n_66));
	notech_xor2 i_30(.A(inb[0]), .B(ina[0]), .Z(n_67));
	notech_xor2 i_21(.A(inb[9]), .B(ina[9]), .Z(n_69));
	notech_xor2 i_22(.A(inb[8]), .B(ina[8]), .Z(n_70));
	notech_xor2 i_23(.A(inb[7]), .B(ina[7]), .Z(n_72));
	notech_xor2 i_24(.A(inb[6]), .B(ina[6]), .Z(n_73));
	notech_or4 i_37(.A(n_73), .B(n_72), .C(n_70), .D(n_69), .Z(n_75));
	notech_nor2 i_2(.A(ina[13]), .B(out2101004), .Z(out));
	notech_or4 i_32(.A(n_67), .B(n_66), .C(n_75), .D(n_65), .Z(out2101004)
		);
	notech_inv i_16092(.A(out2101004), .Z(out2));
endmodule
module cmp14_17(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_xor2 i_25(.A(inb[5]), .B(ina[5]), .Z(n_59));
	notech_xor2 i_26(.A(inb[4]), .B(ina[4]), .Z(n_60));
	notech_xor2 i_27(.A(inb[3]), .B(ina[3]), .Z(n_62));
	notech_xor2 i_28(.A(inb[2]), .B(ina[2]), .Z(n_63));
	notech_or4 i_38(.A(n_63), .B(n_62), .C(n_60), .D(n_59), .Z(n_65));
	notech_xor2 i_29(.A(inb[1]), .B(ina[1]), .Z(n_66));
	notech_xor2 i_30(.A(inb[0]), .B(ina[0]), .Z(n_67));
	notech_xor2 i_21(.A(inb[9]), .B(ina[9]), .Z(n_69));
	notech_xor2 i_22(.A(inb[8]), .B(ina[8]), .Z(n_70));
	notech_xor2 i_23(.A(inb[7]), .B(ina[7]), .Z(n_72));
	notech_xor2 i_24(.A(inb[6]), .B(ina[6]), .Z(n_73));
	notech_or4 i_37(.A(n_73), .B(n_72), .C(n_70), .D(n_69), .Z(n_75));
	notech_nor2 i_2(.A(ina[13]), .B(out2101003), .Z(out));
	notech_or4 i_32(.A(n_67), .B(n_66), .C(n_75), .D(n_65), .Z(out2101003)
		);
	notech_inv i_16076(.A(out2101003), .Z(out2));
endmodule
module cmp14_18(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_xor2 i_25(.A(inb[5]), .B(ina[5]), .Z(n_59));
	notech_xor2 i_26(.A(inb[4]), .B(ina[4]), .Z(n_60));
	notech_xor2 i_27(.A(inb[3]), .B(ina[3]), .Z(n_62));
	notech_xor2 i_28(.A(inb[2]), .B(ina[2]), .Z(n_63));
	notech_or4 i_38(.A(n_63), .B(n_62), .C(n_60), .D(n_59), .Z(n_65));
	notech_xor2 i_29(.A(inb[1]), .B(ina[1]), .Z(n_66));
	notech_xor2 i_30(.A(inb[0]), .B(ina[0]), .Z(n_67));
	notech_xor2 i_21(.A(inb[9]), .B(ina[9]), .Z(n_69));
	notech_xor2 i_22(.A(inb[8]), .B(ina[8]), .Z(n_70));
	notech_xor2 i_23(.A(inb[7]), .B(ina[7]), .Z(n_72));
	notech_xor2 i_24(.A(inb[6]), .B(ina[6]), .Z(n_73));
	notech_or4 i_37(.A(n_73), .B(n_72), .C(n_70), .D(n_69), .Z(n_75));
	notech_nor2 i_2(.A(ina[13]), .B(out2101002), .Z(out));
	notech_or4 i_32(.A(n_67), .B(n_66), .C(n_75), .D(n_65), .Z(out2101002)
		);
	notech_inv i_16060(.A(out2101002), .Z(out2));
endmodule
module cmp14_19(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_xor2 i_25(.A(inb[5]), .B(ina[5]), .Z(n_59));
	notech_xor2 i_26(.A(inb[4]), .B(ina[4]), .Z(n_60));
	notech_xor2 i_27(.A(inb[3]), .B(ina[3]), .Z(n_62));
	notech_xor2 i_28(.A(inb[2]), .B(ina[2]), .Z(n_63));
	notech_or4 i_38(.A(n_63), .B(n_62), .C(n_60), .D(n_59), .Z(n_65));
	notech_xor2 i_29(.A(inb[1]), .B(ina[1]), .Z(n_66));
	notech_xor2 i_30(.A(inb[0]), .B(ina[0]), .Z(n_67));
	notech_xor2 i_21(.A(inb[9]), .B(ina[9]), .Z(n_69));
	notech_xor2 i_22(.A(inb[8]), .B(ina[8]), .Z(n_70));
	notech_xor2 i_23(.A(inb[7]), .B(ina[7]), .Z(n_72));
	notech_xor2 i_24(.A(inb[6]), .B(ina[6]), .Z(n_73));
	notech_or4 i_37(.A(n_73), .B(n_72), .C(n_70), .D(n_69), .Z(n_75));
	notech_nor2 i_2(.A(ina[13]), .B(out2101001), .Z(out));
	notech_or4 i_32(.A(n_67), .B(n_66), .C(n_75), .D(n_65), .Z(out2101001)
		);
	notech_inv i_16044(.A(out2101001), .Z(out2));
endmodule
module Itlb(clk, rstn, addr_phys, cr3, cr0, data_miss, iDaddr, pg_en, iwrite_data
		, owrite_data, iread_req, iread_ack, iwrite_req, iwrite_ack, iread_sz
		, oread_sz, oread_req, oread_ack, owrite_req, owrite_ack, pg_fault
		, wr_fault, cr2, flush_tlb, cs, pt_fault, busy_ram);

	input clk;
	input rstn;
	output [31:0] addr_phys;
	input [31:0] cr3;
	input [31:0] cr0;
	input [31:0] data_miss;
	input [31:0] iDaddr;
	input pg_en;
	input [31:0] iwrite_data;
	output [31:0] owrite_data;
	input iread_req;
	input iread_ack;
	input iwrite_req;
	input iwrite_ack;
	input [1:0] iread_sz;
	output [1:0] oread_sz;
	output oread_req;
	output oread_ack;
	output owrite_req;
	output owrite_ack;
	output pg_fault;
	output wr_fault;
	output [31:0] cr2;
	input flush_tlb;
	input [31:0] cs;
	output pt_fault;
	input busy_ram;

	wire [3:0] fsm;
	wire [31:0] iDaddr_f;
	wire [1:0] nx_dir;
	wire [8:0] fsm5_cnt_0;
	wire [8:0] fsm5_cnt;



	notech_inv i_14829(.A(n_62940), .Z(n_62994));
	notech_inv i_14828(.A(n_62940), .Z(n_62993));
	notech_inv i_14824(.A(n_62940), .Z(n_62989));
	notech_inv i_14820(.A(n_62940), .Z(n_62985));
	notech_inv i_14819(.A(n_62940), .Z(n_62984));
	notech_inv i_14815(.A(n_62940), .Z(n_62980));
	notech_inv i_14811(.A(n_62940), .Z(n_62976));
	notech_inv i_14810(.A(n_62940), .Z(n_62975));
	notech_inv i_14806(.A(n_62940), .Z(n_62971));
	notech_inv i_14801(.A(n_62940), .Z(n_62966));
	notech_inv i_14800(.A(n_62940), .Z(n_62965));
	notech_inv i_14796(.A(n_62940), .Z(n_62961));
	notech_inv i_14792(.A(n_62940), .Z(n_62957));
	notech_inv i_14791(.A(n_62940), .Z(n_62956));
	notech_inv i_14787(.A(n_62940), .Z(n_62952));
	notech_inv i_14783(.A(n_62940), .Z(n_62948));
	notech_inv i_14782(.A(n_62940), .Z(n_62947));
	notech_inv i_14778(.A(n_62940), .Z(n_62943));
	notech_inv i_14775(.A(clk), .Z(n_62940));
	notech_inv i_14773(.A(n_62912), .Z(n_62938));
	notech_inv i_14772(.A(n_62912), .Z(n_62937));
	notech_inv i_14768(.A(n_62912), .Z(n_62933));
	notech_inv i_14764(.A(n_62912), .Z(n_62929));
	notech_inv i_14763(.A(n_62912), .Z(n_62928));
	notech_inv i_14759(.A(n_62912), .Z(n_62924));
	notech_inv i_14755(.A(n_62912), .Z(n_62920));
	notech_inv i_14754(.A(n_62912), .Z(n_62919));
	notech_inv i_14750(.A(n_62912), .Z(n_62915));
	notech_inv i_14747(.A(clk), .Z(n_62912));
	notech_inv i_14745(.A(n_62903), .Z(n_62909));
	notech_inv i_14744(.A(n_62903), .Z(n_62908));
	notech_inv i_14740(.A(n_62903), .Z(n_62904));
	notech_inv i_14739(.A(pg_en), .Z(n_62903));
	notech_inv i_14725(.A(n_62881), .Z(n_62887));
	notech_inv i_14720(.A(n_62881), .Z(n_62882));
	notech_inv i_14719(.A(fsm[0]), .Z(n_62881));
	notech_inv i_14717(.A(n_62865), .Z(n_62878));
	notech_inv i_14715(.A(n_62865), .Z(n_62876));
	notech_inv i_14712(.A(n_62865), .Z(n_62873));
	notech_inv i_14710(.A(n_62865), .Z(n_62871));
	notech_inv i_14707(.A(n_62865), .Z(n_62868));
	notech_inv i_14705(.A(n_62865), .Z(n_62866));
	notech_inv i_14704(.A(n_551), .Z(n_62865));
	notech_inv i_14673(.A(n_62830), .Z(n_62831));
	notech_inv i_14672(.A(n_878), .Z(n_62830));
	notech_inv i_14615(.A(n_62762), .Z(n_62768));
	notech_inv i_14614(.A(n_62762), .Z(n_62767));
	notech_inv i_14610(.A(n_62762), .Z(n_62763));
	notech_inv i_14609(.A(n_886), .Z(n_62762));
	notech_inv i_14602(.A(n_62753), .Z(n_62754));
	notech_inv i_14601(.A(n_993), .Z(n_62753));
	notech_inv i_14594(.A(n_62744), .Z(n_62745));
	notech_inv i_14593(.A(n_15026), .Z(n_62744));
	notech_inv i_14103(.A(n_62206), .Z(n_62260));
	notech_inv i_14102(.A(n_62206), .Z(n_62259));
	notech_inv i_14098(.A(n_62206), .Z(n_62255));
	notech_inv i_14094(.A(n_62206), .Z(n_62251));
	notech_inv i_14093(.A(n_62206), .Z(n_62250));
	notech_inv i_14089(.A(n_62206), .Z(n_62246));
	notech_inv i_14085(.A(n_62206), .Z(n_62242));
	notech_inv i_14084(.A(n_62206), .Z(n_62241));
	notech_inv i_14080(.A(n_62206), .Z(n_62237));
	notech_inv i_14075(.A(n_62206), .Z(n_62232));
	notech_inv i_14074(.A(n_62206), .Z(n_62231));
	notech_inv i_14070(.A(n_62206), .Z(n_62227));
	notech_inv i_14066(.A(n_62206), .Z(n_62223));
	notech_inv i_14065(.A(n_62206), .Z(n_62222));
	notech_inv i_14061(.A(n_62206), .Z(n_62218));
	notech_inv i_14057(.A(n_62206), .Z(n_62214));
	notech_inv i_14056(.A(n_62206), .Z(n_62213));
	notech_inv i_14052(.A(n_62206), .Z(n_62209));
	notech_inv i_14049(.A(rstn), .Z(n_62206));
	notech_inv i_14047(.A(n_62178), .Z(n_62204));
	notech_inv i_14046(.A(n_62178), .Z(n_62203));
	notech_inv i_14042(.A(n_62178), .Z(n_62199));
	notech_inv i_14038(.A(n_62178), .Z(n_62195));
	notech_inv i_14037(.A(n_62178), .Z(n_62194));
	notech_inv i_14033(.A(n_62178), .Z(n_62190));
	notech_inv i_14029(.A(n_62178), .Z(n_62186));
	notech_inv i_14028(.A(n_62178), .Z(n_62185));
	notech_inv i_14024(.A(n_62178), .Z(n_62181));
	notech_inv i_14021(.A(rstn), .Z(n_62178));
	notech_inv i_13944(.A(n_62091), .Z(n_62092));
	notech_inv i_13943(.A(n_885), .Z(n_62091));
	notech_inv i_13936(.A(n_62082), .Z(n_62083));
	notech_inv i_13935(.A(n_890), .Z(n_62082));
	notech_inv i_13418(.A(n_61584), .Z(n_61585));
	notech_inv i_13417(.A(n_853), .Z(n_61584));
	notech_inv i_13414(.A(n_61575), .Z(n_61580));
	notech_inv i_13410(.A(n_61575), .Z(n_61576));
	notech_inv i_13409(.A(data_miss[0]), .Z(n_61575));
	notech_inv i_13198(.A(n_61262), .Z(n_61263));
	notech_inv i_13197(.A(\nbus_14016[0] ), .Z(n_61262));
	notech_inv i_13188(.A(n_61251), .Z(n_61252));
	notech_inv i_13187(.A(\nbus_14023[0] ), .Z(n_61251));
	notech_inv i_13178(.A(n_61240), .Z(n_61241));
	notech_inv i_13177(.A(\nbus_14019[0] ), .Z(n_61240));
	notech_inv i_13168(.A(n_61229), .Z(n_61230));
	notech_inv i_13167(.A(\nbus_14039[0] ), .Z(n_61229));
	notech_inv i_13158(.A(n_61218), .Z(n_61219));
	notech_inv i_13157(.A(\nbus_14025[0] ), .Z(n_61218));
	notech_inv i_13148(.A(n_61207), .Z(n_61208));
	notech_inv i_13147(.A(\nbus_14024[0] ), .Z(n_61207));
	notech_inv i_13138(.A(n_61196), .Z(n_61197));
	notech_inv i_13137(.A(\nbus_14042[0] ), .Z(n_61196));
	notech_inv i_13128(.A(n_61185), .Z(n_61186));
	notech_inv i_13127(.A(\nbus_14038[0] ), .Z(n_61185));
	notech_inv i_13118(.A(n_61174), .Z(n_61175));
	notech_inv i_13117(.A(\nbus_14026[0] ), .Z(n_61174));
	notech_inv i_13108(.A(n_61163), .Z(n_61164));
	notech_inv i_13107(.A(\nbus_14040[0] ), .Z(n_61163));
	notech_inv i_13079(.A(\nbus_14022[0] ), .Z(n_61133));
	notech_inv i_13074(.A(\nbus_14022[0] ), .Z(n_61128));
	notech_inv i_7793(.A(n_55505), .Z(n_55506));
	notech_inv i_7792(.A(n_808), .Z(n_55505));
	notech_ao3 i_68(.A(n_15145), .B(n_15116), .C(hit_adr24), .Z(n_492));
	notech_nor2 i_66(.A(hit_adr24), .B(\nx_tab2[0] ), .Z(n_490));
	notech_nor2 i_468(.A(hit_adr23), .B(n_490), .Z(n_489));
	notech_nor2 i_78(.A(hit_adr22), .B(n_489), .Z(n_487));
	notech_nand3 i_465(.A(n_61580), .B(n_875), .C(n_891), .Z(n_485));
	notech_or4 i_464(.A(n_899), .B(n_919), .C(n_15193), .D(\nx_tab1[1] ), .Z
		(n_484));
	notech_or4 i_463(.A(n_899), .B(n_919), .C(n_15195), .D(\nx_tab1[0] ), .Z
		(n_483));
	notech_or4 i_462(.A(n_899), .B(n_919), .C(n_15195), .D(n_15193), .Z(n_482
		));
	notech_xor2 i_79(.A(\nnx_tab1[1] ), .B(n_15188), .Z(n_478));
	notech_or4 i_73(.A(hit_adr13), .B(hit_adr14), .C(hit_adr12), .D(hit_adr11
		), .Z(n_476));
	notech_ao3 i_69(.A(n_15195), .B(n_15166), .C(hit_adr14), .Z(n_471));
	notech_nor2 i_67(.A(hit_adr14), .B(\nx_tab1[0] ), .Z(n_469));
	notech_nor2 i_452(.A(hit_adr13), .B(n_469), .Z(n_468));
	notech_nor2 i_80(.A(hit_adr12), .B(n_468), .Z(n_466));
	notech_or4 i_449(.A(n_899), .B(n_919), .C(\nx_tab1[1] ), .D(\nx_tab1[0] 
		), .Z(n_464));
	notech_and2 i_61(.A(fsm5_cnt[7]), .B(n_387), .Z(n_463));
	notech_or4 i_448(.A(fsm5_cnt[8]), .B(n_15341), .C(n_930), .D(n_463), .Z(n_462
		));
	notech_nor2 i_74(.A(n_463), .B(fsm5_cnt[8]), .Z(n_461));
	notech_nand2 i_445(.A(fsm[2]), .B(fsm[1]), .Z(n_459));
	notech_and3 i_51(.A(data_miss[5]), .B(iread_req), .C(n_61580), .Z(n_458)
		);
	notech_and2 i_82(.A(data_miss[5]), .B(n_61580), .Z(n_457));
	notech_ao3 i_85(.A(n_905), .B(iread_req), .C(busy_ram), .Z(n_454));
	notech_mux2 i_84(.S(fsm[3]), .A(n_459), .B(n_62887), .Z(n_453));
	notech_ao4 i_83(.A(n_62887), .B(n_889), .C(n_934), .D(n_896), .Z(n_452)
		);
	notech_or2 i_433(.A(iwrite_ack), .B(n_15218), .Z(n_450));
	notech_nor2 i_58(.A(data_miss[5]), .B(n_15284), .Z(n_449));
	notech_nand2 i_87(.A(n_948), .B(n_450), .Z(n_447));
	notech_mux2 i_86(.S(fsm[3]), .A(n_15027), .B(iwrite_ack), .Z(n_445));
	notech_nand3 i_427(.A(n_62887), .B(cr3[31]), .C(n_885), .Z(n_443));
	notech_nand3 i_424(.A(n_62887), .B(n_885), .C(cr3[30]), .Z(n_442));
	notech_nand3 i_421(.A(n_62887), .B(n_885), .C(cr3[29]), .Z(n_441));
	notech_nand3 i_418(.A(n_62887), .B(n_885), .C(cr3[28]), .Z(n_440));
	notech_nand3 i_415(.A(n_62887), .B(n_885), .C(cr3[27]), .Z(n_439));
	notech_nand3 i_412(.A(n_62887), .B(n_885), .C(cr3[26]), .Z(n_438));
	notech_nand3 i_409(.A(n_62887), .B(n_885), .C(cr3[25]), .Z(n_437));
	notech_nand3 i_406(.A(n_62887), .B(n_885), .C(cr3[24]), .Z(n_436));
	notech_nand3 i_403(.A(n_62887), .B(n_885), .C(cr3[23]), .Z(n_435));
	notech_nand3 i_400(.A(n_62887), .B(n_885), .C(cr3[22]), .Z(n_434));
	notech_nand3 i_397(.A(n_62887), .B(n_885), .C(cr3[21]), .Z(n_433));
	notech_nand3 i_394(.A(n_62887), .B(n_62092), .C(cr3[20]), .Z(n_432));
	notech_nand3 i_391(.A(n_62887), .B(n_62092), .C(cr3[19]), .Z(n_431));
	notech_nand3 i_388(.A(n_62887), .B(n_62092), .C(cr3[18]), .Z(n_430));
	notech_nand3 i_385(.A(n_62887), .B(n_62092), .C(cr3[17]), .Z(n_429));
	notech_nand3 i_382(.A(n_62887), .B(n_62092), .C(cr3[16]), .Z(n_428));
	notech_nand3 i_379(.A(n_62887), .B(n_62092), .C(cr3[15]), .Z(n_427));
	notech_nand3 i_376(.A(n_62882), .B(n_885), .C(cr3[14]), .Z(n_426));
	notech_nand3 i_373(.A(n_62882), .B(n_62092), .C(cr3[13]), .Z(n_425));
	notech_nand3 i_370(.A(n_62882), .B(n_62092), .C(cr3[12]), .Z(n_424));
	notech_nand3 i_344(.A(n_62908), .B(\wrA[2] ), .C(n_62768), .Z(n_400));
	notech_nor2 i_27(.A(n_972), .B(n_15341), .Z(n_399));
	notech_nand3 i_341(.A(n_62908), .B(n_62767), .C(\wrA[3] ), .Z(n_398));
	notech_nand3 i_338(.A(n_62909), .B(n_62768), .C(\wrA[4] ), .Z(n_397));
	notech_nand3 i_335(.A(n_62909), .B(n_62768), .C(\wrA[5] ), .Z(n_396));
	notech_nand3 i_332(.A(n_62909), .B(n_62768), .C(\wrA[6] ), .Z(n_395));
	notech_nand3 i_329(.A(n_62908), .B(n_62767), .C(\wrA[7] ), .Z(n_394));
	notech_nand3 i_326(.A(n_62908), .B(n_62767), .C(\wrA[8] ), .Z(n_393));
	notech_nand3 i_323(.A(n_62908), .B(n_62767), .C(\wrA[9] ), .Z(n_392));
	notech_nand3 i_320(.A(n_62908), .B(n_62767), .C(\wrA[10] ), .Z(n_391));
	notech_nand3 i_317(.A(n_62908), .B(n_62767), .C(\wrA[11] ), .Z(n_390));
	notech_nand2 i_81(.A(n_459), .B(n_15218), .Z(n_389));
	notech_nao3 i_21(.A(flush_tlb), .B(n_62909), .C(n_62876), .Z(n_388));
	notech_or2 i_60(.A(fsm5_cnt[6]), .B(n_386), .Z(n_387));
	notech_and3 i_52(.A(fsm5_cnt[4]), .B(fsm5_cnt[5]), .C(n_385), .Z(n_386)
		);
	notech_or2 i_48(.A(fsm5_cnt[2]), .B(fsm5_cnt[3]), .Z(n_385));
	notech_or4 i_72(.A(hit_adr23), .B(hit_adr24), .C(hit_adr22), .D(hit_adr21
		), .Z(n_497));
	notech_xor2 i_77(.A(\nnx_tab2[1] ), .B(n_15138), .Z(n_499));
	notech_nand3 i_478(.A(n_15028), .B(\nx_tab2[1] ), .C(\nx_tab2[0] ), .Z(n_503
		));
	notech_nand3 i_479(.A(n_15028), .B(\nx_tab2[1] ), .C(n_15143), .Z(n_504)
		);
	notech_nand3 i_480(.A(\nx_tab2[0] ), .B(n_15145), .C(n_15028), .Z(n_505)
		);
	notech_nand3 i_483(.A(n_15028), .B(n_15145), .C(n_15143), .Z(n_508));
	notech_or2 i_484(.A(n_876), .B(n_875), .Z(n_509));
	notech_or4 i_503(.A(n_62882), .B(n_875), .C(n_889), .D(n_887), .Z(n_528)
		);
	notech_or4 i_506(.A(nx_dir[0]), .B(nx_dir[1]), .C(n_887), .D(n_890), .Z(n_531
		));
	notech_or4 i_507(.A(n_62882), .B(n_889), .C(n_887), .D(n_61580), .Z(n_532
		));
	notech_or4 i_830043(.A(fsm[1]), .B(fsm[3]), .C(fsm[2]), .D(n_62882), .Z(n_551
		));
	notech_nand2 i_47(.A(n_62909), .B(n_555), .Z(n_553));
	notech_or4 i_528(.A(fsm[2]), .B(n_884), .C(n_62882), .D(n_883), .Z(n_555
		));
	notech_or4 i_75(.A(hit_tab12), .B(hit_tab11), .C(hit_tab13), .D(hit_tab14
		), .Z(n_557));
	notech_or4 i_76(.A(hit_tab22), .B(hit_tab21), .C(hit_tab24), .D(hit_tab23
		), .Z(n_559));
	notech_nao3 i_96(.A(n_973), .B(\addr_miss[31] ), .C(n_62768), .Z(n_564)
		);
	notech_nao3 i_93(.A(n_994), .B(\tab22[29] ), .C(n_993), .Z(n_567));
	notech_nand3 i_90(.A(n_15026), .B(n_986), .C(\tab13[29] ), .Z(n_570));
	notech_nao3 i_107(.A(n_973), .B(\addr_miss[30] ), .C(n_62768), .Z(n_575)
		);
	notech_nao3 i_104(.A(n_994), .B(\tab22[28] ), .C(n_993), .Z(n_578));
	notech_nand3 i_101(.A(n_15026), .B(n_986), .C(\tab13[28] ), .Z(n_581));
	notech_nao3 i_118(.A(n_973), .B(\addr_miss[29] ), .C(n_62768), .Z(n_586)
		);
	notech_nao3 i_115(.A(n_994), .B(\tab22[27] ), .C(n_993), .Z(n_589));
	notech_nand3 i_112(.A(n_15026), .B(n_986), .C(\tab13[27] ), .Z(n_592));
	notech_nao3 i_129(.A(n_973), .B(\addr_miss[28] ), .C(n_62768), .Z(n_597)
		);
	notech_nao3 i_126(.A(n_994), .B(\tab22[26] ), .C(n_993), .Z(n_600));
	notech_nand3 i_123(.A(n_15026), .B(n_986), .C(\tab13[26] ), .Z(n_603));
	notech_nao3 i_140(.A(n_973), .B(\addr_miss[27] ), .C(n_62768), .Z(n_608)
		);
	notech_nao3 i_137(.A(n_994), .B(\tab22[25] ), .C(n_993), .Z(n_611));
	notech_nand3 i_134(.A(n_15026), .B(n_986), .C(\tab13[25] ), .Z(n_614));
	notech_nao3 i_151(.A(n_973), .B(\addr_miss[26] ), .C(n_62768), .Z(n_619)
		);
	notech_nao3 i_148(.A(n_994), .B(\tab22[24] ), .C(n_993), .Z(n_622));
	notech_nand3 i_145(.A(n_15026), .B(n_986), .C(\tab13[24] ), .Z(n_625));
	notech_nao3 i_162(.A(n_973), .B(\addr_miss[25] ), .C(n_62768), .Z(n_630)
		);
	notech_nao3 i_159(.A(n_994), .B(\tab22[23] ), .C(n_993), .Z(n_633));
	notech_nand3 i_156(.A(n_15026), .B(n_986), .C(\tab13[23] ), .Z(n_636));
	notech_nao3 i_173(.A(n_973), .B(\addr_miss[24] ), .C(n_62768), .Z(n_641)
		);
	notech_nao3 i_170(.A(n_994), .B(\tab22[22] ), .C(n_993), .Z(n_644));
	notech_nand3 i_167(.A(n_15026), .B(n_986), .C(\tab13[22] ), .Z(n_647));
	notech_nao3 i_184(.A(n_973), .B(\addr_miss[23] ), .C(n_62768), .Z(n_652)
		);
	notech_nao3 i_181(.A(n_994), .B(\tab22[21] ), .C(n_993), .Z(n_655));
	notech_nand3 i_178(.A(n_15026), .B(n_986), .C(\tab13[21] ), .Z(n_658));
	notech_nao3 i_195(.A(n_973), .B(\addr_miss[22] ), .C(n_62768), .Z(n_663)
		);
	notech_nao3 i_192(.A(n_994), .B(\tab22[20] ), .C(n_993), .Z(n_666));
	notech_nand3 i_189(.A(n_15026), .B(n_986), .C(\tab13[20] ), .Z(n_669));
	notech_nao3 i_206(.A(n_973), .B(\addr_miss[21] ), .C(n_62767), .Z(n_674)
		);
	notech_nao3 i_203(.A(n_994), .B(\tab22[19] ), .C(n_993), .Z(n_677));
	notech_nand3 i_200(.A(n_15026), .B(n_986), .C(\tab13[19] ), .Z(n_680));
	notech_nao3 i_217(.A(n_973), .B(\addr_miss[20] ), .C(n_62763), .Z(n_685)
		);
	notech_nao3 i_214(.A(n_994), .B(\tab22[18] ), .C(n_62754), .Z(n_688));
	notech_nand3 i_211(.A(n_62745), .B(n_986), .C(\tab13[18] ), .Z(n_691));
	notech_nao3 i_228(.A(n_973), .B(\addr_miss[19] ), .C(n_62763), .Z(n_696)
		);
	notech_nao3 i_225(.A(n_994), .B(\tab22[17] ), .C(n_62754), .Z(n_699));
	notech_nand3 i_222(.A(n_62745), .B(n_986), .C(\tab13[17] ), .Z(n_702));
	notech_nao3 i_239(.A(n_973), .B(\addr_miss[18] ), .C(n_62763), .Z(n_707)
		);
	notech_nao3 i_236(.A(n_994), .B(\tab22[16] ), .C(n_62754), .Z(n_710));
	notech_nand3 i_233(.A(n_62745), .B(n_986), .C(\tab13[16] ), .Z(n_713));
	notech_nao3 i_250(.A(n_973), .B(\addr_miss[17] ), .C(n_62763), .Z(n_718)
		);
	notech_nao3 i_247(.A(n_994), .B(\tab22[15] ), .C(n_62754), .Z(n_721));
	notech_nand3 i_244(.A(n_62745), .B(n_986), .C(\tab13[15] ), .Z(n_724));
	notech_nao3 i_261(.A(n_973), .B(\addr_miss[16] ), .C(n_62763), .Z(n_729)
		);
	notech_nao3 i_258(.A(n_994), .B(\tab22[14] ), .C(n_62754), .Z(n_732));
	notech_nand3 i_255(.A(n_62745), .B(n_986), .C(\tab13[14] ), .Z(n_735));
	notech_nao3 i_279(.A(n_973), .B(\addr_miss[15] ), .C(n_62763), .Z(n_740)
		);
	notech_nao3 i_272(.A(n_994), .B(\tab22[13] ), .C(n_62754), .Z(n_743));
	notech_nand3 i_267(.A(n_62745), .B(n_986), .C(\tab13[13] ), .Z(n_746));
	notech_nao3 i_290(.A(n_973), .B(\addr_miss[14] ), .C(n_62763), .Z(n_751)
		);
	notech_nao3 i_287(.A(n_994), .B(\tab22[12] ), .C(n_62754), .Z(n_754));
	notech_nand3 i_284(.A(n_62745), .B(n_986), .C(\tab13[12] ), .Z(n_757));
	notech_nao3 i_301(.A(n_973), .B(\addr_miss[13] ), .C(n_62763), .Z(n_762)
		);
	notech_nao3 i_298(.A(n_994), .B(\tab22[11] ), .C(n_993), .Z(n_765));
	notech_nand3 i_295(.A(n_15026), .B(n_986), .C(\tab13[11] ), .Z(n_768));
	notech_nao3 i_312(.A(\addr_miss[12] ), .B(n_973), .C(n_62763), .Z(n_773)
		);
	notech_nao3 i_309(.A(\tab22[10] ), .B(n_994), .C(n_62754), .Z(n_776));
	notech_nand3 i_306(.A(n_62745), .B(\tab13[10] ), .C(n_986), .Z(n_779));
	notech_and2 i_8(.A(\wrD[7] ), .B(n_62763), .Z(owrite_data[7]));
	notech_and2 i_7(.A(\wrD[6] ), .B(n_62767), .Z(owrite_data[6]));
	notech_and2 i_6(.A(\wrD[5] ), .B(n_62767), .Z(owrite_data[5]));
	notech_and2 i_522138(.A(\wrD[4] ), .B(n_62767), .Z(owrite_data[4]));
	notech_and2 i_4(.A(\wrD[3] ), .B(n_62767), .Z(owrite_data[3]));
	notech_and2 i_3(.A(\wrD[2] ), .B(n_62767), .Z(owrite_data[2]));
	notech_and2 i_222137(.A(\wrD[1] ), .B(n_62763), .Z(owrite_data[1]));
	notech_and2 i_1(.A(\wrD[0] ), .B(n_62763), .Z(owrite_data[0]));
	notech_nao3 i_76767(.A(n_52870), .B(n_15284), .C(n_887), .Z(n_808));
	notech_or4 i_434(.A(n_854), .B(flush_tlb), .C(n_893), .D(n_906), .Z(n_851
		));
	notech_or4 i_435(.A(fsm[2]), .B(fsm[1]), .C(n_15341), .D(n_15218), .Z(n_852
		));
	notech_nand2 i_77895(.A(n_62909), .B(n_52519), .Z(n_853));
	notech_ao4 i_49(.A(hit_dir2), .B(\hit_dir1[7] ), .C(pg_fault), .D(n_15030
		), .Z(n_854));
	notech_or4 i_439(.A(fsm[1]), .B(fsm[3]), .C(fsm[2]), .D(n_454), .Z(n_855
		));
	notech_nao3 i_444(.A(n_15218), .B(n_15027), .C(iwrite_ack), .Z(n_858));
	notech_and2 i_44(.A(iwrite_ack), .B(n_389), .Z(n_861));
	notech_and2 i_76006(.A(n_52870), .B(n_15284), .Z(n_862));
	notech_ao3 i_75994(.A(fsm5_cnt_0[0]), .B(n_929), .C(n_884), .Z(n_863));
	notech_ao3 i_75995(.A(n_929), .B(fsm5_cnt_0[1]), .C(n_884), .Z(n_864));
	notech_ao3 i_75996(.A(n_929), .B(fsm5_cnt_0[2]), .C(n_884), .Z(n_865));
	notech_ao3 i_75997(.A(n_929), .B(fsm5_cnt_0[3]), .C(n_884), .Z(n_866));
	notech_ao3 i_75998(.A(n_929), .B(fsm5_cnt_0[4]), .C(n_884), .Z(n_867));
	notech_ao3 i_75999(.A(n_929), .B(fsm5_cnt_0[5]), .C(n_884), .Z(n_868));
	notech_ao3 i_76000(.A(n_929), .B(fsm5_cnt_0[6]), .C(n_884), .Z(n_869));
	notech_ao3 i_76001(.A(n_929), .B(fsm5_cnt_0[7]), .C(n_884), .Z(n_870));
	notech_ao3 i_76002(.A(n_929), .B(fsm5_cnt_0[8]), .C(n_884), .Z(n_871));
	notech_or4 i_77995(.A(n_906), .B(n_893), .C(n_904), .D(n_905), .Z(n_872)
		);
	notech_nor2 i_76650(.A(n_896), .B(n_15331), .Z(n_873));
	notech_ao3 i_75833(.A(n_61580), .B(\dir1_0[4] ), .C(n_890), .Z(n_874));
	notech_nor2 i_330041(.A(nx_dir[0]), .B(nx_dir[1]), .Z(n_875));
	notech_or4 i_78001(.A(n_62882), .B(n_889), .C(n_887), .D(n_15284), .Z(n_876
		));
	notech_and2 i_75750(.A(iread_ack), .B(n_553), .Z(oread_ack));
	notech_reg nx_dir_reg_0(.CP(n_62971), .D(n_12176), .CD(n_62237), .Q(nx_dir
		[0]));
	notech_mux2 i_16190(.S(n_876), .A(n_875), .B(nx_dir[0]), .Z(n_12176));
	notech_nand3 i_75722(.A(n_15218), .B(n_15027), .C(n_62909), .Z(n_878));
	notech_reg nx_dir_reg_1(.CP(n_62971), .D(n_12185), .CD(n_62237), .Q(nx_dir
		[1]));
	notech_and2 i_16200(.A(n_876), .B(nx_dir[1]), .Z(n_12185));
	notech_reg iDaddr_f_reg_0(.CP(n_62971), .D(n_12188), .CD(n_62237), .Q(iDaddr_f
		[0]));
	notech_mux2 i_16206(.S(n_62876), .A(iDaddr[0]), .B(iDaddr_f[0]), .Z(n_12188
		));
	notech_reg iDaddr_f_reg_1(.CP(n_62971), .D(n_12194), .CD(n_62237), .Q(iDaddr_f
		[1]));
	notech_mux2 i_16214(.S(n_62876), .A(iDaddr[1]), .B(iDaddr_f[1]), .Z(n_12194
		));
	notech_reg iDaddr_f_reg_2(.CP(n_62966), .D(n_12200), .CD(n_62232), .Q(iDaddr_f
		[2]));
	notech_mux2 i_16222(.S(n_62873), .A(iDaddr[2]), .B(iDaddr_f[2]), .Z(n_12200
		));
	notech_reg iDaddr_f_reg_3(.CP(n_62971), .D(n_12206), .CD(n_62237), .Q(iDaddr_f
		[3]));
	notech_mux2 i_16230(.S(n_62873), .A(iDaddr[3]), .B(iDaddr_f[3]), .Z(n_12206
		));
	notech_ao4 i_75580(.A(n_15343), .B(n_15108), .C(n_15340), .D(n_15105), .Z
		(n_883));
	notech_reg iDaddr_f_reg_4(.CP(n_62971), .D(n_12212), .CD(n_62237), .Q(iDaddr_f
		[4]));
	notech_mux2 i_16238(.S(n_62876), .A(iDaddr[4]), .B(iDaddr_f[4]), .Z(n_12212
		));
	notech_or2 i_30(.A(fsm[1]), .B(fsm[3]), .Z(n_884));
	notech_reg iDaddr_f_reg_5(.CP(n_62971), .D(n_12218), .CD(n_62237), .Q(iDaddr_f
		[5]));
	notech_mux2 i_16246(.S(n_62876), .A(iDaddr[5]), .B(iDaddr_f[5]), .Z(n_12218
		));
	notech_nor2 i_59(.A(fsm[2]), .B(n_884), .Z(n_885));
	notech_reg iDaddr_f_reg_6(.CP(n_62971), .D(n_12224), .CD(n_62237), .Q(iDaddr_f
		[6]));
	notech_mux2 i_16254(.S(n_62876), .A(iDaddr[6]), .B(iDaddr_f[6]), .Z(n_12224
		));
	notech_and3 i_20(.A(fsm[2]), .B(fsm[1]), .C(n_15218), .Z(n_886));
	notech_reg iDaddr_f_reg_7(.CP(n_62971), .D(n_12230), .CD(n_62237), .Q(iDaddr_f
		[7]));
	notech_mux2 i_16262(.S(n_62876), .A(iDaddr[7]), .B(iDaddr_f[7]), .Z(n_12230
		));
	notech_nand2 i_31(.A(iread_ack), .B(n_62909), .Z(n_887));
	notech_reg iDaddr_f_reg_8(.CP(n_62971), .D(n_12236), .CD(n_62237), .Q(iDaddr_f
		[8]));
	notech_mux2 i_16270(.S(n_62876), .A(iDaddr[8]), .B(iDaddr_f[8]), .Z(n_12236
		));
	notech_reg iDaddr_f_reg_9(.CP(n_62971), .D(n_12242), .CD(n_62237), .Q(iDaddr_f
		[9]));
	notech_mux2 i_16278(.S(n_62876), .A(iDaddr[9]), .B(iDaddr_f[9]), .Z(n_12242
		));
	notech_nao3 i_18(.A(fsm[1]), .B(n_15218), .C(fsm[2]), .Z(n_889));
	notech_reg iDaddr_f_reg_10(.CP(n_62971), .D(n_12248), .CD(n_62237), .Q(iDaddr_f
		[10]));
	notech_mux2 i_16286(.S(n_62873), .A(iDaddr[10]), .B(iDaddr_f[10]), .Z(n_12248
		));
	notech_nand2 i_32(.A(n_15217), .B(n_15029), .Z(n_890));
	notech_reg iDaddr_f_reg_11(.CP(n_62971), .D(n_12254), .CD(n_62237), .Q(iDaddr_f
		[11]));
	notech_mux2 i_16294(.S(n_62873), .A(iDaddr[11]), .B(iDaddr_f[11]), .Z(n_12254
		));
	notech_ao3 i_55(.A(iread_ack), .B(n_62909), .C(n_890), .Z(n_891));
	notech_reg iDaddr_f_reg_12(.CP(n_62966), .D(\tab11_0[0] ), .CD(n_62232),
		 .Q(iDaddr_f[12]));
	notech_reg iDaddr_f_reg_13(.CP(n_62966), .D(\tab11_0[1] ), .CD(n_62232),
		 .Q(iDaddr_f[13]));
	notech_or4 i_64(.A(fsm[2]), .B(n_884), .C(n_62882), .D(n_15341), .Z(n_893
		));
	notech_reg iDaddr_f_reg_14(.CP(n_62966), .D(\tab11_0[2] ), .CD(n_62232),
		 .Q(iDaddr_f[14]));
	notech_reg iDaddr_f_reg_15(.CP(n_62966), .D(\tab11_0[3] ), .CD(n_62232),
		 .Q(iDaddr_f[15]));
	notech_nand2 i_802(.A(fsm[2]), .B(n_15217), .Z(n_895));
	notech_reg iDaddr_f_reg_16(.CP(n_62966), .D(\tab11_0[4] ), .CD(n_62232),
		 .Q(iDaddr_f[16]));
	notech_or2 i_75698(.A(n_884), .B(n_895), .Z(n_896));
	notech_reg iDaddr_f_reg_17(.CP(n_62966), .D(\tab11_0[5] ), .CD(n_62232),
		 .Q(iDaddr_f[17]));
	notech_reg iDaddr_f_reg_18(.CP(n_62966), .D(\tab11_0[6] ), .CD(n_62232),
		 .Q(iDaddr_f[18]));
	notech_reg iDaddr_f_reg_19(.CP(n_62966), .D(\tab11_0[7] ), .CD(n_62232),
		 .Q(iDaddr_f[19]));
	notech_or4 i_10(.A(n_887), .B(n_884), .C(n_895), .D(n_15284), .Z(n_899)
		);
	notech_reg iDaddr_f_reg_20(.CP(n_62966), .D(\tab11_0[8] ), .CD(n_62232),
		 .Q(iDaddr_f[20]));
	notech_nand2 i_19(.A(hit_dir2), .B(n_15340), .Z(n_900));
	notech_reg iDaddr_f_reg_21(.CP(n_62966), .D(\tab11_0[9] ), .CD(n_62232),
		 .Q(iDaddr_f[21]));
	notech_or4 i_33(.A(n_896), .B(n_887), .C(n_900), .D(n_15284), .Z(n_901)
		);
	notech_reg iDaddr_f_reg_22(.CP(n_62966), .D(\dir1_0[0] ), .CD(n_62232), 
		.Q(iDaddr_f[22]));
	notech_reg iDaddr_f_reg_23(.CP(n_62966), .D(\dir1_0[1] ), .CD(n_62232), 
		.Q(iDaddr_f[23]));
	notech_reg iDaddr_f_reg_24(.CP(n_62966), .D(\dir1_0[2] ), .CD(n_62232), 
		.Q(iDaddr_f[24]));
	notech_nao3 i_798(.A(n_883), .B(n_15344), .C(flush_tlb), .Z(n_904));
	notech_reg iDaddr_f_reg_25(.CP(n_62966), .D(\dir1_0[3] ), .CD(n_62232), 
		.Q(iDaddr_f[25]));
	notech_and2 i_26(.A(n_15343), .B(n_15340), .Z(n_905));
	notech_reg iDaddr_f_reg_26(.CP(n_62966), .D(\dir1_0[4] ), .CD(n_62232), 
		.Q(iDaddr_f[26]));
	notech_or2 i_45(.A(busy_ram), .B(n_15342), .Z(n_906));
	notech_reg iDaddr_f_reg_27(.CP(n_62971), .D(\dir1_0[5] ), .CD(n_62237), 
		.Q(iDaddr_f[27]));
	notech_reg iDaddr_f_reg_28(.CP(n_62975), .D(\dir1_0[6] ), .CD(n_62241), 
		.Q(iDaddr_f[28]));
	notech_reg iDaddr_f_reg_29(.CP(n_62975), .D(\dir1_0[7] ), .CD(n_62241), 
		.Q(iDaddr_f[29]));
	notech_reg iDaddr_f_reg_30(.CP(n_62975), .D(\dir1_0[8] ), .CD(n_62241), 
		.Q(iDaddr_f[30]));
	notech_reg iDaddr_f_reg_31(.CP(n_62975), .D(\dir1_0[9] ), .CD(n_62241), 
		.Q(iDaddr_f[31]));
	notech_reg_set dir1_reg_0(.CP(n_62975), .D(n_12380), .SD(n_62241), .Q(\dir1[0] 
		));
	notech_mux2 i_16462(.S(\nbus_14024[0] ), .A(\dir1[0] ), .B(n_52302), .Z(n_12380
		));
	notech_nand2 i_75694(.A(n_62882), .B(n_15029), .Z(n_912));
	notech_reg_set dir1_reg_1(.CP(n_62975), .D(n_12386), .SD(n_62241), .Q(\dir1[1] 
		));
	notech_mux2 i_16470(.S(\nbus_14024[0] ), .A(\dir1[1] ), .B(n_52308), .Z(n_12386
		));
	notech_nao3 i_29(.A(n_62882), .B(n_62909), .C(n_889), .Z(n_913));
	notech_reg_set dir1_reg_2(.CP(n_62975), .D(n_12392), .SD(n_62241), .Q(\dir1[2] 
		));
	notech_mux2 i_16478(.S(\nbus_14024[0] ), .A(\dir1[2] ), .B(n_52314), .Z(n_12392
		));
	notech_reg_set dir1_reg_3(.CP(n_62976), .D(n_12398), .SD(n_62242), .Q(\dir1[3] 
		));
	notech_mux2 i_16486(.S(\nbus_14024[0] ), .A(\dir1[3] ), .B(n_52320), .Z(n_12398
		));
	notech_reg dir1_reg_4(.CP(n_62976), .D(n_12404), .CD(n_62242), .Q(\dir1[4] 
		));
	notech_mux2 i_16494(.S(\nbus_14024[0] ), .A(\dir1[4] ), .B(n_874), .Z(n_12404
		));
	notech_or2 i_53(.A(n_912), .B(hit_adr21), .Z(n_916));
	notech_reg_set dir1_reg_5(.CP(n_62976), .D(n_12410), .SD(n_62242), .Q(\dir1[5] 
		));
	notech_mux2 i_16502(.S(\nbus_14024[0] ), .A(\dir1[5] ), .B(n_52332), .Z(n_12410
		));
	notech_or2 i_789(.A(hit_adr22), .B(n_916), .Z(n_917));
	notech_reg_set dir1_reg_6(.CP(n_62976), .D(n_12416), .SD(n_62242), .Q(\dir1[6] 
		));
	notech_mux2 i_16510(.S(\nbus_14024[0] ), .A(\dir1[6] ), .B(n_52338), .Z(n_12416
		));
	notech_reg_set dir1_reg_7(.CP(n_62976), .D(n_12422), .SD(n_62242), .Q(\dir1[7] 
		));
	notech_mux2 i_16518(.S(\nbus_14024[0] ), .A(\dir1[7] ), .B(n_52344), .Z(n_12422
		));
	notech_nand2 i_17(.A(\hit_dir1[7] ), .B(n_15343), .Z(n_919));
	notech_reg_set dir1_reg_8(.CP(n_62976), .D(n_12428), .SD(n_62242), .Q(\dir1[8] 
		));
	notech_mux2 i_16526(.S(\nbus_14024[0] ), .A(\dir1[8] ), .B(n_52350), .Z(n_12428
		));
	notech_or4 i_34(.A(n_896), .B(n_887), .C(n_919), .D(n_15284), .Z(n_920)
		);
	notech_reg_set dir1_reg_9(.CP(n_62976), .D(n_12434), .SD(n_62242), .Q(\dir1[9] 
		));
	notech_mux2 i_16534(.S(\nbus_14024[0] ), .A(\dir1[9] ), .B(n_52356), .Z(n_12434
		));
	notech_reg_set dir1_reg_10(.CP(n_62975), .D(n_12440), .SD(n_62241), .Q(\dir1[10] 
		));
	notech_mux2 i_16542(.S(\nbus_14024[0] ), .A(\dir1[10] ), .B(n_52362), .Z
		(n_12440));
	notech_reg_set dir1_reg_11(.CP(n_62975), .D(n_12446), .SD(n_62241), .Q(\dir1[11] 
		));
	notech_mux2 i_16550(.S(\nbus_14024[0] ), .A(\dir1[11] ), .B(n_52368), .Z
		(n_12446));
	notech_reg_set dir1_reg_12(.CP(n_62975), .D(n_12452), .SD(n_62241), .Q(\dir1[12] 
		));
	notech_mux2 i_16558(.S(\nbus_14024[0] ), .A(\dir1[12] ), .B(n_52374), .Z
		(n_12452));
	notech_reg_set dir1_reg_13(.CP(n_62975), .D(n_12458), .SD(n_62241), .Q(\dir1[13] 
		));
	notech_mux2 i_16566(.S(\nbus_14024[0] ), .A(\dir1[13] ), .B(n_52380), .Z
		(n_12458));
	notech_reg_set dir1_reg_14(.CP(n_62971), .D(n_12464), .SD(n_62237), .Q(\dir1[14] 
		));
	notech_mux2 i_16574(.S(\nbus_14024[0] ), .A(\dir1[14] ), .B(n_52386), .Z
		(n_12464));
	notech_or2 i_54(.A(n_912), .B(hit_adr11), .Z(n_926));
	notech_reg_set dir1_reg_15(.CP(n_62971), .D(n_12470), .SD(n_62237), .Q(\dir1[15] 
		));
	notech_mux2 i_16582(.S(\nbus_14024[0] ), .A(\dir1[15] ), .B(n_52392), .Z
		(n_12470));
	notech_or2 i_784(.A(hit_adr12), .B(n_926), .Z(n_927));
	notech_reg_set dir1_reg_16(.CP(n_62971), .D(n_12476), .SD(n_62237), .Q(\dir1[16] 
		));
	notech_mux2 i_16590(.S(n_61208), .A(\dir1[16] ), .B(n_52398), .Z(n_12476
		));
	notech_reg_set dir1_reg_17(.CP(n_62971), .D(n_12482), .SD(n_62237), .Q(\dir1[17] 
		));
	notech_mux2 i_16598(.S(n_61208), .A(\dir1[17] ), .B(n_52404), .Z(n_12482
		));
	notech_and2 i_782(.A(fsm[2]), .B(n_62887), .Z(n_929));
	notech_reg_set dir1_reg_18(.CP(n_62975), .D(n_12488), .SD(n_62241), .Q(\dir1[18] 
		));
	notech_mux2 i_16606(.S(n_61208), .A(\dir1[18] ), .B(n_52410), .Z(n_12488
		));
	notech_nao3 i_75701(.A(fsm[2]), .B(n_62882), .C(n_884), .Z(n_930));
	notech_reg_set dir1_reg_19(.CP(n_62975), .D(n_12494), .SD(n_62241), .Q(\dir1[19] 
		));
	notech_mux2 i_16614(.S(n_61208), .A(\dir1[19] ), .B(n_52416), .Z(n_12494
		));
	notech_reg_set dir1_reg_20(.CP(n_62975), .D(n_12500), .SD(n_62241), .Q(\dir1[20] 
		));
	notech_mux2 i_16622(.S(n_61208), .A(\dir1[20] ), .B(n_52422), .Z(n_12500
		));
	notech_nao3 i_35(.A(n_929), .B(n_62909), .C(n_884), .Z(n_932));
	notech_reg_set dir1_reg_21(.CP(n_62975), .D(n_12506), .SD(n_62241), .Q(\dir1[21] 
		));
	notech_mux2 i_16630(.S(n_61208), .A(\dir1[21] ), .B(n_52428), .Z(n_12506
		));
	notech_reg_set dir1_reg_22(.CP(n_62975), .D(n_12512), .SD(n_62241), .Q(\dir1[22] 
		));
	notech_mux2 i_16638(.S(n_61208), .A(\dir1[22] ), .B(n_52434), .Z(n_12512
		));
	notech_and2 i_28(.A(data_miss[5]), .B(iread_req), .Z(n_934));
	notech_reg_set dir1_reg_23(.CP(n_62975), .D(n_12518), .SD(n_62241), .Q(\dir1[23] 
		));
	notech_mux2 i_16646(.S(n_61208), .A(\dir1[23] ), .B(n_52440), .Z(n_12518
		));
	notech_ao4 i_769(.A(n_896), .B(n_458), .C(n_889), .D(n_457), .Z(n_935)
		);
	notech_reg_set dir1_reg_24(.CP(n_62975), .D(n_12524), .SD(n_62241), .Q(\dir1[24] 
		));
	notech_mux2 i_16654(.S(n_61208), .A(\dir1[24] ), .B(n_52446), .Z(n_12524
		));
	notech_reg_set dir1_reg_25(.CP(n_62957), .D(n_12530), .SD(n_62223), .Q(\dir1[25] 
		));
	notech_mux2 i_16662(.S(n_61208), .A(\dir1[25] ), .B(n_52452), .Z(n_12530
		));
	notech_ao4 i_767(.A(n_453), .B(iwrite_ack), .C(n_452), .D(n_15284), .Z(n_937
		));
	notech_reg_set dir1_reg_26(.CP(n_62957), .D(n_12536), .SD(n_62223), .Q(\dir1[26] 
		));
	notech_mux2 i_16670(.S(n_61208), .A(\dir1[26] ), .B(n_52458), .Z(n_12536
		));
	notech_nand2 i_75687(.A(n_62882), .B(n_62092), .Z(n_938));
	notech_reg_set dir1_reg_27(.CP(n_62961), .D(n_12542), .SD(n_62227), .Q(\dir1[27] 
		));
	notech_mux2 i_16678(.S(n_61208), .A(\dir1[27] ), .B(n_52464), .Z(n_12542
		));
	notech_reg_set dir1_reg_28(.CP(n_62957), .D(n_12548), .SD(n_62223), .Q(\dir1[28] 
		));
	notech_mux2 i_16686(.S(n_61208), .A(\dir1[28] ), .B(n_52470), .Z(n_12548
		));
	notech_reg_set dir1_reg_29(.CP(n_62957), .D(n_12554), .SD(n_62223), .Q(\dir1[29] 
		));
	notech_mux2 i_16694(.S(n_61208), .A(\dir1[29] ), .B(n_52476), .Z(n_12554
		));
	notech_reg_set dir1_reg_33(.CP(n_62957), .D(n_12560), .SD(n_62223), .Q(\dir1[33] 
		));
	notech_mux2 i_16702(.S(n_61208), .A(\dir1[33] ), .B(n_52501), .Z(n_12560
		));
	notech_reg_set dir2_reg_0(.CP(n_62957), .D(n_12566), .SD(n_62223), .Q(\dir2[0] 
		));
	notech_mux2 i_16710(.S(\nbus_14016[0] ), .A(\dir2[0] ), .B(n_52302), .Z(n_12566
		));
	notech_reg_set dir2_reg_1(.CP(n_62961), .D(n_12572), .SD(n_62227), .Q(\dir2[1] 
		));
	notech_mux2 i_16718(.S(\nbus_14016[0] ), .A(\dir2[1] ), .B(n_52308), .Z(n_12572
		));
	notech_reg_set dir2_reg_2(.CP(n_62961), .D(n_12578), .SD(n_62227), .Q(\dir2[2] 
		));
	notech_mux2 i_16726(.S(\nbus_14016[0] ), .A(\dir2[2] ), .B(n_52314), .Z(n_12578
		));
	notech_and3 i_760(.A(n_852), .B(n_851), .C(n_853), .Z(n_945));
	notech_reg_set dir2_reg_3(.CP(n_62961), .D(n_12584), .SD(n_62227), .Q(\dir2[3] 
		));
	notech_mux2 i_16734(.S(\nbus_14016[0] ), .A(\dir2[3] ), .B(n_52320), .Z(n_12584
		));
	notech_reg dir2_reg_4(.CP(n_62961), .D(n_12590), .CD(n_62227), .Q(\dir2[4] 
		));
	notech_mux2 i_16742(.S(\nbus_14016[0] ), .A(\dir2[4] ), .B(n_874), .Z(n_12590
		));
	notech_or2 i_757(.A(fsm[2]), .B(fsm[3]), .Z(n_947));
	notech_reg_set dir2_reg_5(.CP(n_62961), .D(n_12596), .SD(n_62227), .Q(\dir2[5] 
		));
	notech_mux2 i_16750(.S(\nbus_14016[0] ), .A(\dir2[5] ), .B(n_52332), .Z(n_12596
		));
	notech_ao4 i_756(.A(n_458), .B(n_884), .C(n_449), .D(n_947), .Z(n_948)
		);
	notech_reg_set dir2_reg_6(.CP(n_62961), .D(n_12602), .SD(n_62227), .Q(\dir2[6] 
		));
	notech_mux2 i_16758(.S(\nbus_14016[0] ), .A(\dir2[6] ), .B(n_52338), .Z(n_12602
		));
	notech_or2 i_15(.A(\hit_dir1[7] ), .B(n_912), .Z(n_949));
	notech_reg_set dir2_reg_7(.CP(n_62961), .D(n_12608), .SD(n_62227), .Q(\dir2[7] 
		));
	notech_mux2 i_16766(.S(\nbus_14016[0] ), .A(\dir2[7] ), .B(n_52344), .Z(n_12608
		));
	notech_nao3 i_11(.A(n_62882), .B(\hit_dir1[7] ), .C(n_889), .Z(n_950));
	notech_reg_set dir2_reg_8(.CP(n_62957), .D(n_12614), .SD(n_62223), .Q(\dir2[8] 
		));
	notech_mux2 i_16774(.S(\nbus_14016[0] ), .A(\dir2[8] ), .B(n_52350), .Z(n_12614
		));
	notech_ao4 i_755(.A(n_950), .B(n_15050), .C(n_949), .D(n_15070), .Z(n_951
		));
	notech_reg_set dir2_reg_9(.CP(n_62957), .D(n_12620), .SD(n_62223), .Q(\dir2[9] 
		));
	notech_mux2 i_16782(.S(\nbus_14016[0] ), .A(\dir2[9] ), .B(n_52356), .Z(n_12620
		));
	notech_ao4 i_754(.A(n_950), .B(n_15049), .C(n_949), .D(n_15069), .Z(n_952
		));
	notech_reg_set dir2_reg_10(.CP(n_62957), .D(n_12626), .SD(n_62223), .Q(\dir2[10] 
		));
	notech_mux2 i_16790(.S(\nbus_14016[0] ), .A(\dir2[10] ), .B(n_52362), .Z
		(n_12626));
	notech_ao4 i_753(.A(n_950), .B(n_15048), .C(n_949), .D(n_15068), .Z(n_953
		));
	notech_reg_set dir2_reg_11(.CP(n_62957), .D(n_12632), .SD(n_62223), .Q(\dir2[11] 
		));
	notech_mux2 i_16798(.S(\nbus_14016[0] ), .A(\dir2[11] ), .B(n_52368), .Z
		(n_12632));
	notech_ao4 i_752(.A(n_950), .B(n_15047), .C(n_949), .D(n_15067), .Z(n_954
		));
	notech_reg_set dir2_reg_12(.CP(n_62957), .D(n_12638), .SD(n_62223), .Q(\dir2[12] 
		));
	notech_mux2 i_16806(.S(\nbus_14016[0] ), .A(\dir2[12] ), .B(n_52374), .Z
		(n_12638));
	notech_ao4 i_751(.A(n_950), .B(n_15046), .C(n_949), .D(n_15066), .Z(n_955
		));
	notech_reg_set dir2_reg_13(.CP(n_62956), .D(n_12644), .SD(n_62222), .Q(\dir2[13] 
		));
	notech_mux2 i_16814(.S(\nbus_14016[0] ), .A(\dir2[13] ), .B(n_52380), .Z
		(n_12644));
	notech_ao4 i_750(.A(n_950), .B(n_15045), .C(n_949), .D(n_15065), .Z(n_956
		));
	notech_reg_set dir2_reg_14(.CP(n_62956), .D(n_12650), .SD(n_62222), .Q(\dir2[14] 
		));
	notech_mux2 i_16822(.S(\nbus_14016[0] ), .A(\dir2[14] ), .B(n_52386), .Z
		(n_12650));
	notech_ao4 i_749(.A(n_950), .B(n_15044), .C(n_949), .D(n_15064), .Z(n_957
		));
	notech_reg_set dir2_reg_15(.CP(n_62956), .D(n_12656), .SD(n_62222), .Q(\dir2[15] 
		));
	notech_mux2 i_16830(.S(\nbus_14016[0] ), .A(\dir2[15] ), .B(n_52392), .Z
		(n_12656));
	notech_ao4 i_748(.A(n_950), .B(n_15043), .C(n_949), .D(n_15063), .Z(n_958
		));
	notech_reg_set dir2_reg_16(.CP(n_62957), .D(n_12662), .SD(n_62223), .Q(\dir2[16] 
		));
	notech_mux2 i_16838(.S(n_61263), .A(\dir2[16] ), .B(n_52398), .Z(n_12662
		));
	notech_ao4 i_747(.A(n_950), .B(n_15042), .C(n_949), .D(n_15062), .Z(n_959
		));
	notech_reg_set dir2_reg_17(.CP(n_62957), .D(n_12668), .SD(n_62223), .Q(\dir2[17] 
		));
	notech_mux2 i_16846(.S(n_61263), .A(\dir2[17] ), .B(n_52404), .Z(n_12668
		));
	notech_ao4 i_746(.A(n_950), .B(n_15041), .C(n_949), .D(n_15061), .Z(n_960
		));
	notech_reg_set dir2_reg_18(.CP(n_62957), .D(n_12674), .SD(n_62223), .Q(\dir2[18] 
		));
	notech_mux2 i_16854(.S(n_61263), .A(\dir2[18] ), .B(n_52410), .Z(n_12674
		));
	notech_ao4 i_745(.A(n_950), .B(n_15040), .C(n_949), .D(n_15060), .Z(n_961
		));
	notech_reg_set dir2_reg_19(.CP(n_62957), .D(n_12680), .SD(n_62223), .Q(\dir2[19] 
		));
	notech_mux2 i_16862(.S(n_61263), .A(\dir2[19] ), .B(n_52416), .Z(n_12680
		));
	notech_ao4 i_744(.A(n_950), .B(n_15039), .C(n_949), .D(n_15059), .Z(n_962
		));
	notech_reg_set dir2_reg_20(.CP(n_62957), .D(n_12686), .SD(n_62223), .Q(\dir2[20] 
		));
	notech_mux2 i_16870(.S(n_61263), .A(\dir2[20] ), .B(n_52422), .Z(n_12686
		));
	notech_ao4 i_743(.A(n_950), .B(n_15038), .C(n_949), .D(n_15058), .Z(n_963
		));
	notech_reg_set dir2_reg_21(.CP(n_62957), .D(n_12692), .SD(n_62223), .Q(\dir2[21] 
		));
	notech_mux2 i_16878(.S(n_61263), .A(\dir2[21] ), .B(n_52428), .Z(n_12692
		));
	notech_ao4 i_742(.A(n_950), .B(n_15037), .C(n_949), .D(n_15057), .Z(n_964
		));
	notech_reg_set dir2_reg_22(.CP(n_62957), .D(n_12698), .SD(n_62223), .Q(\dir2[22] 
		));
	notech_mux2 i_16886(.S(n_61263), .A(\dir2[22] ), .B(n_52434), .Z(n_12698
		));
	notech_ao4 i_741(.A(n_950), .B(n_15036), .C(n_949), .D(n_15056), .Z(n_965
		));
	notech_reg_set dir2_reg_23(.CP(n_62961), .D(n_12704), .SD(n_62227), .Q(\dir2[23] 
		));
	notech_mux2 i_16894(.S(n_61263), .A(\dir2[23] ), .B(n_52440), .Z(n_12704
		));
	notech_ao4 i_740(.A(n_950), .B(n_15035), .C(n_949), .D(n_15055), .Z(n_966
		));
	notech_reg_set dir2_reg_24(.CP(n_62965), .D(n_12710), .SD(n_62231), .Q(\dir2[24] 
		));
	notech_mux2 i_16902(.S(n_61263), .A(\dir2[24] ), .B(n_52446), .Z(n_12710
		));
	notech_ao4 i_739(.A(n_950), .B(n_15034), .C(n_949), .D(n_15054), .Z(n_967
		));
	notech_reg_set dir2_reg_25(.CP(n_62965), .D(n_12716), .SD(n_62231), .Q(\dir2[25] 
		));
	notech_mux2 i_16910(.S(n_61263), .A(\dir2[25] ), .B(n_52452), .Z(n_12716
		));
	notech_ao4 i_738(.A(n_950), .B(n_15033), .C(n_949), .D(n_15053), .Z(n_968
		));
	notech_reg_set dir2_reg_26(.CP(n_62965), .D(n_12722), .SD(n_62231), .Q(\dir2[26] 
		));
	notech_mux2 i_16918(.S(n_61263), .A(\dir2[26] ), .B(n_52458), .Z(n_12722
		));
	notech_ao4 i_737(.A(n_950), .B(n_15032), .C(n_949), .D(n_15052), .Z(n_969
		));
	notech_reg_set dir2_reg_27(.CP(n_62965), .D(n_12728), .SD(n_62231), .Q(\dir2[27] 
		));
	notech_mux2 i_16926(.S(n_61263), .A(\dir2[27] ), .B(n_52464), .Z(n_12728
		));
	notech_ao4 i_736(.A(n_950), .B(n_15031), .C(n_949), .D(n_15051), .Z(n_970
		));
	notech_reg_set dir2_reg_28(.CP(n_62965), .D(n_12734), .SD(n_62231), .Q(\dir2[28] 
		));
	notech_mux2 i_16934(.S(n_61263), .A(\dir2[28] ), .B(n_52470), .Z(n_12734
		));
	notech_reg_set dir2_reg_29(.CP(n_62965), .D(n_12740), .SD(n_62231), .Q(\dir2[29] 
		));
	notech_mux2 i_16942(.S(n_61263), .A(\dir2[29] ), .B(n_52476), .Z(n_12740
		));
	notech_ao3 i_031242(.A(n_62909), .B(n_15030), .C(n_62763), .Z(n_972));
	notech_reg_set dir2_reg_33(.CP(n_62965), .D(n_12746), .SD(n_62231), .Q(\dir2[33] 
		));
	notech_mux2 i_16950(.S(n_61263), .A(\dir2[33] ), .B(n_52501), .Z(n_12746
		));
	notech_and2 i_725(.A(n_62909), .B(n_883), .Z(n_973));
	notech_reg_set tab21_reg_0(.CP(n_62965), .D(n_12752), .SD(n_62231), .Q(\tab21[0] 
		));
	notech_mux2 i_16958(.S(\nbus_14019[0] ), .A(\tab21[0] ), .B(n_52574), .Z
		(n_12752));
	notech_nao3 i_9(.A(n_62909), .B(n_883), .C(n_62767), .Z(n_974));
	notech_reg_set tab21_reg_1(.CP(n_62966), .D(n_12758), .SD(n_62232), .Q(\tab21[1] 
		));
	notech_mux2 i_16966(.S(\nbus_14019[0] ), .A(\tab21[1] ), .B(n_52580), .Z
		(n_12758));
	notech_ao4 i_724(.A(n_974), .B(n_15229), .C(n_399), .D(n_15285), .Z(n_975
		));
	notech_reg_set tab21_reg_2(.CP(n_62966), .D(n_12764), .SD(n_62232), .Q(\tab21[2] 
		));
	notech_mux2 i_16974(.S(\nbus_14019[0] ), .A(\tab21[2] ), .B(n_52586), .Z
		(n_12764));
	notech_ao4 i_723(.A(n_974), .B(n_15230), .C(n_399), .D(n_15286), .Z(n_976
		));
	notech_reg_set tab21_reg_3(.CP(n_62965), .D(n_12770), .SD(n_62231), .Q(\tab21[3] 
		));
	notech_mux2 i_16982(.S(\nbus_14019[0] ), .A(\tab21[3] ), .B(n_52592), .Z
		(n_12770));
	notech_ao4 i_722(.A(n_974), .B(n_15231), .C(n_399), .D(n_15287), .Z(n_977
		));
	notech_reg tab21_reg_4(.CP(n_62965), .D(n_12776), .CD(n_62231), .Q(\tab21[4] 
		));
	notech_mux2 i_16990(.S(\nbus_14019[0] ), .A(\tab21[4] ), .B(n_873), .Z(n_12776
		));
	notech_ao4 i_721(.A(n_974), .B(n_15232), .C(n_399), .D(n_15288), .Z(n_978
		));
	notech_reg_set tab21_reg_5(.CP(n_62965), .D(n_12782), .SD(n_62231), .Q(\tab21[5] 
		));
	notech_mux2 i_16998(.S(\nbus_14019[0] ), .A(\tab21[5] ), .B(n_52604), .Z
		(n_12782));
	notech_ao4 i_720(.A(n_974), .B(n_15233), .C(n_399), .D(n_15289), .Z(n_979
		));
	notech_reg_set tab21_reg_6(.CP(n_62965), .D(n_12788), .SD(n_62231), .Q(\tab21[6] 
		));
	notech_mux2 i_17006(.S(\nbus_14019[0] ), .A(\tab21[6] ), .B(n_52610), .Z
		(n_12788));
	notech_ao4 i_719(.A(n_974), .B(n_15234), .C(n_399), .D(n_15290), .Z(n_980
		));
	notech_reg_set tab21_reg_7(.CP(n_62965), .D(n_12794), .SD(n_62231), .Q(\tab21[7] 
		));
	notech_mux2 i_17014(.S(\nbus_14019[0] ), .A(\tab21[7] ), .B(n_52616), .Z
		(n_12794));
	notech_ao4 i_718(.A(n_974), .B(n_15235), .C(n_399), .D(n_15291), .Z(n_981
		));
	notech_reg_set tab21_reg_8(.CP(n_62961), .D(n_12800), .SD(n_62227), .Q(\tab21[8] 
		));
	notech_mux2 i_17022(.S(\nbus_14019[0] ), .A(\tab21[8] ), .B(n_52622), .Z
		(n_12800));
	notech_ao4 i_717(.A(n_974), .B(n_15236), .C(n_399), .D(n_15292), .Z(n_982
		));
	notech_reg_set tab21_reg_9(.CP(n_62961), .D(n_12806), .SD(n_62227), .Q(\tab21[9] 
		));
	notech_mux2 i_17030(.S(\nbus_14019[0] ), .A(\tab21[9] ), .B(n_52628), .Z
		(n_12806));
	notech_ao4 i_716(.A(n_974), .B(n_15237), .C(n_399), .D(n_15293), .Z(n_983
		));
	notech_reg_set tab21_reg_10(.CP(n_62961), .D(n_12812), .SD(n_62227), .Q(\tab21[10] 
		));
	notech_mux2 i_17038(.S(\nbus_14019[0] ), .A(\tab21[10] ), .B(n_52634), .Z
		(n_12812));
	notech_ao4 i_715(.A(n_974), .B(n_15238), .C(n_399), .D(n_15294), .Z(n_984
		));
	notech_reg_set tab21_reg_11(.CP(n_62961), .D(n_12818), .SD(n_62227), .Q(\tab21[11] 
		));
	notech_mux2 i_17046(.S(\nbus_14019[0] ), .A(\tab21[11] ), .B(n_52640), .Z
		(n_12818));
	notech_nand2 i_63(.A(\hit_dir1[7] ), .B(n_972), .Z(n_985));
	notech_reg_set tab21_reg_12(.CP(n_62961), .D(n_12824), .SD(n_62227), .Q(\tab21[12] 
		));
	notech_mux2 i_17054(.S(\nbus_14019[0] ), .A(\tab21[12] ), .B(n_52646), .Z
		(n_12824));
	notech_ao3 i_713(.A(hit_tab13), .B(n_15339), .C(hit_tab11), .Z(n_986));
	notech_reg_set tab21_reg_13(.CP(n_62961), .D(n_12830), .SD(n_62227), .Q(\tab21[13] 
		));
	notech_mux2 i_17062(.S(\nbus_14019[0] ), .A(\tab21[13] ), .B(n_52652), .Z
		(n_12830));
	notech_reg_set tab21_reg_14(.CP(n_62961), .D(n_12836), .SD(n_62227), .Q(\tab21[14] 
		));
	notech_mux2 i_17070(.S(\nbus_14019[0] ), .A(\tab21[14] ), .B(n_52658), .Z
		(n_12836));
	notech_or4 i_25(.A(hit_tab12), .B(hit_tab11), .C(hit_tab13), .D(n_985), 
		.Z(n_988));
	notech_reg_set tab21_reg_15(.CP(n_62965), .D(n_12842), .SD(n_62231), .Q(\tab21[15] 
		));
	notech_mux2 i_17078(.S(\nbus_14019[0] ), .A(\tab21[15] ), .B(n_52664), .Z
		(n_12842));
	notech_reg_set tab21_reg_16(.CP(n_62965), .D(n_12848), .SD(n_62231), .Q(\tab21[16] 
		));
	notech_mux2 i_17086(.S(n_61241), .A(\tab21[16] ), .B(n_52670), .Z(n_12848
		));
	notech_nao3 i_24(.A(hit_tab12), .B(n_62745), .C(hit_tab11), .Z(n_990));
	notech_reg_set tab21_reg_17(.CP(n_62965), .D(n_12854), .SD(n_62231), .Q(\tab21[17] 
		));
	notech_mux2 i_17094(.S(n_61241), .A(\tab21[17] ), .B(n_52676), .Z(n_12854
		));
	notech_ao4 i_708(.A(n_15146), .B(n_990), .C(n_988), .D(n_15167), .Z(n_991
		));
	notech_reg_set tab21_reg_18(.CP(n_62965), .D(n_12860), .SD(n_62231), .Q(\tab21[18] 
		));
	notech_mux2 i_17102(.S(n_61241), .A(\tab21[18] ), .B(n_52682), .Z(n_12860
		));
	notech_reg_set tab21_reg_19(.CP(n_62961), .D(n_12866), .SD(n_62227), .Q(\tab21[19] 
		));
	notech_mux2 i_17110(.S(n_61241), .A(\tab21[19] ), .B(n_52688), .Z(n_12866
		));
	notech_or4 i_62(.A(n_62767), .B(\hit_dir1[7] ), .C(n_15341), .D(n_883), 
		.Z(n_993));
	notech_reg_set tab21_reg_20(.CP(n_62961), .D(n_12872), .SD(n_62227), .Q(\tab21[20] 
		));
	notech_mux2 i_17118(.S(n_61241), .A(\tab21[20] ), .B(n_52694), .Z(n_12872
		));
	notech_and2 i_711(.A(hit_tab22), .B(n_15337), .Z(n_994));
	notech_reg_set tab21_reg_21(.CP(n_62965), .D(n_12878), .SD(n_62231), .Q(\tab21[21] 
		));
	notech_mux2 i_17126(.S(n_61241), .A(\tab21[21] ), .B(n_52700), .Z(n_12878
		));
	notech_reg_set tab21_reg_22(.CP(n_62976), .D(n_12884), .SD(n_62242), .Q(\tab21[22] 
		));
	notech_mux2 i_17134(.S(n_61241), .A(\tab21[22] ), .B(n_52706), .Z(n_12884
		));
	notech_nand2 i_22(.A(hit_tab11), .B(n_62745), .Z(n_996));
	notech_reg_set tab21_reg_23(.CP(n_62989), .D(n_12890), .SD(n_62255), .Q(\tab21[23] 
		));
	notech_mux2 i_17142(.S(n_61241), .A(\tab21[23] ), .B(n_52712), .Z(n_12890
		));
	notech_reg_set tab21_reg_24(.CP(n_62989), .D(n_12896), .SD(n_62255), .Q(\tab21[24] 
		));
	notech_mux2 i_17150(.S(n_61241), .A(\tab21[24] ), .B(n_52718), .Z(n_12896
		));
	notech_or4 i_16(.A(hit_tab22), .B(hit_tab21), .C(n_62754), .D(n_15338), 
		.Z(n_998));
	notech_reg_set tab21_reg_25(.CP(n_62989), .D(n_12902), .SD(n_62255), .Q(\tab21[25] 
		));
	notech_mux2 i_17158(.S(n_61241), .A(\tab21[25] ), .B(n_52724), .Z(n_12902
		));
	notech_ao4 i_706(.A(n_998), .B(n_15093), .C(n_996), .D(n_15196), .Z(n_999
		));
	notech_reg_set tab21_reg_26(.CP(n_62989), .D(n_12908), .SD(n_62255), .Q(\tab21[26] 
		));
	notech_mux2 i_17166(.S(n_61241), .A(\tab21[26] ), .B(n_52730), .Z(n_12908
		));
	notech_reg_set tab21_reg_27(.CP(n_62989), .D(n_12914), .SD(n_62255), .Q(\tab21[27] 
		));
	notech_mux2 i_17174(.S(n_61241), .A(\tab21[27] ), .B(n_52736), .Z(n_12914
		));
	notech_and4 i_710(.A(n_999), .B(n_991), .C(n_776), .D(n_779), .Z(n_1001)
		);
	notech_reg_set tab21_reg_28(.CP(n_62989), .D(n_12920), .SD(n_62255), .Q(\tab21[28] 
		));
	notech_mux2 i_17182(.S(n_61241), .A(\tab21[28] ), .B(n_52742), .Z(n_12920
		));
	notech_nao3 i_13(.A(hit_tab21), .B(n_972), .C(\hit_dir1[7] ), .Z(n_1002)
		);
	notech_reg_set tab21_reg_29(.CP(n_62989), .D(n_12926), .SD(n_62255), .Q(\tab21[29] 
		));
	notech_mux2 i_17190(.S(n_61241), .A(\tab21[29] ), .B(n_52748), .Z(n_12926
		));
	notech_or4 i_12(.A(hit_tab22), .B(hit_tab21), .C(hit_tab23), .D(n_62754)
		, .Z(n_1003));
	notech_reg_set tab21_reg_33(.CP(n_62993), .D(n_12932), .SD(n_62259), .Q(\tab21[33] 
		));
	notech_mux2 i_17198(.S(n_61241), .A(\tab21[33] ), .B(n_52772), .Z(n_12932
		));
	notech_ao4 i_703(.A(n_1003), .B(n_15117), .C(n_1002), .D(n_15072), .Z(n_1004
		));
	notech_reg hit_adr21_reg(.CP(n_62993), .D(n_12938), .CD(n_62259), .Q(hit_adr21
		));
	notech_mux2 i_17206(.S(n_872), .A(hit_add21), .B(hit_adr21), .Z(n_12938)
		);
	notech_reg_set tab22_reg_0(.CP(n_62993), .D(n_12944), .SD(n_62259), .Q(\tab22[0] 
		));
	notech_mux2 i_17214(.S(\nbus_14023[0] ), .A(\tab22[0] ), .B(n_52574), .Z
		(n_12944));
	notech_ao4 i_702(.A(n_62904), .B(n_15295), .C(n_878), .D(n_15239), .Z(n_1006
		));
	notech_reg_set tab22_reg_1(.CP(n_62993), .D(n_12950), .SD(n_62259), .Q(\tab22[1] 
		));
	notech_mux2 i_17222(.S(\nbus_14023[0] ), .A(\tab22[1] ), .B(n_52580), .Z
		(n_12950));
	notech_reg_set tab22_reg_2(.CP(n_62989), .D(n_12956), .SD(n_62255), .Q(\tab22[2] 
		));
	notech_mux2 i_17230(.S(\nbus_14023[0] ), .A(\tab22[2] ), .B(n_52586), .Z
		(n_12956));
	notech_ao4 i_699(.A(n_990), .B(n_15147), .C(n_988), .D(n_15168), .Z(n_1008
		));
	notech_reg_set tab22_reg_3(.CP(n_62993), .D(n_12962), .SD(n_62259), .Q(\tab22[3] 
		));
	notech_mux2 i_17238(.S(\nbus_14023[0] ), .A(\tab22[3] ), .B(n_52592), .Z
		(n_12962));
	notech_reg tab22_reg_4(.CP(n_62993), .D(n_12968), .CD(n_62259), .Q(\tab22[4] 
		));
	notech_mux2 i_17246(.S(\nbus_14023[0] ), .A(\tab22[4] ), .B(n_873), .Z(n_12968
		));
	notech_ao4 i_697(.A(n_998), .B(n_15094), .C(n_996), .D(n_15197), .Z(n_1010
		));
	notech_reg_set tab22_reg_5(.CP(n_62989), .D(n_12974), .SD(n_62255), .Q(\tab22[5] 
		));
	notech_mux2 i_17254(.S(\nbus_14023[0] ), .A(\tab22[5] ), .B(n_52604), .Z
		(n_12974));
	notech_reg_set tab22_reg_6(.CP(n_62985), .D(n_12980), .SD(n_62251), .Q(\tab22[6] 
		));
	notech_mux2 i_17262(.S(\nbus_14023[0] ), .A(\tab22[6] ), .B(n_52610), .Z
		(n_12980));
	notech_and4 i_701(.A(n_1010), .B(n_1008), .C(n_765), .D(n_768), .Z(n_1012
		));
	notech_reg_set tab22_reg_7(.CP(n_62989), .D(n_12986), .SD(n_62255), .Q(\tab22[7] 
		));
	notech_mux2 i_17270(.S(\nbus_14023[0] ), .A(\tab22[7] ), .B(n_52616), .Z
		(n_12986));
	notech_ao4 i_694(.A(n_1003), .B(n_15118), .C(n_1002), .D(n_15073), .Z(n_1013
		));
	notech_reg_set tab22_reg_8(.CP(n_62989), .D(n_12992), .SD(n_62255), .Q(\tab22[8] 
		));
	notech_mux2 i_17278(.S(\nbus_14023[0] ), .A(\tab22[8] ), .B(n_52622), .Z
		(n_12992));
	notech_reg_set tab22_reg_9(.CP(n_62985), .D(n_12998), .SD(n_62251), .Q(\tab22[9] 
		));
	notech_mux2 i_17286(.S(\nbus_14023[0] ), .A(\tab22[9] ), .B(n_52628), .Z
		(n_12998));
	notech_ao4 i_693(.A(n_62904), .B(n_15296), .C(n_878), .D(n_15240), .Z(n_1015
		));
	notech_reg_set tab22_reg_10(.CP(n_62985), .D(n_13004), .SD(n_62251), .Q(\tab22[10] 
		));
	notech_mux2 i_17294(.S(\nbus_14023[0] ), .A(\tab22[10] ), .B(n_52634), .Z
		(n_13004));
	notech_reg_set tab22_reg_11(.CP(n_62985), .D(n_13010), .SD(n_62251), .Q(\tab22[11] 
		));
	notech_mux2 i_17302(.S(\nbus_14023[0] ), .A(\tab22[11] ), .B(n_52640), .Z
		(n_13010));
	notech_ao4 i_690(.A(n_990), .B(n_15148), .C(n_988), .D(n_15169), .Z(n_1017
		));
	notech_reg_set tab22_reg_12(.CP(n_62985), .D(n_13016), .SD(n_62251), .Q(\tab22[12] 
		));
	notech_mux2 i_17310(.S(\nbus_14023[0] ), .A(\tab22[12] ), .B(n_52646), .Z
		(n_13016));
	notech_reg_set tab22_reg_13(.CP(n_62989), .D(n_13022), .SD(n_62255), .Q(\tab22[13] 
		));
	notech_mux2 i_17318(.S(\nbus_14023[0] ), .A(\tab22[13] ), .B(n_52652), .Z
		(n_13022));
	notech_ao4 i_688(.A(n_998), .B(n_15095), .C(n_996), .D(n_15198), .Z(n_1019
		));
	notech_reg_set tab22_reg_14(.CP(n_62989), .D(n_13028), .SD(n_62255), .Q(\tab22[14] 
		));
	notech_mux2 i_17326(.S(\nbus_14023[0] ), .A(\tab22[14] ), .B(n_52658), .Z
		(n_13028));
	notech_reg_set tab22_reg_15(.CP(n_62989), .D(n_13034), .SD(n_62255), .Q(\tab22[15] 
		));
	notech_mux2 i_17334(.S(\nbus_14023[0] ), .A(\tab22[15] ), .B(n_52664), .Z
		(n_13034));
	notech_and4 i_692(.A(n_1019), .B(n_1017), .C(n_754), .D(n_757), .Z(n_1021
		));
	notech_reg_set tab22_reg_16(.CP(n_62989), .D(n_13040), .SD(n_62255), .Q(\tab22[16] 
		));
	notech_mux2 i_17342(.S(n_61252), .A(\tab22[16] ), .B(n_52670), .Z(n_13040
		));
	notech_ao4 i_685(.A(n_1003), .B(n_15119), .C(n_1002), .D(n_15074), .Z(n_1022
		));
	notech_reg_set tab22_reg_17(.CP(n_62989), .D(n_13046), .SD(n_62255), .Q(\tab22[17] 
		));
	notech_mux2 i_17350(.S(n_61252), .A(\tab22[17] ), .B(n_52676), .Z(n_13046
		));
	notech_reg_set tab22_reg_18(.CP(n_62989), .D(n_13052), .SD(n_62255), .Q(\tab22[18] 
		));
	notech_mux2 i_17358(.S(n_61252), .A(\tab22[18] ), .B(n_52682), .Z(n_13052
		));
	notech_ao4 i_684(.A(n_62904), .B(n_15297), .C(n_878), .D(n_15241), .Z(n_1024
		));
	notech_reg_set tab22_reg_19(.CP(n_62989), .D(n_13058), .SD(n_62255), .Q(\tab22[19] 
		));
	notech_mux2 i_17366(.S(n_61252), .A(\tab22[19] ), .B(n_52688), .Z(n_13058
		));
	notech_reg_set tab22_reg_20(.CP(n_62993), .D(n_13064), .SD(n_62259), .Q(\tab22[20] 
		));
	notech_mux2 i_17374(.S(n_61252), .A(\tab22[20] ), .B(n_52694), .Z(n_13064
		));
	notech_ao4 i_681(.A(n_990), .B(n_15149), .C(n_988), .D(n_15170), .Z(n_1026
		));
	notech_reg_set tab22_reg_21(.CP(n_62994), .D(n_13070), .SD(n_62260), .Q(\tab22[21] 
		));
	notech_mux2 i_17382(.S(n_61252), .A(\tab22[21] ), .B(n_52700), .Z(n_13070
		));
	notech_reg_set tab22_reg_22(.CP(n_62994), .D(n_13076), .SD(n_62260), .Q(\tab22[22] 
		));
	notech_mux2 i_17390(.S(n_61252), .A(\tab22[22] ), .B(n_52706), .Z(n_13076
		));
	notech_ao4 i_679(.A(n_998), .B(n_15096), .C(n_996), .D(n_15199), .Z(n_1028
		));
	notech_reg_set tab22_reg_23(.CP(n_62994), .D(n_13082), .SD(n_62260), .Q(\tab22[23] 
		));
	notech_mux2 i_17398(.S(n_61252), .A(\tab22[23] ), .B(n_52712), .Z(n_13082
		));
	notech_reg_set tab22_reg_24(.CP(n_62994), .D(n_13088), .SD(n_62260), .Q(\tab22[24] 
		));
	notech_mux2 i_17406(.S(n_61252), .A(\tab22[24] ), .B(n_52718), .Z(n_13088
		));
	notech_and4 i_683(.A(n_1028), .B(n_1026), .C(n_743), .D(n_746), .Z(n_1030
		));
	notech_reg_set tab22_reg_25(.CP(n_62994), .D(n_13094), .SD(n_62260), .Q(\tab22[25] 
		));
	notech_mux2 i_17414(.S(n_61252), .A(\tab22[25] ), .B(n_52724), .Z(n_13094
		));
	notech_ao4 i_676(.A(n_1003), .B(n_15120), .C(n_1002), .D(n_15075), .Z(n_1031
		));
	notech_reg_set tab22_reg_26(.CP(n_62994), .D(n_13100), .SD(n_62260), .Q(\tab22[26] 
		));
	notech_mux2 i_17422(.S(n_61252), .A(\tab22[26] ), .B(n_52730), .Z(n_13100
		));
	notech_reg_set tab22_reg_27(.CP(n_62994), .D(n_13106), .SD(n_62260), .Q(\tab22[27] 
		));
	notech_mux2 i_17430(.S(n_61252), .A(\tab22[27] ), .B(n_52736), .Z(n_13106
		));
	notech_ao4 i_675(.A(n_62904), .B(n_15298), .C(n_878), .D(n_15242), .Z(n_1033
		));
	notech_reg_set tab22_reg_28(.CP(n_62994), .D(n_13112), .SD(n_62260), .Q(\tab22[28] 
		));
	notech_mux2 i_17438(.S(n_61252), .A(\tab22[28] ), .B(n_52742), .Z(n_13112
		));
	notech_reg_set tab22_reg_29(.CP(n_62994), .D(n_13118), .SD(n_62260), .Q(\tab22[29] 
		));
	notech_mux2 i_17446(.S(n_61252), .A(\tab22[29] ), .B(n_52748), .Z(n_13118
		));
	notech_ao4 i_672(.A(n_990), .B(n_15150), .C(n_988), .D(n_15171), .Z(n_1035
		));
	notech_reg_set tab22_reg_33(.CP(n_62994), .D(n_13124), .SD(n_62260), .Q(\tab22[33] 
		));
	notech_mux2 i_17454(.S(n_61252), .A(\tab22[33] ), .B(n_52772), .Z(n_13124
		));
	notech_reg hit_adr22_reg(.CP(n_62994), .D(n_13130), .CD(n_62260), .Q(hit_adr22
		));
	notech_mux2 i_17462(.S(n_872), .A(hit_add22), .B(hit_adr22), .Z(n_13130)
		);
	notech_ao4 i_670(.A(n_998), .B(n_15097), .C(n_996), .D(n_15200), .Z(n_1037
		));
	notech_reg_set tab23_reg_0(.CP(n_62994), .D(n_13136), .SD(n_62260), .Q(\tab23[0] 
		));
	notech_mux2 i_17470(.S(\nbus_14025[0] ), .A(\tab23[0] ), .B(n_52574), .Z
		(n_13136));
	notech_reg_set tab23_reg_1(.CP(n_62994), .D(n_13142), .SD(n_62260), .Q(\tab23[1] 
		));
	notech_mux2 i_17478(.S(\nbus_14025[0] ), .A(\tab23[1] ), .B(n_52580), .Z
		(n_13142));
	notech_and4 i_674(.A(n_1037), .B(n_1035), .C(n_732), .D(n_735), .Z(n_1039
		));
	notech_reg_set tab23_reg_2(.CP(n_62994), .D(n_13148), .SD(n_62260), .Q(\tab23[2] 
		));
	notech_mux2 i_17486(.S(\nbus_14025[0] ), .A(\tab23[2] ), .B(n_52586), .Z
		(n_13148));
	notech_ao4 i_667(.A(n_1003), .B(n_15121), .C(n_1002), .D(n_15076), .Z(n_1040
		));
	notech_reg_set tab23_reg_3(.CP(n_62994), .D(n_13154), .SD(n_62260), .Q(\tab23[3] 
		));
	notech_mux2 i_17494(.S(\nbus_14025[0] ), .A(\tab23[3] ), .B(n_52592), .Z
		(n_13154));
	notech_reg tab23_reg_4(.CP(n_62993), .D(n_13160), .CD(n_62259), .Q(\tab23[4] 
		));
	notech_mux2 i_17502(.S(\nbus_14025[0] ), .A(\tab23[4] ), .B(n_873), .Z(n_13160
		));
	notech_ao4 i_666(.A(n_62904), .B(n_15299), .C(n_878), .D(n_15243), .Z(n_1042
		));
	notech_reg_set tab23_reg_5(.CP(n_62993), .D(n_13166), .SD(n_62259), .Q(\tab23[5] 
		));
	notech_mux2 i_17510(.S(\nbus_14025[0] ), .A(\tab23[5] ), .B(n_52604), .Z
		(n_13166));
	notech_reg_set tab23_reg_6(.CP(n_62993), .D(n_13172), .SD(n_62259), .Q(\tab23[6] 
		));
	notech_mux2 i_17518(.S(\nbus_14025[0] ), .A(\tab23[6] ), .B(n_52610), .Z
		(n_13172));
	notech_ao4 i_663(.A(n_990), .B(n_15151), .C(n_988), .D(n_15172), .Z(n_1044
		));
	notech_reg_set tab23_reg_7(.CP(n_62993), .D(n_13178), .SD(n_62259), .Q(\tab23[7] 
		));
	notech_mux2 i_17526(.S(\nbus_14025[0] ), .A(\tab23[7] ), .B(n_52616), .Z
		(n_13178));
	notech_reg_set tab23_reg_8(.CP(n_62993), .D(n_13184), .SD(n_62259), .Q(\tab23[8] 
		));
	notech_mux2 i_17534(.S(\nbus_14025[0] ), .A(\tab23[8] ), .B(n_52622), .Z
		(n_13184));
	notech_ao4 i_661(.A(n_998), .B(n_15098), .C(n_996), .D(n_15201), .Z(n_1046
		));
	notech_reg_set tab23_reg_9(.CP(n_62993), .D(n_13190), .SD(n_62259), .Q(\tab23[9] 
		));
	notech_mux2 i_17542(.S(\nbus_14025[0] ), .A(\tab23[9] ), .B(n_52628), .Z
		(n_13190));
	notech_reg_set tab23_reg_10(.CP(n_62993), .D(n_13196), .SD(n_62259), .Q(\tab23[10] 
		));
	notech_mux2 i_17550(.S(\nbus_14025[0] ), .A(\tab23[10] ), .B(n_52634), .Z
		(n_13196));
	notech_and4 i_665(.A(n_1046), .B(n_1044), .C(n_721), .D(n_724), .Z(n_1048
		));
	notech_reg_set tab23_reg_11(.CP(n_62994), .D(n_13202), .SD(n_62260), .Q(\tab23[11] 
		));
	notech_mux2 i_17558(.S(\nbus_14025[0] ), .A(\tab23[11] ), .B(n_52640), .Z
		(n_13202));
	notech_ao4 i_658(.A(n_1003), .B(n_15122), .C(n_1002), .D(n_15077), .Z(n_1049
		));
	notech_reg_set tab23_reg_12(.CP(n_62994), .D(n_13208), .SD(n_62260), .Q(\tab23[12] 
		));
	notech_mux2 i_17566(.S(\nbus_14025[0] ), .A(\tab23[12] ), .B(n_52646), .Z
		(n_13208));
	notech_reg_set tab23_reg_13(.CP(n_62994), .D(n_13214), .SD(n_62260), .Q(\tab23[13] 
		));
	notech_mux2 i_17574(.S(\nbus_14025[0] ), .A(\tab23[13] ), .B(n_52652), .Z
		(n_13214));
	notech_ao4 i_657(.A(n_62904), .B(n_15300), .C(n_878), .D(n_15244), .Z(n_1051
		));
	notech_reg_set tab23_reg_14(.CP(n_62993), .D(n_13220), .SD(n_62259), .Q(\tab23[14] 
		));
	notech_mux2 i_17582(.S(\nbus_14025[0] ), .A(\tab23[14] ), .B(n_52658), .Z
		(n_13220));
	notech_reg_set tab23_reg_15(.CP(n_62993), .D(n_13226), .SD(n_62259), .Q(\tab23[15] 
		));
	notech_mux2 i_17590(.S(\nbus_14025[0] ), .A(\tab23[15] ), .B(n_52664), .Z
		(n_13226));
	notech_ao4 i_654(.A(n_990), .B(n_15152), .C(n_988), .D(n_15173), .Z(n_1053
		));
	notech_reg_set tab23_reg_16(.CP(n_62993), .D(n_13232), .SD(n_62259), .Q(\tab23[16] 
		));
	notech_mux2 i_17598(.S(n_61219), .A(\tab23[16] ), .B(n_52670), .Z(n_13232
		));
	notech_reg_set tab23_reg_17(.CP(n_62993), .D(n_13238), .SD(n_62259), .Q(\tab23[17] 
		));
	notech_mux2 i_17606(.S(n_61219), .A(\tab23[17] ), .B(n_52676), .Z(n_13238
		));
	notech_ao4 i_652(.A(n_998), .B(n_15099), .C(n_996), .D(n_15202), .Z(n_1055
		));
	notech_reg_set tab23_reg_18(.CP(n_62980), .D(n_13244), .SD(n_62246), .Q(\tab23[18] 
		));
	notech_mux2 i_17614(.S(n_61219), .A(\tab23[18] ), .B(n_52682), .Z(n_13244
		));
	notech_reg_set tab23_reg_19(.CP(n_62980), .D(n_13250), .SD(n_62246), .Q(\tab23[19] 
		));
	notech_mux2 i_17622(.S(n_61219), .A(\tab23[19] ), .B(n_52688), .Z(n_13250
		));
	notech_and4 i_656(.A(n_1055), .B(n_1053), .C(n_710), .D(n_713), .Z(n_1057
		));
	notech_reg_set tab23_reg_20(.CP(n_62980), .D(n_13256), .SD(n_62246), .Q(\tab23[20] 
		));
	notech_mux2 i_17630(.S(n_61219), .A(\tab23[20] ), .B(n_52694), .Z(n_13256
		));
	notech_ao4 i_649(.A(n_1003), .B(n_15123), .C(n_1002), .D(n_15078), .Z(n_1058
		));
	notech_reg_set tab23_reg_21(.CP(n_62980), .D(n_13262), .SD(n_62246), .Q(\tab23[21] 
		));
	notech_mux2 i_17638(.S(n_61219), .A(\tab23[21] ), .B(n_52700), .Z(n_13262
		));
	notech_reg_set tab23_reg_22(.CP(n_62980), .D(n_13268), .SD(n_62246), .Q(\tab23[22] 
		));
	notech_mux2 i_17646(.S(n_61219), .A(\tab23[22] ), .B(n_52706), .Z(n_13268
		));
	notech_ao4 i_648(.A(n_62904), .B(n_15301), .C(n_878), .D(n_15245), .Z(n_1060
		));
	notech_reg_set tab23_reg_23(.CP(n_62980), .D(n_13274), .SD(n_62246), .Q(\tab23[23] 
		));
	notech_mux2 i_17654(.S(n_61219), .A(\tab23[23] ), .B(n_52712), .Z(n_13274
		));
	notech_reg_set tab23_reg_24(.CP(n_62980), .D(n_13280), .SD(n_62246), .Q(\tab23[24] 
		));
	notech_mux2 i_17662(.S(n_61219), .A(\tab23[24] ), .B(n_52718), .Z(n_13280
		));
	notech_ao4 i_645(.A(n_990), .B(n_15153), .C(n_988), .D(n_15174), .Z(n_1062
		));
	notech_reg_set tab23_reg_25(.CP(n_62980), .D(n_13286), .SD(n_62246), .Q(\tab23[25] 
		));
	notech_mux2 i_17670(.S(n_61219), .A(\tab23[25] ), .B(n_52724), .Z(n_13286
		));
	notech_reg_set tab23_reg_26(.CP(n_62980), .D(n_13292), .SD(n_62246), .Q(\tab23[26] 
		));
	notech_mux2 i_17678(.S(n_61219), .A(\tab23[26] ), .B(n_52730), .Z(n_13292
		));
	notech_ao4 i_643(.A(n_998), .B(n_15101), .C(n_996), .D(n_15203), .Z(n_1064
		));
	notech_reg_set tab23_reg_27(.CP(n_62984), .D(n_13298), .SD(n_62250), .Q(\tab23[27] 
		));
	notech_mux2 i_17686(.S(n_61219), .A(\tab23[27] ), .B(n_52736), .Z(n_13298
		));
	notech_reg_set tab23_reg_28(.CP(n_62980), .D(n_13304), .SD(n_62246), .Q(\tab23[28] 
		));
	notech_mux2 i_17694(.S(n_61219), .A(\tab23[28] ), .B(n_52742), .Z(n_13304
		));
	notech_and4 i_647(.A(n_1064), .B(n_1062), .C(n_699), .D(n_702), .Z(n_1066
		));
	notech_reg_set tab23_reg_29(.CP(n_62980), .D(n_13310), .SD(n_62246), .Q(\tab23[29] 
		));
	notech_mux2 i_17702(.S(n_61219), .A(\tab23[29] ), .B(n_52748), .Z(n_13310
		));
	notech_ao4 i_640(.A(n_1003), .B(n_15124), .C(n_1002), .D(n_15079), .Z(n_1067
		));
	notech_reg_set tab23_reg_33(.CP(n_62980), .D(n_13316), .SD(n_62246), .Q(\tab23[33] 
		));
	notech_mux2 i_17710(.S(n_61219), .A(\tab23[33] ), .B(n_52772), .Z(n_13316
		));
	notech_reg hit_adr23_reg(.CP(n_62980), .D(n_13322), .CD(n_62246), .Q(hit_adr23
		));
	notech_mux2 i_17718(.S(n_872), .A(hit_add23), .B(hit_adr23), .Z(n_13322)
		);
	notech_ao4 i_639(.A(n_62904), .B(n_15302), .C(n_878), .D(n_15246), .Z(n_1069
		));
	notech_reg_set tab24_reg_0(.CP(n_62980), .D(n_13328), .SD(n_62246), .Q(\tab24[0] 
		));
	notech_mux2 i_17726(.S(\nbus_14039[0] ), .A(\tab24[0] ), .B(n_52574), .Z
		(n_13328));
	notech_reg_set tab24_reg_1(.CP(n_62976), .D(n_13334), .SD(n_62242), .Q(\tab24[1] 
		));
	notech_mux2 i_17734(.S(\nbus_14039[0] ), .A(\tab24[1] ), .B(n_52580), .Z
		(n_13334));
	notech_ao4 i_636(.A(n_990), .B(n_15154), .C(n_988), .D(n_15175), .Z(n_1071
		));
	notech_reg_set tab24_reg_2(.CP(n_62976), .D(n_13340), .SD(n_62242), .Q(\tab24[2] 
		));
	notech_mux2 i_17742(.S(\nbus_14039[0] ), .A(\tab24[2] ), .B(n_52586), .Z
		(n_13340));
	notech_reg_set tab24_reg_3(.CP(n_62976), .D(n_13346), .SD(n_62242), .Q(\tab24[3] 
		));
	notech_mux2 i_17750(.S(\nbus_14039[0] ), .A(\tab24[3] ), .B(n_52592), .Z
		(n_13346));
	notech_ao4 i_634(.A(n_998), .B(n_15102), .C(n_996), .D(n_15204), .Z(n_1073
		));
	notech_reg tab24_reg_4(.CP(n_62976), .D(n_13352), .CD(n_62242), .Q(\tab24[4] 
		));
	notech_mux2 i_17758(.S(\nbus_14039[0] ), .A(\tab24[4] ), .B(n_873), .Z(n_13352
		));
	notech_reg_set tab24_reg_5(.CP(n_62976), .D(n_13358), .SD(n_62242), .Q(\tab24[5] 
		));
	notech_mux2 i_17766(.S(\nbus_14039[0] ), .A(\tab24[5] ), .B(n_52604), .Z
		(n_13358));
	notech_and4 i_638(.A(n_1073), .B(n_1071), .C(n_688), .D(n_691), .Z(n_1075
		));
	notech_reg_set tab24_reg_6(.CP(n_62976), .D(n_13364), .SD(n_62242), .Q(\tab24[6] 
		));
	notech_mux2 i_17774(.S(\nbus_14039[0] ), .A(\tab24[6] ), .B(n_52610), .Z
		(n_13364));
	notech_ao4 i_631(.A(n_1003), .B(n_15125), .C(n_1002), .D(n_15080), .Z(n_1076
		));
	notech_reg_set tab24_reg_7(.CP(n_62976), .D(n_13370), .SD(n_62242), .Q(\tab24[7] 
		));
	notech_mux2 i_17782(.S(\nbus_14039[0] ), .A(\tab24[7] ), .B(n_52616), .Z
		(n_13370));
	notech_reg_set tab24_reg_8(.CP(n_62980), .D(n_13376), .SD(n_62246), .Q(\tab24[8] 
		));
	notech_mux2 i_17790(.S(\nbus_14039[0] ), .A(\tab24[8] ), .B(n_52622), .Z
		(n_13376));
	notech_ao4 i_630(.A(n_62904), .B(n_15303), .C(n_878), .D(n_15247), .Z(n_1078
		));
	notech_reg_set tab24_reg_9(.CP(n_62980), .D(n_13382), .SD(n_62246), .Q(\tab24[9] 
		));
	notech_mux2 i_17798(.S(\nbus_14039[0] ), .A(\tab24[9] ), .B(n_52628), .Z
		(n_13382));
	notech_reg_set tab24_reg_10(.CP(n_62980), .D(n_13388), .SD(n_62246), .Q(\tab24[10] 
		));
	notech_mux2 i_17806(.S(\nbus_14039[0] ), .A(\tab24[10] ), .B(n_52634), .Z
		(n_13388));
	notech_ao4 i_627(.A(n_990), .B(n_15155), .C(n_988), .D(n_15176), .Z(n_1080
		));
	notech_reg_set tab24_reg_11(.CP(n_62980), .D(n_13394), .SD(n_62246), .Q(\tab24[11] 
		));
	notech_mux2 i_17814(.S(\nbus_14039[0] ), .A(\tab24[11] ), .B(n_52640), .Z
		(n_13394));
	notech_reg_set tab24_reg_12(.CP(n_62976), .D(n_13400), .SD(n_62242), .Q(\tab24[12] 
		));
	notech_mux2 i_17822(.S(\nbus_14039[0] ), .A(\tab24[12] ), .B(n_52646), .Z
		(n_13400));
	notech_ao4 i_625(.A(n_998), .B(n_15103), .C(n_996), .D(n_15205), .Z(n_1082
		));
	notech_reg_set tab24_reg_13(.CP(n_62976), .D(n_13406), .SD(n_62242), .Q(\tab24[13] 
		));
	notech_mux2 i_17830(.S(\nbus_14039[0] ), .A(\tab24[13] ), .B(n_52652), .Z
		(n_13406));
	notech_reg_set tab24_reg_14(.CP(n_62976), .D(n_13412), .SD(n_62242), .Q(\tab24[14] 
		));
	notech_mux2 i_17838(.S(\nbus_14039[0] ), .A(\tab24[14] ), .B(n_52658), .Z
		(n_13412));
	notech_and4 i_629(.A(n_1082), .B(n_1080), .C(n_677), .D(n_680), .Z(n_1084
		));
	notech_reg_set tab24_reg_15(.CP(n_62984), .D(n_13418), .SD(n_62250), .Q(\tab24[15] 
		));
	notech_mux2 i_17846(.S(\nbus_14039[0] ), .A(\tab24[15] ), .B(n_52664), .Z
		(n_13418));
	notech_ao4 i_622(.A(n_1003), .B(n_15126), .C(n_1002), .D(n_15081), .Z(n_1085
		));
	notech_reg_set tab24_reg_16(.CP(n_62985), .D(n_13424), .SD(n_62251), .Q(\tab24[16] 
		));
	notech_mux2 i_17854(.S(n_61230), .A(\tab24[16] ), .B(n_52670), .Z(n_13424
		));
	notech_reg_set tab24_reg_17(.CP(n_62985), .D(n_13430), .SD(n_62251), .Q(\tab24[17] 
		));
	notech_mux2 i_17862(.S(n_61230), .A(\tab24[17] ), .B(n_52676), .Z(n_13430
		));
	notech_ao4 i_621(.A(n_62904), .B(n_15304), .C(n_878), .D(n_15248), .Z(n_1087
		));
	notech_reg_set tab24_reg_18(.CP(n_62985), .D(n_13436), .SD(n_62251), .Q(\tab24[18] 
		));
	notech_mux2 i_17870(.S(n_61230), .A(\tab24[18] ), .B(n_52682), .Z(n_13436
		));
	notech_reg_set tab24_reg_19(.CP(n_62985), .D(n_13442), .SD(n_62251), .Q(\tab24[19] 
		));
	notech_mux2 i_17878(.S(n_61230), .A(\tab24[19] ), .B(n_52688), .Z(n_13442
		));
	notech_ao4 i_618(.A(n_990), .B(n_15156), .C(n_988), .D(n_15177), .Z(n_1089
		));
	notech_reg_set tab24_reg_20(.CP(n_62984), .D(n_13448), .SD(n_62250), .Q(\tab24[20] 
		));
	notech_mux2 i_17886(.S(n_61230), .A(\tab24[20] ), .B(n_52694), .Z(n_13448
		));
	notech_reg_set tab24_reg_21(.CP(n_62985), .D(n_13454), .SD(n_62251), .Q(\tab24[21] 
		));
	notech_mux2 i_17894(.S(n_61230), .A(\tab24[21] ), .B(n_52700), .Z(n_13454
		));
	notech_ao4 i_616(.A(n_998), .B(n_15104), .C(n_996), .D(n_15206), .Z(n_1091
		));
	notech_reg_set tab24_reg_22(.CP(n_62985), .D(n_13460), .SD(n_62251), .Q(\tab24[22] 
		));
	notech_mux2 i_17902(.S(n_61230), .A(\tab24[22] ), .B(n_52706), .Z(n_13460
		));
	notech_reg_set tab24_reg_23(.CP(n_62985), .D(n_13466), .SD(n_62251), .Q(\tab24[23] 
		));
	notech_mux2 i_17910(.S(n_61230), .A(\tab24[23] ), .B(n_52712), .Z(n_13466
		));
	notech_and4 i_620(.A(n_1091), .B(n_1089), .C(n_666), .D(n_669), .Z(n_1093
		));
	notech_reg_set tab24_reg_24(.CP(n_62985), .D(n_13472), .SD(n_62251), .Q(\tab24[24] 
		));
	notech_mux2 i_17918(.S(n_61230), .A(\tab24[24] ), .B(n_52718), .Z(n_13472
		));
	notech_ao4 i_613(.A(n_1003), .B(n_15127), .C(n_1002), .D(n_15082), .Z(n_1094
		));
	notech_reg_set tab24_reg_25(.CP(n_62985), .D(n_13478), .SD(n_62251), .Q(\tab24[25] 
		));
	notech_mux2 i_17926(.S(n_61230), .A(\tab24[25] ), .B(n_52724), .Z(n_13478
		));
	notech_reg_set tab24_reg_26(.CP(n_62985), .D(n_13484), .SD(n_62251), .Q(\tab24[26] 
		));
	notech_mux2 i_17934(.S(n_61230), .A(\tab24[26] ), .B(n_52730), .Z(n_13484
		));
	notech_ao4 i_612(.A(n_62904), .B(n_15305), .C(n_878), .D(n_15249), .Z(n_1096
		));
	notech_reg_set tab24_reg_27(.CP(n_62985), .D(n_13490), .SD(n_62251), .Q(\tab24[27] 
		));
	notech_mux2 i_17942(.S(n_61230), .A(\tab24[27] ), .B(n_52736), .Z(n_13490
		));
	notech_reg_set tab24_reg_28(.CP(n_62985), .D(n_13496), .SD(n_62251), .Q(\tab24[28] 
		));
	notech_mux2 i_17950(.S(n_61230), .A(\tab24[28] ), .B(n_52742), .Z(n_13496
		));
	notech_ao4 i_609(.A(n_990), .B(n_15157), .C(n_988), .D(n_15178), .Z(n_1098
		));
	notech_reg_set tab24_reg_29(.CP(n_62985), .D(n_13502), .SD(n_62251), .Q(\tab24[29] 
		));
	notech_mux2 i_17958(.S(n_61230), .A(\tab24[29] ), .B(n_52748), .Z(n_13502
		));
	notech_reg_set tab24_reg_33(.CP(n_62984), .D(n_13508), .SD(n_62250), .Q(\tab24[33] 
		));
	notech_mux2 i_17966(.S(n_61230), .A(\tab24[33] ), .B(n_52772), .Z(n_13508
		));
	notech_ao4 i_607(.A(n_998), .B(n_15106), .C(n_996), .D(n_15207), .Z(n_1100
		));
	notech_reg_set nnx_tab2_reg_0(.CP(n_62984), .D(n_13514), .SD(n_62250), .Q
		(\nnx_tab2[0] ));
	notech_mux2 i_17974(.S(n_15141), .A(\nnx_tab2[0] ), .B(n_15137), .Z(n_13514
		));
	notech_reg nnx_tab2_reg_1(.CP(n_62984), .D(n_13520), .CD(n_62250), .Q(\nnx_tab2[1] 
		));
	notech_mux2 i_17982(.S(n_15141), .A(\nnx_tab2[1] ), .B(n_15139), .Z(n_13520
		));
	notech_and4 i_611(.A(n_1100), .B(n_1098), .C(n_655), .D(n_658), .Z(n_1102
		));
	notech_reg hit_adr24_reg(.CP(n_62984), .D(n_13526), .CD(n_62250), .Q(hit_adr24
		));
	notech_mux2 i_17990(.S(n_872), .A(hit_add24), .B(hit_adr24), .Z(n_13526)
		);
	notech_ao4 i_604(.A(n_1003), .B(n_15128), .C(n_1002), .D(n_15083), .Z(n_1103
		));
	notech_reg nx_tab2_reg_0(.CP(n_62984), .D(n_13532), .CD(n_62250), .Q(\nx_tab2[0] 
		));
	notech_mux2 i_17998(.S(\nbus_14015[0] ), .A(\nx_tab2[0] ), .B(n_15142), 
		.Z(n_13532));
	notech_reg nx_tab2_reg_1(.CP(n_62984), .D(n_13538), .CD(n_62250), .Q(\nx_tab2[1] 
		));
	notech_mux2 i_18006(.S(\nbus_14015[0] ), .A(\nx_tab2[1] ), .B(n_15144), 
		.Z(n_13538));
	notech_ao4 i_603(.A(n_62908), .B(n_15306), .C(n_62831), .D(n_15250), .Z(n_1105
		));
	notech_reg hit_adr11_reg(.CP(n_62984), .D(n_13544), .CD(n_62250), .Q(hit_adr11
		));
	notech_mux2 i_18014(.S(n_872), .A(hit_add11), .B(hit_adr11), .Z(n_13544)
		);
	notech_reg_set tab12_reg_0(.CP(n_62984), .D(n_13550), .SD(n_62250), .Q(\tab12[0] 
		));
	notech_mux2 i_18022(.S(\nbus_14042[0] ), .A(\tab12[0] ), .B(n_52574), .Z
		(n_13550));
	notech_ao4 i_600(.A(n_990), .B(n_15158), .C(n_988), .D(n_15179), .Z(n_1107
		));
	notech_reg_set tab12_reg_1(.CP(n_62984), .D(n_13556), .SD(n_62250), .Q(\tab12[1] 
		));
	notech_mux2 i_18030(.S(\nbus_14042[0] ), .A(\tab12[1] ), .B(n_52580), .Z
		(n_13556));
	notech_reg_set tab12_reg_2(.CP(n_62984), .D(n_13562), .SD(n_62250), .Q(\tab12[2] 
		));
	notech_mux2 i_18038(.S(\nbus_14042[0] ), .A(\tab12[2] ), .B(n_52586), .Z
		(n_13562));
	notech_ao4 i_598(.A(n_998), .B(n_15107), .C(n_996), .D(n_15208), .Z(n_1109
		));
	notech_reg_set tab12_reg_3(.CP(n_62984), .D(n_13568), .SD(n_62250), .Q(\tab12[3] 
		));
	notech_mux2 i_18046(.S(\nbus_14042[0] ), .A(\tab12[3] ), .B(n_52592), .Z
		(n_13568));
	notech_reg tab12_reg_4(.CP(n_62984), .D(n_13574), .CD(n_62250), .Q(\tab12[4] 
		));
	notech_mux2 i_18054(.S(\nbus_14042[0] ), .A(\tab12[4] ), .B(n_873), .Z(n_13574
		));
	notech_and4 i_602(.A(n_1109), .B(n_1107), .C(n_644), .D(n_647), .Z(n_1111
		));
	notech_reg_set tab12_reg_5(.CP(n_62984), .D(n_13580), .SD(n_62250), .Q(\tab12[5] 
		));
	notech_mux2 i_18062(.S(\nbus_14042[0] ), .A(\tab12[5] ), .B(n_52604), .Z
		(n_13580));
	notech_ao4 i_595(.A(n_1003), .B(n_15129), .C(n_1002), .D(n_15084), .Z(n_1112
		));
	notech_reg_set tab12_reg_6(.CP(n_62984), .D(n_13586), .SD(n_62250), .Q(\tab12[6] 
		));
	notech_mux2 i_18070(.S(\nbus_14042[0] ), .A(\tab12[6] ), .B(n_52610), .Z
		(n_13586));
	notech_reg_set tab12_reg_7(.CP(n_62984), .D(n_13592), .SD(n_62250), .Q(\tab12[7] 
		));
	notech_mux2 i_18078(.S(\nbus_14042[0] ), .A(\tab12[7] ), .B(n_52616), .Z
		(n_13592));
	notech_ao4 i_594(.A(n_62908), .B(n_15307), .C(n_62831), .D(n_15251), .Z(n_1114
		));
	notech_reg_set tab12_reg_8(.CP(n_62956), .D(n_13598), .SD(n_62222), .Q(\tab12[8] 
		));
	notech_mux2 i_18086(.S(\nbus_14042[0] ), .A(\tab12[8] ), .B(n_52622), .Z
		(n_13598));
	notech_reg_set tab12_reg_9(.CP(n_62928), .D(n_13604), .SD(n_62194), .Q(\tab12[9] 
		));
	notech_mux2 i_18094(.S(\nbus_14042[0] ), .A(\tab12[9] ), .B(n_52628), .Z
		(n_13604));
	notech_ao4 i_591(.A(n_990), .B(n_15159), .C(n_988), .D(n_15180), .Z(n_1116
		));
	notech_reg_set tab12_reg_10(.CP(n_62928), .D(n_13610), .SD(n_62194), .Q(\tab12[10] 
		));
	notech_mux2 i_18102(.S(\nbus_14042[0] ), .A(\tab12[10] ), .B(n_52634), .Z
		(n_13610));
	notech_reg_set tab12_reg_11(.CP(n_62929), .D(n_13616), .SD(n_62195), .Q(\tab12[11] 
		));
	notech_mux2 i_18110(.S(\nbus_14042[0] ), .A(\tab12[11] ), .B(n_52640), .Z
		(n_13616));
	notech_ao4 i_589(.A(n_998), .B(n_15109), .C(n_996), .D(n_15209), .Z(n_1118
		));
	notech_reg_set tab12_reg_12(.CP(n_62928), .D(n_13622), .SD(n_62194), .Q(\tab12[12] 
		));
	notech_mux2 i_18118(.S(\nbus_14042[0] ), .A(\tab12[12] ), .B(n_52646), .Z
		(n_13622));
	notech_reg_set tab12_reg_13(.CP(n_62928), .D(n_13628), .SD(n_62194), .Q(\tab12[13] 
		));
	notech_mux2 i_18126(.S(\nbus_14042[0] ), .A(\tab12[13] ), .B(n_52652), .Z
		(n_13628));
	notech_and4 i_593(.A(n_1118), .B(n_1116), .C(n_633), .D(n_636), .Z(n_1120
		));
	notech_reg_set tab12_reg_14(.CP(n_62928), .D(n_13634), .SD(n_62194), .Q(\tab12[14] 
		));
	notech_mux2 i_18134(.S(\nbus_14042[0] ), .A(\tab12[14] ), .B(n_52658), .Z
		(n_13634));
	notech_ao4 i_586(.A(n_1003), .B(n_15130), .C(n_1002), .D(n_15085), .Z(n_1121
		));
	notech_reg_set tab12_reg_15(.CP(n_62928), .D(n_13640), .SD(n_62194), .Q(\tab12[15] 
		));
	notech_mux2 i_18142(.S(\nbus_14042[0] ), .A(\tab12[15] ), .B(n_52664), .Z
		(n_13640));
	notech_reg_set tab12_reg_16(.CP(n_62929), .D(n_13646), .SD(n_62195), .Q(\tab12[16] 
		));
	notech_mux2 i_18150(.S(n_61197), .A(\tab12[16] ), .B(n_52670), .Z(n_13646
		));
	notech_ao4 i_585(.A(n_62908), .B(n_15308), .C(n_62831), .D(n_15252), .Z(n_1123
		));
	notech_reg_set tab12_reg_17(.CP(n_62929), .D(n_13652), .SD(n_62195), .Q(\tab12[17] 
		));
	notech_mux2 i_18158(.S(n_61197), .A(\tab12[17] ), .B(n_52676), .Z(n_13652
		));
	notech_reg_set tab12_reg_18(.CP(n_62929), .D(n_13658), .SD(n_62195), .Q(\tab12[18] 
		));
	notech_mux2 i_18166(.S(n_61197), .A(\tab12[18] ), .B(n_52682), .Z(n_13658
		));
	notech_ao4 i_582(.A(n_990), .B(n_15160), .C(n_988), .D(n_15181), .Z(n_1125
		));
	notech_reg_set tab12_reg_19(.CP(n_62929), .D(n_13664), .SD(n_62195), .Q(\tab12[19] 
		));
	notech_mux2 i_18174(.S(n_61197), .A(\tab12[19] ), .B(n_52688), .Z(n_13664
		));
	notech_reg_set tab12_reg_20(.CP(n_62929), .D(n_13670), .SD(n_62195), .Q(\tab12[20] 
		));
	notech_mux2 i_18182(.S(n_61197), .A(\tab12[20] ), .B(n_52694), .Z(n_13670
		));
	notech_ao4 i_580(.A(n_998), .B(n_15110), .C(n_996), .D(n_15210), .Z(n_1127
		));
	notech_reg_set tab12_reg_21(.CP(n_62929), .D(n_13676), .SD(n_62195), .Q(\tab12[21] 
		));
	notech_mux2 i_18190(.S(n_61197), .A(\tab12[21] ), .B(n_52700), .Z(n_13676
		));
	notech_reg_set tab12_reg_22(.CP(n_62929), .D(n_13682), .SD(n_62195), .Q(\tab12[22] 
		));
	notech_mux2 i_18198(.S(n_61197), .A(\tab12[22] ), .B(n_52706), .Z(n_13682
		));
	notech_and4 i_584(.A(n_1127), .B(n_1125), .C(n_622), .D(n_625), .Z(n_1129
		));
	notech_reg_set tab12_reg_23(.CP(n_62928), .D(n_13688), .SD(n_62194), .Q(\tab12[23] 
		));
	notech_mux2 i_18206(.S(n_61197), .A(\tab12[23] ), .B(n_52712), .Z(n_13688
		));
	notech_ao4 i_577(.A(n_1003), .B(n_15131), .C(n_1002), .D(n_15087), .Z(n_1130
		));
	notech_reg_set tab12_reg_24(.CP(n_62924), .D(n_13694), .SD(n_62190), .Q(\tab12[24] 
		));
	notech_mux2 i_18214(.S(n_61197), .A(\tab12[24] ), .B(n_52718), .Z(n_13694
		));
	notech_reg_set tab12_reg_25(.CP(n_62928), .D(n_13700), .SD(n_62194), .Q(\tab12[25] 
		));
	notech_mux2 i_18222(.S(n_61197), .A(\tab12[25] ), .B(n_52724), .Z(n_13700
		));
	notech_ao4 i_576(.A(n_62908), .B(n_15309), .C(n_62831), .D(n_15253), .Z(n_1132
		));
	notech_reg_set tab12_reg_26(.CP(n_62928), .D(n_13706), .SD(n_62194), .Q(\tab12[26] 
		));
	notech_mux2 i_18230(.S(n_61197), .A(\tab12[26] ), .B(n_52730), .Z(n_13706
		));
	notech_reg_set tab12_reg_27(.CP(n_62924), .D(n_13712), .SD(n_62190), .Q(\tab12[27] 
		));
	notech_mux2 i_18238(.S(n_61197), .A(\tab12[27] ), .B(n_52736), .Z(n_13712
		));
	notech_ao4 i_573(.A(n_990), .B(n_15161), .C(n_988), .D(n_15182), .Z(n_1134
		));
	notech_reg_set tab12_reg_28(.CP(n_62924), .D(n_13718), .SD(n_62190), .Q(\tab12[28] 
		));
	notech_mux2 i_18246(.S(n_61197), .A(\tab12[28] ), .B(n_52742), .Z(n_13718
		));
	notech_reg_set tab12_reg_29(.CP(n_62924), .D(n_13724), .SD(n_62190), .Q(\tab12[29] 
		));
	notech_mux2 i_18254(.S(n_61197), .A(\tab12[29] ), .B(n_52748), .Z(n_13724
		));
	notech_ao4 i_571(.A(n_998), .B(n_15111), .C(n_996), .D(n_15211), .Z(n_1136
		));
	notech_reg_set tab12_reg_33(.CP(n_62924), .D(n_13730), .SD(n_62190), .Q(\tab12[33] 
		));
	notech_mux2 i_18262(.S(n_61197), .A(\tab12[33] ), .B(n_52772), .Z(n_13730
		));
	notech_reg hit_adr12_reg(.CP(n_62928), .D(n_13736), .CD(n_62194), .Q(hit_adr12
		));
	notech_mux2 i_18270(.S(n_872), .A(hit_add12), .B(hit_adr12), .Z(n_13736)
		);
	notech_and4 i_575(.A(n_1136), .B(n_1134), .C(n_611), .D(n_614), .Z(n_1138
		));
	notech_reg_set tab13_reg_0(.CP(n_62928), .D(n_13742), .SD(n_62194), .Q(\tab13[0] 
		));
	notech_mux2 i_18278(.S(\nbus_14026[0] ), .A(\tab13[0] ), .B(n_52574), .Z
		(n_13742));
	notech_ao4 i_568(.A(n_1003), .B(n_15132), .C(n_1002), .D(n_15088), .Z(n_1139
		));
	notech_reg_set tab13_reg_1(.CP(n_62928), .D(n_13748), .SD(n_62194), .Q(\tab13[1] 
		));
	notech_mux2 i_18286(.S(\nbus_14026[0] ), .A(\tab13[1] ), .B(n_52580), .Z
		(n_13748));
	notech_reg_set tab13_reg_2(.CP(n_62928), .D(n_13754), .SD(n_62194), .Q(\tab13[2] 
		));
	notech_mux2 i_18294(.S(\nbus_14026[0] ), .A(\tab13[2] ), .B(n_52586), .Z
		(n_13754));
	notech_ao4 i_567(.A(n_62908), .B(n_15310), .C(n_62831), .D(n_15254), .Z(n_1141
		));
	notech_reg_set tab13_reg_3(.CP(n_62928), .D(n_13760), .SD(n_62194), .Q(\tab13[3] 
		));
	notech_mux2 i_18302(.S(\nbus_14026[0] ), .A(\tab13[3] ), .B(n_52592), .Z
		(n_13760));
	notech_reg tab13_reg_4(.CP(n_62928), .D(n_13766), .CD(n_62194), .Q(\tab13[4] 
		));
	notech_mux2 i_18310(.S(\nbus_14026[0] ), .A(\tab13[4] ), .B(n_873), .Z(n_13766
		));
	notech_ao4 i_564(.A(n_990), .B(n_15162), .C(n_988), .D(n_15183), .Z(n_1143
		));
	notech_reg_set tab13_reg_5(.CP(n_62928), .D(n_13772), .SD(n_62194), .Q(\tab13[5] 
		));
	notech_mux2 i_18318(.S(\nbus_14026[0] ), .A(\tab13[5] ), .B(n_52604), .Z
		(n_13772));
	notech_reg_set tab13_reg_6(.CP(n_62929), .D(n_13778), .SD(n_62195), .Q(\tab13[6] 
		));
	notech_mux2 i_18326(.S(\nbus_14026[0] ), .A(\tab13[6] ), .B(n_52610), .Z
		(n_13778));
	notech_ao4 i_562(.A(n_998), .B(n_15112), .C(n_996), .D(n_15212), .Z(n_1145
		));
	notech_reg_set tab13_reg_7(.CP(n_62933), .D(n_13784), .SD(n_62199), .Q(\tab13[7] 
		));
	notech_mux2 i_18334(.S(\nbus_14026[0] ), .A(\tab13[7] ), .B(n_52616), .Z
		(n_13784));
	notech_reg_set tab13_reg_8(.CP(n_62933), .D(n_13790), .SD(n_62199), .Q(\tab13[8] 
		));
	notech_mux2 i_18342(.S(\nbus_14026[0] ), .A(\tab13[8] ), .B(n_52622), .Z
		(n_13790));
	notech_and4 i_566(.A(n_1145), .B(n_1143), .C(n_600), .D(n_603), .Z(n_1147
		));
	notech_reg_set tab13_reg_9(.CP(n_62933), .D(n_13796), .SD(n_62199), .Q(\tab13[9] 
		));
	notech_mux2 i_18350(.S(\nbus_14026[0] ), .A(\tab13[9] ), .B(n_52628), .Z
		(n_13796));
	notech_ao4 i_559(.A(n_1003), .B(n_15133), .C(n_1002), .D(n_15089), .Z(n_1148
		));
	notech_reg_set tab13_reg_10(.CP(n_62933), .D(n_13802), .SD(n_62199), .Q(\tab13[10] 
		));
	notech_mux2 i_18358(.S(\nbus_14026[0] ), .A(\tab13[10] ), .B(n_52634), .Z
		(n_13802));
	notech_reg_set tab13_reg_11(.CP(n_62933), .D(n_13808), .SD(n_62199), .Q(\tab13[11] 
		));
	notech_mux2 i_18366(.S(\nbus_14026[0] ), .A(\tab13[11] ), .B(n_52640), .Z
		(n_13808));
	notech_ao4 i_558(.A(n_62904), .B(n_15311), .C(n_62831), .D(n_15255), .Z(n_1150
		));
	notech_reg_set tab13_reg_12(.CP(n_62933), .D(n_13814), .SD(n_62199), .Q(\tab13[12] 
		));
	notech_mux2 i_18374(.S(\nbus_14026[0] ), .A(\tab13[12] ), .B(n_52646), .Z
		(n_13814));
	notech_reg_set tab13_reg_13(.CP(n_62933), .D(n_13820), .SD(n_62199), .Q(\tab13[13] 
		));
	notech_mux2 i_18382(.S(\nbus_14026[0] ), .A(\tab13[13] ), .B(n_52652), .Z
		(n_13820));
	notech_ao4 i_555(.A(n_990), .B(n_15163), .C(n_988), .D(n_15184), .Z(n_1152
		));
	notech_reg_set tab13_reg_14(.CP(n_62937), .D(n_13826), .SD(n_62203), .Q(\tab13[14] 
		));
	notech_mux2 i_18390(.S(\nbus_14026[0] ), .A(\tab13[14] ), .B(n_52658), .Z
		(n_13826));
	notech_reg_set tab13_reg_15(.CP(n_62937), .D(n_13832), .SD(n_62203), .Q(\tab13[15] 
		));
	notech_mux2 i_18398(.S(\nbus_14026[0] ), .A(\tab13[15] ), .B(n_52664), .Z
		(n_13832));
	notech_ao4 i_553(.A(n_998), .B(n_15113), .C(n_996), .D(n_15213), .Z(n_1154
		));
	notech_reg_set tab13_reg_16(.CP(n_62937), .D(n_13838), .SD(n_62203), .Q(\tab13[16] 
		));
	notech_mux2 i_18406(.S(n_61175), .A(\tab13[16] ), .B(n_52670), .Z(n_13838
		));
	notech_reg_set tab13_reg_17(.CP(n_62933), .D(n_13844), .SD(n_62199), .Q(\tab13[17] 
		));
	notech_mux2 i_18414(.S(n_61175), .A(\tab13[17] ), .B(n_52676), .Z(n_13844
		));
	notech_and4 i_557(.A(n_1154), .B(n_1152), .C(n_589), .D(n_592), .Z(n_1156
		));
	notech_reg_set tab13_reg_18(.CP(n_62933), .D(n_13850), .SD(n_62199), .Q(\tab13[18] 
		));
	notech_mux2 i_18422(.S(n_61175), .A(\tab13[18] ), .B(n_52682), .Z(n_13850
		));
	notech_ao4 i_550(.A(n_1003), .B(n_15134), .C(n_1002), .D(n_15090), .Z(n_1157
		));
	notech_reg_set tab13_reg_19(.CP(n_62933), .D(n_13856), .SD(n_62199), .Q(\tab13[19] 
		));
	notech_mux2 i_18430(.S(n_61175), .A(\tab13[19] ), .B(n_52688), .Z(n_13856
		));
	notech_reg_set tab13_reg_20(.CP(n_62933), .D(n_13862), .SD(n_62199), .Q(\tab13[20] 
		));
	notech_mux2 i_18438(.S(n_61175), .A(\tab13[20] ), .B(n_52694), .Z(n_13862
		));
	notech_ao4 i_549(.A(n_62904), .B(n_15312), .C(n_62831), .D(n_15256), .Z(n_1159
		));
	notech_reg_set tab13_reg_21(.CP(n_62933), .D(n_13868), .SD(n_62199), .Q(\tab13[21] 
		));
	notech_mux2 i_18446(.S(n_61175), .A(\tab13[21] ), .B(n_52700), .Z(n_13868
		));
	notech_reg_set tab13_reg_22(.CP(n_62929), .D(n_13874), .SD(n_62195), .Q(\tab13[22] 
		));
	notech_mux2 i_18454(.S(n_61175), .A(\tab13[22] ), .B(n_52706), .Z(n_13874
		));
	notech_ao4 i_546(.A(n_990), .B(n_15164), .C(n_988), .D(n_15185), .Z(n_1161
		));
	notech_reg_set tab13_reg_23(.CP(n_62929), .D(n_13880), .SD(n_62195), .Q(\tab13[23] 
		));
	notech_mux2 i_18462(.S(n_61175), .A(\tab13[23] ), .B(n_52712), .Z(n_13880
		));
	notech_reg_set tab13_reg_24(.CP(n_62929), .D(n_13886), .SD(n_62195), .Q(\tab13[24] 
		));
	notech_mux2 i_18470(.S(n_61175), .A(\tab13[24] ), .B(n_52718), .Z(n_13886
		));
	notech_ao4 i_544(.A(n_998), .B(n_15114), .C(n_996), .D(n_15214), .Z(n_1163
		));
	notech_reg_set tab13_reg_25(.CP(n_62929), .D(n_13892), .SD(n_62195), .Q(\tab13[25] 
		));
	notech_mux2 i_18478(.S(n_61175), .A(\tab13[25] ), .B(n_52724), .Z(n_13892
		));
	notech_reg_set tab13_reg_26(.CP(n_62929), .D(n_13898), .SD(n_62195), .Q(\tab13[26] 
		));
	notech_mux2 i_18486(.S(n_61175), .A(\tab13[26] ), .B(n_52730), .Z(n_13898
		));
	notech_and4 i_548(.A(n_1163), .B(n_1161), .C(n_578), .D(n_581), .Z(n_1165
		));
	notech_reg_set tab13_reg_27(.CP(n_62929), .D(n_13904), .SD(n_62195), .Q(\tab13[27] 
		));
	notech_mux2 i_18494(.S(n_61175), .A(\tab13[27] ), .B(n_52736), .Z(n_13904
		));
	notech_ao4 i_541(.A(n_1003), .B(n_15135), .C(n_1002), .D(n_15091), .Z(n_1166
		));
	notech_reg_set tab13_reg_28(.CP(n_62929), .D(n_13910), .SD(n_62195), .Q(\tab13[28] 
		));
	notech_mux2 i_18502(.S(n_61175), .A(\tab13[28] ), .B(n_52742), .Z(n_13910
		));
	notech_reg_set tab13_reg_29(.CP(n_62933), .D(n_13916), .SD(n_62199), .Q(\tab13[29] 
		));
	notech_mux2 i_18510(.S(n_61175), .A(\tab13[29] ), .B(n_52748), .Z(n_13916
		));
	notech_ao4 i_540(.A(n_62904), .B(n_15313), .C(n_878), .D(n_15257), .Z(n_1168
		));
	notech_reg_set tab13_reg_33(.CP(n_62933), .D(n_13922), .SD(n_62199), .Q(\tab13[33] 
		));
	notech_mux2 i_18518(.S(n_61175), .A(\tab13[33] ), .B(n_52772), .Z(n_13922
		));
	notech_reg hit_adr13_reg(.CP(n_62933), .D(n_13928), .CD(n_62199), .Q(hit_adr13
		));
	notech_mux2 i_18526(.S(n_872), .A(hit_add13), .B(hit_adr13), .Z(n_13928)
		);
	notech_ao4 i_537(.A(n_990), .B(n_15165), .C(n_988), .D(n_15186), .Z(n_1170
		));
	notech_reg_set tab14_reg_0(.CP(n_62933), .D(n_13934), .SD(n_62199), .Q(\tab14[0] 
		));
	notech_mux2 i_18534(.S(\nbus_14040[0] ), .A(\tab14[0] ), .B(n_52574), .Z
		(n_13934));
	notech_reg_set tab14_reg_1(.CP(n_62929), .D(n_13940), .SD(n_62195), .Q(\tab14[1] 
		));
	notech_mux2 i_18542(.S(\nbus_14040[0] ), .A(\tab14[1] ), .B(n_52580), .Z
		(n_13940));
	notech_ao4 i_535(.A(n_998), .B(n_15115), .C(n_996), .D(n_15215), .Z(n_1172
		));
	notech_reg_set tab14_reg_2(.CP(n_62933), .D(n_13946), .SD(n_62199), .Q(\tab14[2] 
		));
	notech_mux2 i_18550(.S(\nbus_14040[0] ), .A(\tab14[2] ), .B(n_52586), .Z
		(n_13946));
	notech_reg_set tab14_reg_3(.CP(n_62933), .D(n_13952), .SD(n_62199), .Q(\tab14[3] 
		));
	notech_mux2 i_18558(.S(\nbus_14040[0] ), .A(\tab14[3] ), .B(n_52592), .Z
		(n_13952));
	notech_and4 i_539(.A(n_1172), .B(n_1170), .C(n_567), .D(n_570), .Z(n_1174
		));
	notech_reg tab14_reg_4(.CP(n_62919), .D(n_13958), .CD(n_62185), .Q(\tab14[4] 
		));
	notech_mux2 i_18566(.S(\nbus_14040[0] ), .A(\tab14[4] ), .B(n_873), .Z(n_13958
		));
	notech_ao4 i_532(.A(n_1003), .B(n_15136), .C(n_1002), .D(n_15092), .Z(n_1175
		));
	notech_reg_set tab14_reg_5(.CP(n_62919), .D(n_13964), .SD(n_62185), .Q(\tab14[5] 
		));
	notech_mux2 i_18574(.S(\nbus_14040[0] ), .A(\tab14[5] ), .B(n_52604), .Z
		(n_13964));
	notech_reg_set tab14_reg_6(.CP(n_62919), .D(n_13970), .SD(n_62185), .Q(\tab14[6] 
		));
	notech_mux2 i_18582(.S(\nbus_14040[0] ), .A(\tab14[6] ), .B(n_52610), .Z
		(n_13970));
	notech_ao4 i_531(.A(n_62908), .B(n_15314), .C(n_62831), .D(n_15258), .Z(n_1177
		));
	notech_reg_set tab14_reg_7(.CP(n_62919), .D(n_13976), .SD(n_62185), .Q(\tab14[7] 
		));
	notech_mux2 i_18590(.S(\nbus_14040[0] ), .A(\tab14[7] ), .B(n_52616), .Z
		(n_13976));
	notech_reg_set tab14_reg_8(.CP(n_62915), .D(n_13982), .SD(n_62181), .Q(\tab14[8] 
		));
	notech_mux2 i_18598(.S(\nbus_14040[0] ), .A(\tab14[8] ), .B(n_52622), .Z
		(n_13982));
	notech_ao4 i_75720(.A(n_15262), .B(n_15341), .C(n_15100), .D(n_15342), .Z
		(oread_req101009));
	notech_reg_set tab14_reg_9(.CP(n_62919), .D(n_13988), .SD(n_62185), .Q(\tab14[9] 
		));
	notech_mux2 i_18606(.S(\nbus_14040[0] ), .A(\tab14[9] ), .B(n_52628), .Z
		(n_13988));
	notech_nand3 i_77553(.A(n_532), .B(n_388), .C(n_531), .Z(\nbus_14024[0] 
		));
	notech_reg_set tab14_reg_10(.CP(n_62919), .D(n_13994), .SD(n_62185), .Q(\tab14[10] 
		));
	notech_mux2 i_18614(.S(\nbus_14040[0] ), .A(\tab14[10] ), .B(n_52634), .Z
		(n_13994));
	notech_nand3 i_77031(.A(n_532), .B(n_388), .C(n_528), .Z(\nbus_14016[0] 
		));
	notech_reg_set tab14_reg_11(.CP(n_62919), .D(n_14000), .SD(n_62185), .Q(\tab14[11] 
		));
	notech_mux2 i_18622(.S(\nbus_14040[0] ), .A(\tab14[11] ), .B(n_52640), .Z
		(n_14000));
	notech_nand3 i_77181(.A(n_509), .B(n_388), .C(n_508), .Z(\nbus_14019[0] 
		));
	notech_reg_set tab14_reg_12(.CP(n_62919), .D(n_14006), .SD(n_62185), .Q(\tab14[12] 
		));
	notech_mux2 i_18630(.S(\nbus_14040[0] ), .A(\tab14[12] ), .B(n_52646), .Z
		(n_14006));
	notech_nand3 i_77444(.A(n_509), .B(n_388), .C(n_505), .Z(\nbus_14023[0] 
		));
	notech_reg_set tab14_reg_13(.CP(n_62919), .D(n_14012), .SD(n_62185), .Q(\tab14[13] 
		));
	notech_mux2 i_18638(.S(\nbus_14040[0] ), .A(\tab14[13] ), .B(n_52652), .Z
		(n_14012));
	notech_nand3 i_77672(.A(n_509), .B(n_388), .C(n_504), .Z(\nbus_14025[0] 
		));
	notech_reg_set tab14_reg_14(.CP(n_62919), .D(n_14018), .SD(n_62185), .Q(\tab14[14] 
		));
	notech_mux2 i_18646(.S(\nbus_14040[0] ), .A(\tab14[14] ), .B(n_52658), .Z
		(n_14018));
	notech_nand3 i_78139(.A(n_509), .B(n_388), .C(n_503), .Z(\nbus_14039[0] 
		));
	notech_reg_set tab14_reg_15(.CP(n_62919), .D(n_14024), .SD(n_62185), .Q(\tab14[15] 
		));
	notech_mux2 i_18654(.S(\nbus_14040[0] ), .A(\tab14[15] ), .B(n_52664), .Z
		(n_14024));
	notech_ao4 i_78400(.A(n_899), .B(n_900), .C(n_913), .D(n_15086), .Z(\nbus_14041[0] 
		));
	notech_reg_set tab14_reg_16(.CP(n_62919), .D(n_14030), .SD(n_62185), .Q(\tab14[16] 
		));
	notech_mux2 i_18662(.S(n_61164), .A(\tab14[16] ), .B(n_52670), .Z(n_14030
		));
	notech_nand2 i_77001(.A(n_913), .B(n_901), .Z(\nbus_14015[0] ));
	notech_reg_set tab14_reg_17(.CP(n_62919), .D(n_14036), .SD(n_62185), .Q(\tab14[17] 
		));
	notech_mux2 i_18670(.S(n_61164), .A(\tab14[17] ), .B(n_52676), .Z(n_14036
		));
	notech_nand3 i_78419(.A(n_485), .B(n_388), .C(n_484), .Z(\nbus_14042[0] 
		));
	notech_reg_set tab14_reg_18(.CP(n_62915), .D(n_14042), .SD(n_62181), .Q(\tab14[18] 
		));
	notech_mux2 i_18678(.S(n_61164), .A(\tab14[18] ), .B(n_52682), .Z(n_14042
		));
	notech_nand3 i_77784(.A(n_485), .B(n_388), .C(n_483), .Z(\nbus_14026[0] 
		));
	notech_reg_set tab14_reg_19(.CP(n_62915), .D(n_14048), .SD(n_62181), .Q(\tab14[19] 
		));
	notech_mux2 i_18686(.S(n_61164), .A(\tab14[19] ), .B(n_52688), .Z(n_14048
		));
	notech_nand3 i_78251(.A(n_485), .B(n_388), .C(n_482), .Z(\nbus_14040[0] 
		));
	notech_reg_set tab14_reg_20(.CP(n_62915), .D(n_14054), .SD(n_62181), .Q(\tab14[20] 
		));
	notech_mux2 i_18694(.S(n_61164), .A(\tab14[20] ), .B(n_52694), .Z(n_14054
		));
	notech_ao4 i_76878(.A(n_899), .B(n_919), .C(n_913), .D(n_15071), .Z(\nbus_14014[0] 
		));
	notech_reg_set tab14_reg_21(.CP(n_62915), .D(n_14060), .SD(n_62181), .Q(\tab14[21] 
		));
	notech_mux2 i_18702(.S(n_61164), .A(\tab14[21] ), .B(n_52700), .Z(n_14060
		));
	notech_nand2 i_77291(.A(n_913), .B(n_920), .Z(\nbus_14020[0] ));
	notech_reg_set tab14_reg_22(.CP(n_62915), .D(n_14066), .SD(n_62181), .Q(\tab14[22] 
		));
	notech_mux2 i_18710(.S(n_61164), .A(\tab14[22] ), .B(n_52706), .Z(n_14066
		));
	notech_nand3 i_78017(.A(n_485), .B(n_388), .C(n_464), .Z(\nbus_14038[0] 
		));
	notech_reg_set tab14_reg_23(.CP(n_62915), .D(n_14072), .SD(n_62181), .Q(\tab14[23] 
		));
	notech_mux2 i_18718(.S(n_61164), .A(\tab14[23] ), .B(n_52712), .Z(n_14072
		));
	notech_nand2 i_77303(.A(n_893), .B(n_462), .Z(\nbus_14021[0] ));
	notech_reg_set tab14_reg_24(.CP(n_62915), .D(n_14078), .SD(n_62181), .Q(\tab14[24] 
		));
	notech_mux2 i_18726(.S(n_61164), .A(\tab14[24] ), .B(n_52718), .Z(n_14078
		));
	notech_ao4 i_76990(.A(n_461), .B(n_932), .C(n_887), .D(n_15259), .Z(n_52233
		));
	notech_reg_set tab14_reg_25(.CP(n_62915), .D(n_14084), .SD(n_62181), .Q(\tab14[25] 
		));
	notech_mux2 i_18734(.S(n_61164), .A(\tab14[25] ), .B(n_52724), .Z(n_14084
		));
	notech_nand3 i_77159(.A(n_62831), .B(n_52233), .C(n_945), .Z(\nbus_14018[0] 
		));
	notech_reg_set tab14_reg_26(.CP(n_62915), .D(n_14090), .SD(n_62181), .Q(\tab14[26] 
		));
	notech_mux2 i_18742(.S(n_61164), .A(\tab14[26] ), .B(n_52730), .Z(n_14090
		));
	notech_nand2 i_76210(.A(n_938), .B(n_912), .Z(n_52519));
	notech_reg_set tab14_reg_27(.CP(n_62915), .D(n_14096), .SD(n_62181), .Q(\tab14[27] 
		));
	notech_mux2 i_18750(.S(n_61164), .A(\tab14[27] ), .B(n_52736), .Z(n_14096
		));
	notech_ao4 i_77338(.A(n_876), .B(data_miss[5]), .C(n_899), .D(n_934), .Z
		(\nbus_14022[0] ));
	notech_reg_set tab14_reg_28(.CP(n_62915), .D(n_14102), .SD(n_62181), .Q(\tab14[28] 
		));
	notech_mux2 i_18758(.S(n_61164), .A(\tab14[28] ), .B(n_52742), .Z(n_14102
		));
	notech_ao4 i_77139(.A(n_15341), .B(n_15261), .C(n_887), .D(n_15259), .Z(n_52516
		));
	notech_reg_set tab14_reg_29(.CP(n_62915), .D(n_14108), .SD(n_62181), .Q(\tab14[29] 
		));
	notech_mux2 i_18766(.S(n_61164), .A(\tab14[29] ), .B(n_52748), .Z(n_14108
		));
	notech_nand2 i_322205(.A(n_975), .B(n_400), .Z(addr_phys[2]));
	notech_reg_set tab14_reg_33(.CP(n_62915), .D(n_14114), .SD(n_62181), .Q(\tab14[33] 
		));
	notech_mux2 i_18774(.S(n_61164), .A(\tab14[33] ), .B(n_52772), .Z(n_14114
		));
	notech_nand2 i_422206(.A(n_976), .B(n_398), .Z(addr_phys[3]));
	notech_reg hit_adr14_reg(.CP(n_62915), .D(n_14120), .CD(n_62181), .Q(hit_adr14
		));
	notech_mux2 i_18782(.S(n_872), .A(hit_add14), .B(hit_adr14), .Z(n_14120)
		);
	notech_nand2 i_522207(.A(n_977), .B(n_397), .Z(addr_phys[4]));
	notech_reg_set nnx_tab1_reg_0(.CP(n_62915), .D(n_14126), .SD(n_62181), .Q
		(\nnx_tab1[0] ));
	notech_mux2 i_18790(.S(n_15191), .A(\nnx_tab1[0] ), .B(n_15187), .Z(n_14126
		));
	notech_nand2 i_622208(.A(n_978), .B(n_396), .Z(addr_phys[5]));
	notech_reg nnx_tab1_reg_1(.CP(n_62919), .D(n_14132), .CD(n_62185), .Q(\nnx_tab1[1] 
		));
	notech_mux2 i_18798(.S(n_15191), .A(\nnx_tab1[1] ), .B(n_15189), .Z(n_14132
		));
	notech_nand2 i_722209(.A(n_979), .B(n_395), .Z(addr_phys[6]));
	notech_reg nx_tab1_reg_0(.CP(n_62924), .D(n_14138), .CD(n_62190), .Q(\nx_tab1[0] 
		));
	notech_mux2 i_18806(.S(\nbus_14020[0] ), .A(\nx_tab1[0] ), .B(n_15192), 
		.Z(n_14138));
	notech_nand2 i_822210(.A(n_980), .B(n_394), .Z(addr_phys[7]));
	notech_reg nx_tab1_reg_1(.CP(n_62924), .D(n_14144), .CD(n_62190), .Q(\nx_tab1[1] 
		));
	notech_mux2 i_18814(.S(\nbus_14020[0] ), .A(\nx_tab1[1] ), .B(n_15194), 
		.Z(n_14144));
	notech_nand2 i_922211(.A(n_981), .B(n_393), .Z(addr_phys[8]));
	notech_reg_set tab11_reg_0(.CP(n_62924), .D(n_14150), .SD(n_62190), .Q(\tab11[0] 
		));
	notech_mux2 i_18822(.S(\nbus_14038[0] ), .A(\tab11[0] ), .B(n_52574), .Z
		(n_14150));
	notech_nand2 i_1022212(.A(n_982), .B(n_392), .Z(addr_phys[9]));
	notech_reg_set tab11_reg_1(.CP(n_62924), .D(n_14156), .SD(n_62190), .Q(\tab11[1] 
		));
	notech_mux2 i_18830(.S(\nbus_14038[0] ), .A(\tab11[1] ), .B(n_52580), .Z
		(n_14156));
	notech_nand2 i_1122213(.A(n_983), .B(n_391), .Z(addr_phys[10]));
	notech_reg_set tab11_reg_2(.CP(n_62920), .D(n_14162), .SD(n_62186), .Q(\tab11[2] 
		));
	notech_mux2 i_18838(.S(\nbus_14038[0] ), .A(\tab11[2] ), .B(n_52586), .Z
		(n_14162));
	notech_nand2 i_1222214(.A(n_984), .B(n_390), .Z(addr_phys[11]));
	notech_reg_set tab11_reg_3(.CP(n_62920), .D(n_14168), .SD(n_62186), .Q(\tab11[3] 
		));
	notech_mux2 i_18846(.S(\nbus_14038[0] ), .A(\tab11[3] ), .B(n_52592), .Z
		(n_14168));
	notech_and4 i_1322215(.A(n_1004), .B(n_1006), .C(n_1001), .D(n_773), .Z(addr_phys_12101010
		));
	notech_reg tab11_reg_4(.CP(n_62920), .D(n_14174), .CD(n_62186), .Q(\tab11[4] 
		));
	notech_mux2 i_18854(.S(\nbus_14038[0] ), .A(\tab11[4] ), .B(n_873), .Z(n_14174
		));
	notech_and4 i_1422216(.A(n_1013), .B(n_1015), .C(n_1012), .D(n_762), .Z(addr_phys_13101011
		));
	notech_reg_set tab11_reg_5(.CP(n_62924), .D(n_14180), .SD(n_62190), .Q(\tab11[5] 
		));
	notech_mux2 i_18862(.S(\nbus_14038[0] ), .A(\tab11[5] ), .B(n_52604), .Z
		(n_14180));
	notech_and4 i_1522217(.A(n_1022), .B(n_1024), .C(n_1021), .D(n_751), .Z(addr_phys_14101012
		));
	notech_reg_set tab11_reg_6(.CP(n_62924), .D(n_14186), .SD(n_62190), .Q(\tab11[6] 
		));
	notech_mux2 i_18870(.S(\nbus_14038[0] ), .A(\tab11[6] ), .B(n_52610), .Z
		(n_14186));
	notech_and4 i_1622218(.A(n_1031), .B(n_1033), .C(n_1030), .D(n_740), .Z(addr_phys_15101013
		));
	notech_reg_set tab11_reg_7(.CP(n_62924), .D(n_14192), .SD(n_62190), .Q(\tab11[7] 
		));
	notech_mux2 i_18878(.S(\nbus_14038[0] ), .A(\tab11[7] ), .B(n_52616), .Z
		(n_14192));
	notech_and4 i_1722219(.A(n_1040), .B(n_1042), .C(n_1039), .D(n_729), .Z(addr_phys_16101014
		));
	notech_reg_set tab11_reg_8(.CP(n_62924), .D(n_14198), .SD(n_62190), .Q(\tab11[8] 
		));
	notech_mux2 i_18886(.S(\nbus_14038[0] ), .A(\tab11[8] ), .B(n_52622), .Z
		(n_14198));
	notech_and4 i_1822220(.A(n_1049), .B(n_1051), .C(n_1048), .D(n_718), .Z(addr_phys_17101015
		));
	notech_reg_set tab11_reg_9(.CP(n_62924), .D(n_14204), .SD(n_62190), .Q(\tab11[9] 
		));
	notech_mux2 i_18894(.S(\nbus_14038[0] ), .A(\tab11[9] ), .B(n_52628), .Z
		(n_14204));
	notech_and4 i_1922221(.A(n_1058), .B(n_1060), .C(n_1057), .D(n_707), .Z(addr_phys_18101016
		));
	notech_reg_set tab11_reg_10(.CP(n_62924), .D(n_14210), .SD(n_62190), .Q(\tab11[10] 
		));
	notech_mux2 i_18902(.S(\nbus_14038[0] ), .A(\tab11[10] ), .B(n_52634), .Z
		(n_14210));
	notech_and4 i_2022222(.A(n_1067), .B(n_1069), .C(n_1066), .D(n_696), .Z(addr_phys_19101017
		));
	notech_reg_set tab11_reg_11(.CP(n_62924), .D(n_14216), .SD(n_62190), .Q(\tab11[11] 
		));
	notech_mux2 i_18910(.S(\nbus_14038[0] ), .A(\tab11[11] ), .B(n_52640), .Z
		(n_14216));
	notech_and4 i_2122223(.A(n_1076), .B(n_1078), .C(n_1075), .D(n_685), .Z(addr_phys_20101018
		));
	notech_reg_set tab11_reg_12(.CP(n_62920), .D(n_14222), .SD(n_62186), .Q(\tab11[12] 
		));
	notech_mux2 i_18918(.S(\nbus_14038[0] ), .A(\tab11[12] ), .B(n_52646), .Z
		(n_14222));
	notech_and4 i_2222224(.A(n_1085), .B(n_1087), .C(n_1084), .D(n_674), .Z(addr_phys_21101019
		));
	notech_reg_set tab11_reg_13(.CP(n_62920), .D(n_14228), .SD(n_62186), .Q(\tab11[13] 
		));
	notech_mux2 i_18926(.S(\nbus_14038[0] ), .A(\tab11[13] ), .B(n_52652), .Z
		(n_14228));
	notech_and4 i_2322225(.A(n_1094), .B(n_1096), .C(n_1093), .D(n_663), .Z(addr_phys_22101020
		));
	notech_reg_set tab11_reg_14(.CP(n_62920), .D(n_14234), .SD(n_62186), .Q(\tab11[14] 
		));
	notech_mux2 i_18934(.S(\nbus_14038[0] ), .A(\tab11[14] ), .B(n_52658), .Z
		(n_14234));
	notech_and4 i_2422226(.A(n_1103), .B(n_1105), .C(n_1102), .D(n_652), .Z(addr_phys_23101021
		));
	notech_reg_set tab11_reg_15(.CP(n_62920), .D(n_14240), .SD(n_62186), .Q(\tab11[15] 
		));
	notech_mux2 i_18942(.S(\nbus_14038[0] ), .A(\tab11[15] ), .B(n_52664), .Z
		(n_14240));
	notech_and4 i_2522227(.A(n_1112), .B(n_1114), .C(n_1111), .D(n_641), .Z(addr_phys_24101022
		));
	notech_reg_set tab11_reg_16(.CP(n_62920), .D(n_14246), .SD(n_62186), .Q(\tab11[16] 
		));
	notech_mux2 i_18950(.S(n_61186), .A(\tab11[16] ), .B(n_52670), .Z(n_14246
		));
	notech_and4 i_2622228(.A(n_1121), .B(n_1123), .C(n_1120), .D(n_630), .Z(addr_phys_25101023
		));
	notech_reg_set tab11_reg_17(.CP(n_62919), .D(n_14252), .SD(n_62185), .Q(\tab11[17] 
		));
	notech_mux2 i_18958(.S(n_61186), .A(\tab11[17] ), .B(n_52676), .Z(n_14252
		));
	notech_and4 i_2722229(.A(n_1130), .B(n_1132), .C(n_1129), .D(n_619), .Z(addr_phys_26101024
		));
	notech_reg_set tab11_reg_18(.CP(n_62919), .D(n_14258), .SD(n_62185), .Q(\tab11[18] 
		));
	notech_mux2 i_18966(.S(n_61186), .A(\tab11[18] ), .B(n_52682), .Z(n_14258
		));
	notech_and4 i_2822230(.A(n_1139), .B(n_1141), .C(n_1138), .D(n_608), .Z(addr_phys_27101025
		));
	notech_reg_set tab11_reg_19(.CP(n_62920), .D(n_14264), .SD(n_62186), .Q(\tab11[19] 
		));
	notech_mux2 i_18974(.S(n_61186), .A(\tab11[19] ), .B(n_52688), .Z(n_14264
		));
	notech_and4 i_2922231(.A(n_1148), .B(n_1150), .C(n_1147), .D(n_597), .Z(addr_phys_28101026
		));
	notech_reg_set tab11_reg_20(.CP(n_62920), .D(n_14270), .SD(n_62186), .Q(\tab11[20] 
		));
	notech_mux2 i_18982(.S(n_61186), .A(\tab11[20] ), .B(n_52694), .Z(n_14270
		));
	notech_and4 i_3022232(.A(n_1157), .B(n_1159), .C(n_1156), .D(n_586), .Z(addr_phys_29101027
		));
	notech_reg_set tab11_reg_21(.CP(n_62920), .D(n_14276), .SD(n_62186), .Q(\tab11[21] 
		));
	notech_mux2 i_18990(.S(n_61186), .A(\tab11[21] ), .B(n_52700), .Z(n_14276
		));
	notech_and4 i_3122233(.A(n_1166), .B(n_1168), .C(n_1165), .D(n_575), .Z(addr_phys_30101028
		));
	notech_reg_set tab11_reg_22(.CP(n_62920), .D(n_14282), .SD(n_62186), .Q(\tab11[22] 
		));
	notech_mux2 i_18998(.S(n_61186), .A(\tab11[22] ), .B(n_52706), .Z(n_14282
		));
	notech_and4 i_3222234(.A(n_1175), .B(n_1177), .C(n_1174), .D(n_564), .Z(addr_phys_31101029
		));
	notech_reg_set tab11_reg_23(.CP(n_62920), .D(n_14288), .SD(n_62186), .Q(\tab11[23] 
		));
	notech_mux2 i_19006(.S(n_61186), .A(\tab11[23] ), .B(n_52712), .Z(n_14288
		));
	notech_mux2 i_122728(.S(n_62873), .A(iDaddr[12]), .B(iDaddr_f[12]), .Z(\tab11_0[0] 
		));
	notech_reg_set tab11_reg_24(.CP(n_62920), .D(n_14294), .SD(n_62186), .Q(\tab11[24] 
		));
	notech_mux2 i_19014(.S(n_61186), .A(\tab11[24] ), .B(n_52718), .Z(n_14294
		));
	notech_mux2 i_222729(.S(n_62873), .A(iDaddr[13]), .B(iDaddr_f[13]), .Z(\tab11_0[1] 
		));
	notech_reg_set tab11_reg_25(.CP(n_62920), .D(n_14300), .SD(n_62186), .Q(\tab11[25] 
		));
	notech_mux2 i_19022(.S(n_61186), .A(\tab11[25] ), .B(n_52724), .Z(n_14300
		));
	notech_mux2 i_322730(.S(n_62873), .A(iDaddr[14]), .B(iDaddr_f[14]), .Z(\tab11_0[2] 
		));
	notech_reg_set tab11_reg_26(.CP(n_62920), .D(n_14306), .SD(n_62186), .Q(\tab11[26] 
		));
	notech_mux2 i_19030(.S(n_61186), .A(\tab11[26] ), .B(n_52730), .Z(n_14306
		));
	notech_mux2 i_422731(.S(n_62873), .A(iDaddr[15]), .B(iDaddr_f[15]), .Z(\tab11_0[3] 
		));
	notech_reg_set tab11_reg_27(.CP(n_62937), .D(n_14312), .SD(n_62203), .Q(\tab11[27] 
		));
	notech_mux2 i_19038(.S(n_61186), .A(\tab11[27] ), .B(n_52736), .Z(n_14312
		));
	notech_mux2 i_522732(.S(n_62873), .A(iDaddr[16]), .B(iDaddr_f[16]), .Z(\tab11_0[4] 
		));
	notech_reg_set tab11_reg_28(.CP(n_62948), .D(n_14318), .SD(n_62214), .Q(\tab11[28] 
		));
	notech_mux2 i_19046(.S(n_61186), .A(\tab11[28] ), .B(n_52742), .Z(n_14318
		));
	notech_mux2 i_622733(.S(n_62873), .A(iDaddr[17]), .B(iDaddr_f[17]), .Z(\tab11_0[5] 
		));
	notech_reg_set tab11_reg_29(.CP(n_62948), .D(n_14324), .SD(n_62214), .Q(\tab11[29] 
		));
	notech_mux2 i_19054(.S(n_61186), .A(\tab11[29] ), .B(n_52748), .Z(n_14324
		));
	notech_mux2 i_722734(.S(n_62873), .A(iDaddr[18]), .B(iDaddr_f[18]), .Z(\tab11_0[6] 
		));
	notech_reg_set tab11_reg_33(.CP(n_62948), .D(n_14330), .SD(n_62214), .Q(\tab11[33] 
		));
	notech_mux2 i_19062(.S(n_61186), .A(\tab11[33] ), .B(n_52772), .Z(n_14330
		));
	notech_mux2 i_822735(.S(n_62873), .A(iDaddr[19]), .B(iDaddr_f[19]), .Z(\tab11_0[7] 
		));
	notech_reg fsm5_cnt_reg_0(.CP(n_62948), .D(n_14336), .CD(n_62214), .Q(fsm5_cnt
		[0]));
	notech_mux2 i_19070(.S(\nbus_14021[0] ), .A(fsm5_cnt[0]), .B(n_863), .Z(n_14336
		));
	notech_mux2 i_922736(.S(n_62873), .A(iDaddr[20]), .B(iDaddr_f[20]), .Z(\tab11_0[8] 
		));
	notech_reg fsm5_cnt_reg_1(.CP(n_62948), .D(n_14342), .CD(n_62214), .Q(fsm5_cnt
		[1]));
	notech_mux2 i_19078(.S(\nbus_14021[0] ), .A(fsm5_cnt[1]), .B(n_864), .Z(n_14342
		));
	notech_mux2 i_1022737(.S(n_62873), .A(iDaddr[21]), .B(iDaddr_f[21]), .Z(\tab11_0[9] 
		));
	notech_reg fsm5_cnt_reg_2(.CP(n_62948), .D(n_14348), .CD(n_62214), .Q(fsm5_cnt
		[2]));
	notech_mux2 i_19086(.S(\nbus_14021[0] ), .A(fsm5_cnt[2]), .B(n_865), .Z(n_14348
		));
	notech_mux2 i_1122738(.S(n_62878), .A(iDaddr[22]), .B(iDaddr_f[22]), .Z(\dir1_0[0] 
		));
	notech_reg fsm5_cnt_reg_3(.CP(n_62948), .D(n_14354), .CD(n_62214), .Q(fsm5_cnt
		[3]));
	notech_mux2 i_19094(.S(\nbus_14021[0] ), .A(fsm5_cnt[3]), .B(n_866), .Z(n_14354
		));
	notech_mux2 i_1222739(.S(n_62878), .A(iDaddr[23]), .B(iDaddr_f[23]), .Z(\dir1_0[1] 
		));
	notech_reg fsm5_cnt_reg_4(.CP(n_62948), .D(n_14360), .CD(n_62214), .Q(fsm5_cnt
		[4]));
	notech_mux2 i_19102(.S(\nbus_14021[0] ), .A(fsm5_cnt[4]), .B(n_867), .Z(n_14360
		));
	notech_mux2 i_1322740(.S(n_62878), .A(iDaddr[24]), .B(iDaddr_f[24]), .Z(\dir1_0[2] 
		));
	notech_reg fsm5_cnt_reg_5(.CP(n_62952), .D(n_14366), .CD(n_62218), .Q(fsm5_cnt
		[5]));
	notech_mux2 i_19110(.S(\nbus_14021[0] ), .A(fsm5_cnt[5]), .B(n_868), .Z(n_14366
		));
	notech_mux2 i_1422741(.S(n_62878), .A(iDaddr[25]), .B(iDaddr_f[25]), .Z(\dir1_0[3] 
		));
	notech_reg fsm5_cnt_reg_6(.CP(n_62952), .D(n_14372), .CD(n_62218), .Q(fsm5_cnt
		[6]));
	notech_mux2 i_19118(.S(\nbus_14021[0] ), .A(fsm5_cnt[6]), .B(n_869), .Z(n_14372
		));
	notech_mux2 i_1522742(.S(n_62878), .A(iDaddr[26]), .B(iDaddr_f[26]), .Z(\dir1_0[4] 
		));
	notech_reg fsm5_cnt_reg_7(.CP(n_62948), .D(n_14378), .CD(n_62214), .Q(fsm5_cnt
		[7]));
	notech_mux2 i_19126(.S(\nbus_14021[0] ), .A(fsm5_cnt[7]), .B(n_870), .Z(n_14378
		));
	notech_mux2 i_1622743(.S(n_62878), .A(iDaddr[27]), .B(iDaddr_f[27]), .Z(\dir1_0[5] 
		));
	notech_reg fsm5_cnt_reg_8(.CP(n_62948), .D(n_14384), .CD(n_62214), .Q(fsm5_cnt
		[8]));
	notech_mux2 i_19134(.S(\nbus_14021[0] ), .A(fsm5_cnt[8]), .B(n_871), .Z(n_14384
		));
	notech_mux2 i_1722744(.S(n_62878), .A(iDaddr[28]), .B(iDaddr_f[28]), .Z(\dir1_0[6] 
		));
	notech_reg pg_fault_reg(.CP(n_62948), .D(n_14390), .CD(n_62214), .Q(pg_fault
		));
	notech_mux2 i_19142(.S(n_15216), .A(pg_fault), .B(n_862), .Z(n_14390));
	notech_mux2 i_1822745(.S(n_62878), .A(iDaddr[29]), .B(iDaddr_f[29]), .Z(\dir1_0[7] 
		));
	notech_reg fsm_reg_0(.CP(n_62948), .D(n_14396), .CD(n_62214), .Q(fsm[0])
		);
	notech_mux2 i_19150(.S(\nbus_14018[0] ), .A(n_62882), .B(n_52541), .Z(n_14396
		));
	notech_mux2 i_1922746(.S(n_62878), .A(iDaddr[30]), .B(iDaddr_f[30]), .Z(\dir1_0[8] 
		));
	notech_reg fsm_reg_1(.CP(n_62948), .D(n_14402), .CD(n_62214), .Q(fsm[1])
		);
	notech_mux2 i_19158(.S(\nbus_14018[0] ), .A(fsm[1]), .B(n_52547), .Z(n_14402
		));
	notech_mux2 i_2022747(.S(n_62878), .A(iDaddr[31]), .B(iDaddr_f[31]), .Z(\dir1_0[9] 
		));
	notech_reg fsm_reg_2(.CP(n_62947), .D(n_14408), .CD(n_62213), .Q(fsm[2])
		);
	notech_mux2 i_19166(.S(\nbus_14018[0] ), .A(fsm[2]), .B(n_52553), .Z(n_14408
		));
	notech_nand3 i_75826(.A(n_61580), .B(n_62878), .C(n_15325), .Z(n_52302)
		);
	notech_reg fsm_reg_3(.CP(n_62947), .D(n_14414), .CD(n_62213), .Q(fsm[3])
		);
	notech_mux2 i_19174(.S(\nbus_14018[0] ), .A(fsm[3]), .B(n_861), .Z(n_14414
		));
	notech_nand3 i_75828(.A(n_61580), .B(n_62878), .C(n_15324), .Z(n_52308)
		);
	notech_reg addr_miss_reg_2(.CP(n_62947), .D(n_14420), .CD(n_62213), .Q(\addr_miss[2] 
		));
	notech_mux2 i_19182(.S(n_853), .A(n_15219), .B(\addr_miss[2] ), .Z(n_14420
		));
	notech_nand3 i_75830(.A(n_61580), .B(n_62876), .C(n_15323), .Z(n_52314)
		);
	notech_reg addr_miss_reg_3(.CP(n_62947), .D(n_14426), .CD(n_62213), .Q(\addr_miss[3] 
		));
	notech_mux2 i_19190(.S(n_853), .A(n_15220), .B(\addr_miss[3] ), .Z(n_14426
		));
	notech_nand3 i_75832(.A(n_61580), .B(n_62876), .C(n_15322), .Z(n_52320)
		);
	notech_reg addr_miss_reg_4(.CP(n_62947), .D(n_14432), .CD(n_62213), .Q(\addr_miss[4] 
		));
	notech_mux2 i_19198(.S(n_853), .A(n_15221), .B(\addr_miss[4] ), .Z(n_14432
		));
	notech_nand3 i_75836(.A(n_61580), .B(n_62876), .C(n_15320), .Z(n_52332)
		);
	notech_reg addr_miss_reg_5(.CP(n_62947), .D(n_14438), .CD(n_62213), .Q(\addr_miss[5] 
		));
	notech_mux2 i_19206(.S(n_853), .A(n_15222), .B(\addr_miss[5] ), .Z(n_14438
		));
	notech_nand3 i_75838(.A(n_61580), .B(n_62876), .C(n_15319), .Z(n_52338)
		);
	notech_reg addr_miss_reg_6(.CP(n_62947), .D(n_14444), .CD(n_62213), .Q(\addr_miss[6] 
		));
	notech_mux2 i_19214(.S(n_853), .A(n_15223), .B(\addr_miss[6] ), .Z(n_14444
		));
	notech_nand3 i_75840(.A(n_61580), .B(n_62876), .C(n_15318), .Z(n_52344)
		);
	notech_reg addr_miss_reg_7(.CP(n_62948), .D(n_14450), .CD(n_62214), .Q(\addr_miss[7] 
		));
	notech_mux2 i_19222(.S(n_853), .A(n_15224), .B(\addr_miss[7] ), .Z(n_14450
		));
	notech_nand3 i_75842(.A(n_61580), .B(n_62876), .C(n_15317), .Z(n_52350)
		);
	notech_reg addr_miss_reg_8(.CP(n_62948), .D(n_14456), .CD(n_62214), .Q(\addr_miss[8] 
		));
	notech_mux2 i_19230(.S(n_853), .A(n_15225), .B(\addr_miss[8] ), .Z(n_14456
		));
	notech_nand3 i_75844(.A(n_61580), .B(n_62878), .C(n_15316), .Z(n_52356)
		);
	notech_reg addr_miss_reg_9(.CP(n_62948), .D(n_14462), .CD(n_62214), .Q(\addr_miss[9] 
		));
	notech_mux2 i_19238(.S(n_853), .A(n_15226), .B(\addr_miss[9] ), .Z(n_14462
		));
	notech_nao3 i_75846(.A(n_62878), .B(n_61580), .C(data_miss[12]), .Z(n_52362
		));
	notech_reg addr_miss_reg_10(.CP(n_62948), .D(n_14468), .CD(n_62214), .Q(\addr_miss[10] 
		));
	notech_mux2 i_19246(.S(n_853), .A(n_15227), .B(\addr_miss[10] ), .Z(n_14468
		));
	notech_nao3 i_75848(.A(n_62878), .B(n_61580), .C(data_miss[13]), .Z(n_52368
		));
	notech_reg addr_miss_reg_11(.CP(n_62947), .D(n_14474), .CD(n_62213), .Q(\addr_miss[11] 
		));
	notech_mux2 i_19254(.S(n_853), .A(n_15228), .B(\addr_miss[11] ), .Z(n_14474
		));
	notech_nao3 i_75850(.A(n_62876), .B(n_61580), .C(data_miss[14]), .Z(n_52374
		));
	notech_reg addr_miss_reg_12(.CP(n_62947), .D(n_14480), .CD(n_62213), .Q(\addr_miss[12] 
		));
	notech_mux2 i_19262(.S(n_853), .A(n_54015), .B(\addr_miss[12] ), .Z(n_14480
		));
	notech_nao3 i_75852(.A(n_62878), .B(n_61580), .C(data_miss[15]), .Z(n_52380
		));
	notech_reg addr_miss_reg_13(.CP(n_62948), .D(n_14486), .CD(n_62214), .Q(\addr_miss[13] 
		));
	notech_mux2 i_19270(.S(n_853), .A(n_54021), .B(\addr_miss[13] ), .Z(n_14486
		));
	notech_nao3 i_75854(.A(n_62873), .B(n_61576), .C(data_miss[16]), .Z(n_52386
		));
	notech_reg addr_miss_reg_14(.CP(n_62952), .D(n_14492), .CD(n_62218), .Q(\addr_miss[14] 
		));
	notech_mux2 i_19278(.S(n_853), .A(n_54027), .B(\addr_miss[14] ), .Z(n_14492
		));
	notech_nao3 i_75856(.A(n_62868), .B(n_61576), .C(data_miss[17]), .Z(n_52392
		));
	notech_reg addr_miss_reg_15(.CP(n_62956), .D(n_14498), .CD(n_62222), .Q(\addr_miss[15] 
		));
	notech_mux2 i_19286(.S(n_853), .A(n_54033), .B(\addr_miss[15] ), .Z(n_14498
		));
	notech_nao3 i_75858(.A(n_62868), .B(n_61576), .C(data_miss[18]), .Z(n_52398
		));
	notech_reg addr_miss_reg_16(.CP(n_62956), .D(n_14504), .CD(n_62222), .Q(\addr_miss[16] 
		));
	notech_mux2 i_19294(.S(n_853), .A(n_54039), .B(\addr_miss[16] ), .Z(n_14504
		));
	notech_nao3 i_75860(.A(n_62868), .B(n_61576), .C(data_miss[19]), .Z(n_52404
		));
	notech_reg addr_miss_reg_17(.CP(n_62956), .D(n_14510), .CD(n_62222), .Q(\addr_miss[17] 
		));
	notech_mux2 i_19302(.S(n_61585), .A(n_54045), .B(\addr_miss[17] ), .Z(n_14510
		));
	notech_nao3 i_75862(.A(n_62866), .B(n_61576), .C(data_miss[20]), .Z(n_52410
		));
	notech_reg addr_miss_reg_18(.CP(n_62956), .D(n_14516), .CD(n_62222), .Q(\addr_miss[18] 
		));
	notech_mux2 i_19310(.S(n_61585), .A(n_54051), .B(\addr_miss[18] ), .Z(n_14516
		));
	notech_nao3 i_75864(.A(n_62866), .B(n_61576), .C(data_miss[21]), .Z(n_52416
		));
	notech_reg addr_miss_reg_19(.CP(n_62956), .D(n_14522), .CD(n_62222), .Q(\addr_miss[19] 
		));
	notech_mux2 i_19318(.S(n_61585), .A(n_54057), .B(\addr_miss[19] ), .Z(n_14522
		));
	notech_nao3 i_75866(.A(n_62868), .B(n_61576), .C(data_miss[22]), .Z(n_52422
		));
	notech_reg addr_miss_reg_20(.CP(n_62956), .D(n_14528), .CD(n_62222), .Q(\addr_miss[20] 
		));
	notech_mux2 i_19326(.S(n_61585), .A(n_54063), .B(\addr_miss[20] ), .Z(n_14528
		));
	notech_nao3 i_75868(.A(n_62868), .B(n_61576), .C(data_miss[23]), .Z(n_52428
		));
	notech_reg addr_miss_reg_21(.CP(n_62956), .D(n_14534), .CD(n_62222), .Q(\addr_miss[21] 
		));
	notech_mux2 i_19334(.S(n_61585), .A(n_54069), .B(\addr_miss[21] ), .Z(n_14534
		));
	notech_nao3 i_75870(.A(n_62868), .B(n_61576), .C(data_miss[24]), .Z(n_52434
		));
	notech_reg addr_miss_reg_22(.CP(n_62956), .D(n_14540), .CD(n_62222), .Q(\addr_miss[22] 
		));
	notech_mux2 i_19342(.S(n_61585), .A(n_54075), .B(\addr_miss[22] ), .Z(n_14540
		));
	notech_nao3 i_75872(.A(n_62868), .B(n_61576), .C(data_miss[25]), .Z(n_52440
		));
	notech_reg addr_miss_reg_23(.CP(n_62956), .D(n_14546), .CD(n_62222), .Q(\addr_miss[23] 
		));
	notech_mux2 i_19350(.S(n_61585), .A(n_54081), .B(\addr_miss[23] ), .Z(n_14546
		));
	notech_nao3 i_75874(.A(n_62868), .B(n_61576), .C(data_miss[26]), .Z(n_52446
		));
	notech_reg addr_miss_reg_24(.CP(n_62956), .D(n_14552), .CD(n_62222), .Q(\addr_miss[24] 
		));
	notech_mux2 i_19358(.S(n_61585), .A(n_54087), .B(\addr_miss[24] ), .Z(n_14552
		));
	notech_nao3 i_75876(.A(n_62868), .B(n_61576), .C(data_miss[27]), .Z(n_52452
		));
	notech_reg addr_miss_reg_25(.CP(n_62956), .D(n_14558), .CD(n_62222), .Q(\addr_miss[25] 
		));
	notech_mux2 i_19366(.S(n_61585), .A(n_54093), .B(\addr_miss[25] ), .Z(n_14558
		));
	notech_nao3 i_75878(.A(n_62866), .B(n_61576), .C(data_miss[28]), .Z(n_52458
		));
	notech_reg addr_miss_reg_26(.CP(n_62956), .D(n_14564), .CD(n_62222), .Q(\addr_miss[26] 
		));
	notech_mux2 i_19374(.S(n_61585), .A(n_54099), .B(\addr_miss[26] ), .Z(n_14564
		));
	notech_nao3 i_75880(.A(n_62866), .B(n_61576), .C(data_miss[29]), .Z(n_52464
		));
	notech_reg addr_miss_reg_27(.CP(n_62956), .D(n_14570), .CD(n_62222), .Q(\addr_miss[27] 
		));
	notech_mux2 i_19382(.S(n_61585), .A(n_54105), .B(\addr_miss[27] ), .Z(n_14570
		));
	notech_nao3 i_75882(.A(n_62866), .B(n_61576), .C(data_miss[30]), .Z(n_52470
		));
	notech_reg addr_miss_reg_28(.CP(n_62956), .D(n_14576), .CD(n_62222), .Q(\addr_miss[28] 
		));
	notech_mux2 i_19390(.S(n_61585), .A(n_54111), .B(\addr_miss[28] ), .Z(n_14576
		));
	notech_nao3 i_75884(.A(n_62866), .B(n_61576), .C(data_miss[31]), .Z(n_52476
		));
	notech_reg addr_miss_reg_29(.CP(n_62952), .D(n_14582), .CD(n_62218), .Q(\addr_miss[29] 
		));
	notech_mux2 i_19398(.S(n_61585), .A(n_54117), .B(\addr_miss[29] ), .Z(n_14582
		));
	notech_nand2 i_75890(.A(n_62866), .B(n_61576), .Z(n_52501));
	notech_reg addr_miss_reg_30(.CP(n_62952), .D(n_14588), .CD(n_62218), .Q(\addr_miss[30] 
		));
	notech_mux2 i_19406(.S(n_61585), .A(n_54123), .B(\addr_miss[30] ), .Z(n_14588
		));
	notech_nand2 i_76130(.A(n_896), .B(n_890), .Z(n_52870));
	notech_reg addr_miss_reg_31(.CP(n_62952), .D(n_14594), .CD(n_62218), .Q(\addr_miss[31] 
		));
	notech_mux2 i_19414(.S(n_61585), .A(n_54129), .B(\addr_miss[31] ), .Z(n_14594
		));
	notech_ao4 i_76020(.A(n_938), .B(n_15325), .C(n_912), .D(n_15335), .Z(n_53955
		));
	notech_reg wrA_reg_2(.CP(n_62952), .D(n_14600), .CD(n_62218), .Q(\wrA[2] 
		));
	notech_mux2 i_19422(.S(n_61133), .A(\wrA[2] ), .B(\addr_miss[2] ), .Z(n_14600
		));
	notech_ao4 i_76023(.A(n_938), .B(n_15324), .C(n_912), .D(n_15334), .Z(n_53961
		));
	notech_reg wrA_reg_3(.CP(n_62952), .D(n_14606), .CD(n_62218), .Q(\wrA[3] 
		));
	notech_mux2 i_19430(.S(n_61133), .A(\wrA[3] ), .B(\addr_miss[3] ), .Z(n_14606
		));
	notech_ao4 i_76026(.A(n_938), .B(n_15323), .C(n_912), .D(n_15333), .Z(n_53967
		));
	notech_reg wrA_reg_4(.CP(n_62952), .D(n_14612), .CD(n_62218), .Q(\wrA[4] 
		));
	notech_mux2 i_19438(.S(n_61133), .A(\wrA[4] ), .B(\addr_miss[4] ), .Z(n_14612
		));
	notech_ao4 i_76029(.A(n_938), .B(n_15322), .C(n_912), .D(n_15332), .Z(n_53973
		));
	notech_reg wrA_reg_5(.CP(n_62952), .D(n_14618), .CD(n_62218), .Q(\wrA[5] 
		));
	notech_mux2 i_19446(.S(n_61133), .A(\wrA[5] ), .B(\addr_miss[5] ), .Z(n_14618
		));
	notech_ao4 i_76032(.A(n_938), .B(n_15321), .C(n_912), .D(n_15331), .Z(n_53979
		));
	notech_reg wrA_reg_6(.CP(n_62952), .D(n_14624), .CD(n_62218), .Q(\wrA[6] 
		));
	notech_mux2 i_19454(.S(n_61133), .A(\wrA[6] ), .B(\addr_miss[6] ), .Z(n_14624
		));
	notech_ao4 i_76035(.A(n_938), .B(n_15320), .C(n_912), .D(n_15330), .Z(n_53985
		));
	notech_reg wrA_reg_7(.CP(n_62952), .D(n_14630), .CD(n_62218), .Q(\wrA[7] 
		));
	notech_mux2 i_19462(.S(n_61133), .A(\wrA[7] ), .B(\addr_miss[7] ), .Z(n_14630
		));
	notech_ao4 i_76038(.A(n_938), .B(n_15319), .C(n_912), .D(n_15329), .Z(n_53991
		));
	notech_reg wrA_reg_8(.CP(n_62952), .D(n_14636), .CD(n_62218), .Q(\wrA[8] 
		));
	notech_mux2 i_19470(.S(n_61133), .A(\wrA[8] ), .B(\addr_miss[8] ), .Z(n_14636
		));
	notech_ao4 i_76041(.A(n_938), .B(n_15318), .C(n_912), .D(n_15328), .Z(n_53997
		));
	notech_reg wrA_reg_9(.CP(n_62952), .D(n_14642), .CD(n_62218), .Q(\wrA[9] 
		));
	notech_mux2 i_19478(.S(n_61133), .A(\wrA[9] ), .B(\addr_miss[9] ), .Z(n_14642
		));
	notech_ao4 i_76044(.A(n_938), .B(n_15317), .C(n_912), .D(n_15327), .Z(n_54003
		));
	notech_reg wrA_reg_10(.CP(n_62952), .D(n_14648), .CD(n_62218), .Q(\wrA[10] 
		));
	notech_mux2 i_19486(.S(n_61133), .A(\wrA[10] ), .B(\addr_miss[10] ), .Z(n_14648
		));
	notech_ao4 i_76047(.A(n_938), .B(n_15316), .C(n_912), .D(n_15326), .Z(n_54009
		));
	notech_reg wrA_reg_11(.CP(n_62952), .D(n_14654), .CD(n_62218), .Q(\wrA[11] 
		));
	notech_mux2 i_19494(.S(n_61133), .A(\wrA[11] ), .B(\addr_miss[11] ), .Z(n_14654
		));
	notech_nand2 i_76050(.A(n_970), .B(n_424), .Z(n_54015));
	notech_reg wrA_reg_12(.CP(n_62952), .D(n_14660), .CD(n_62218), .Q(\wrA[12] 
		));
	notech_mux2 i_19502(.S(n_61133), .A(\wrA[12] ), .B(\addr_miss[12] ), .Z(n_14660
		));
	notech_nand2 i_76053(.A(n_969), .B(n_425), .Z(n_54021));
	notech_reg wrA_reg_13(.CP(n_62952), .D(n_14666), .CD(n_62218), .Q(\wrA[13] 
		));
	notech_mux2 i_19510(.S(n_61133), .A(\wrA[13] ), .B(\addr_miss[13] ), .Z(n_14666
		));
	notech_nand2 i_76056(.A(n_968), .B(n_426), .Z(n_54027));
	notech_reg wrA_reg_14(.CP(n_62938), .D(n_14672), .CD(n_62204), .Q(\wrA[14] 
		));
	notech_mux2 i_19518(.S(n_61133), .A(\wrA[14] ), .B(\addr_miss[14] ), .Z(n_14672
		));
	notech_nand2 i_76059(.A(n_967), .B(n_427), .Z(n_54033));
	notech_reg wrA_reg_15(.CP(n_62938), .D(n_14678), .CD(n_62204), .Q(\wrA[15] 
		));
	notech_mux2 i_19526(.S(n_61133), .A(\wrA[15] ), .B(\addr_miss[15] ), .Z(n_14678
		));
	notech_nand2 i_76062(.A(n_966), .B(n_428), .Z(n_54039));
	notech_reg wrA_reg_16(.CP(n_62938), .D(n_14684), .CD(n_62204), .Q(\wrA[16] 
		));
	notech_mux2 i_19534(.S(n_61133), .A(\wrA[16] ), .B(\addr_miss[16] ), .Z(n_14684
		));
	notech_nand2 i_76065(.A(n_965), .B(n_429), .Z(n_54045));
	notech_reg wrA_reg_17(.CP(n_62938), .D(n_14690), .CD(n_62204), .Q(\wrA[17] 
		));
	notech_mux2 i_19542(.S(n_61133), .A(\wrA[17] ), .B(\addr_miss[17] ), .Z(n_14690
		));
	notech_nand2 i_76068(.A(n_964), .B(n_430), .Z(n_54051));
	notech_reg wrA_reg_18(.CP(n_62938), .D(n_14696), .CD(n_62204), .Q(\wrA[18] 
		));
	notech_mux2 i_19550(.S(n_61133), .A(\wrA[18] ), .B(\addr_miss[18] ), .Z(n_14696
		));
	notech_nand2 i_76071(.A(n_963), .B(n_431), .Z(n_54057));
	notech_reg wrA_reg_19(.CP(n_62938), .D(n_14702), .CD(n_62204), .Q(\wrA[19] 
		));
	notech_mux2 i_19558(.S(n_61133), .A(\wrA[19] ), .B(\addr_miss[19] ), .Z(n_14702
		));
	notech_nand2 i_76074(.A(n_962), .B(n_432), .Z(n_54063));
	notech_reg wrA_reg_20(.CP(n_62938), .D(n_14708), .CD(n_62204), .Q(\wrA[20] 
		));
	notech_mux2 i_19566(.S(n_61133), .A(\wrA[20] ), .B(\addr_miss[20] ), .Z(n_14708
		));
	notech_nand2 i_76077(.A(n_961), .B(n_433), .Z(n_54069));
	notech_reg wrA_reg_21(.CP(n_62938), .D(n_14714), .CD(n_62204), .Q(\wrA[21] 
		));
	notech_mux2 i_19574(.S(n_61128), .A(\wrA[21] ), .B(\addr_miss[21] ), .Z(n_14714
		));
	notech_nand2 i_76080(.A(n_960), .B(n_434), .Z(n_54075));
	notech_reg wrA_reg_22(.CP(n_62938), .D(n_14720), .CD(n_62204), .Q(\wrA[22] 
		));
	notech_mux2 i_19582(.S(n_61128), .A(\wrA[22] ), .B(\addr_miss[22] ), .Z(n_14720
		));
	notech_nand2 i_76083(.A(n_959), .B(n_435), .Z(n_54081));
	notech_reg wrA_reg_23(.CP(n_62938), .D(n_14726), .CD(n_62204), .Q(\wrA[23] 
		));
	notech_mux2 i_19590(.S(n_61128), .A(\wrA[23] ), .B(\addr_miss[23] ), .Z(n_14726
		));
	notech_nand2 i_76086(.A(n_958), .B(n_436), .Z(n_54087));
	notech_reg wrA_reg_24(.CP(n_62938), .D(n_14732), .CD(n_62204), .Q(\wrA[24] 
		));
	notech_mux2 i_19598(.S(n_61128), .A(\wrA[24] ), .B(\addr_miss[24] ), .Z(n_14732
		));
	notech_nand2 i_76089(.A(n_957), .B(n_437), .Z(n_54093));
	notech_reg wrA_reg_25(.CP(n_62938), .D(n_14738), .CD(n_62204), .Q(\wrA[25] 
		));
	notech_mux2 i_19606(.S(n_61128), .A(\wrA[25] ), .B(\addr_miss[25] ), .Z(n_14738
		));
	notech_nand2 i_76092(.A(n_956), .B(n_438), .Z(n_54099));
	notech_reg wrA_reg_26(.CP(n_62938), .D(n_14744), .CD(n_62204), .Q(\wrA[26] 
		));
	notech_mux2 i_19614(.S(n_61128), .A(\wrA[26] ), .B(\addr_miss[26] ), .Z(n_14744
		));
	notech_nand2 i_76095(.A(n_955), .B(n_439), .Z(n_54105));
	notech_reg wrA_reg_27(.CP(n_62938), .D(n_14750), .CD(n_62204), .Q(\wrA[27] 
		));
	notech_mux2 i_19622(.S(n_61128), .A(\wrA[27] ), .B(\addr_miss[27] ), .Z(n_14750
		));
	notech_nand2 i_76098(.A(n_954), .B(n_440), .Z(n_54111));
	notech_reg wrA_reg_28(.CP(n_62938), .D(n_14756), .CD(n_62204), .Q(\wrA[28] 
		));
	notech_mux2 i_19630(.S(n_61128), .A(\wrA[28] ), .B(\addr_miss[28] ), .Z(n_14756
		));
	notech_nand2 i_76101(.A(n_953), .B(n_441), .Z(n_54117));
	notech_reg wrA_reg_29(.CP(n_62937), .D(n_14762), .CD(n_62203), .Q(\wrA[29] 
		));
	notech_mux2 i_19638(.S(n_61128), .A(\wrA[29] ), .B(\addr_miss[29] ), .Z(n_14762
		));
	notech_nand2 i_76104(.A(n_952), .B(n_442), .Z(n_54123));
	notech_reg wrA_reg_30(.CP(n_62937), .D(n_14768), .CD(n_62203), .Q(\wrA[30] 
		));
	notech_mux2 i_19646(.S(n_61128), .A(\wrA[30] ), .B(\addr_miss[30] ), .Z(n_14768
		));
	notech_nand2 i_76107(.A(n_951), .B(n_443), .Z(n_54129));
	notech_reg wrA_reg_31(.CP(n_62937), .D(n_14774), .CD(n_62203), .Q(\wrA[31] 
		));
	notech_mux2 i_19654(.S(n_61128), .A(\wrA[31] ), .B(\addr_miss[31] ), .Z(n_14774
		));
	notech_ao4 i_76486(.A(n_912), .B(n_15143), .C(n_896), .D(\nnx_tab2[0] ),
		 .Z(n_54839));
	notech_reg wrD_reg_0(.CP(n_62937), .D(n_14780), .CD(n_62203), .Q(\wrD[0] 
		));
	notech_mux2 i_19662(.S(n_61128), .A(\wrD[0] ), .B(n_52870), .Z(n_14780)
		);
	notech_ao4 i_76489(.A(n_912), .B(n_15145), .C(n_896), .D(n_499), .Z(n_54845
		));
	notech_reg wrD_reg_1(.CP(n_62937), .D(n_14786), .CD(n_62203), .Q(\wrD[1] 
		));
	notech_mux2 i_19670(.S(n_61133), .A(\wrD[1] ), .B(data_miss[1]), .Z(n_14786
		));
	notech_ao4 i_76500(.A(n_896), .B(n_15138), .C(n_487), .D(n_916), .Z(n_52255
		));
	notech_reg wrD_reg_2(.CP(n_62937), .D(n_14792), .CD(n_62203), .Q(\wrD[2] 
		));
	notech_mux2 i_19678(.S(n_61128), .A(\wrD[2] ), .B(data_miss[2]), .Z(n_14792
		));
	notech_ao4 i_76503(.A(n_896), .B(n_15140), .C(n_492), .D(n_917), .Z(n_52261
		));
	notech_reg wrD_reg_3(.CP(n_62937), .D(n_14798), .CD(n_62203), .Q(\wrD[3] 
		));
	notech_mux2 i_19686(.S(n_61128), .A(\wrD[3] ), .B(data_miss[3]), .Z(n_14798
		));
	notech_nand3 i_76643(.A(n_890), .B(n_62866), .C(n_15335), .Z(n_52574));
	notech_reg wrD_reg_4(.CP(n_62937), .D(n_14804), .CD(n_62203), .Q(\wrD[4] 
		));
	notech_mux2 i_19694(.S(n_61128), .A(\wrD[4] ), .B(data_miss[4]), .Z(n_14804
		));
	notech_nand3 i_76645(.A(n_890), .B(n_62866), .C(n_15334), .Z(n_52580));
	notech_reg wrD_reg_5(.CP(n_62937), .D(n_14810), .CD(n_62203), .Q(\wrD[5] 
		));
	notech_mux2 i_19702(.S(n_61128), .A(\wrD[5] ), .B(n_52870), .Z(n_14810)
		);
	notech_nand3 i_76647(.A(n_890), .B(n_62866), .C(n_15333), .Z(n_52586));
	notech_reg wrD_reg_6(.CP(n_62937), .D(n_14816), .CD(n_62203), .Q(\wrD[6] 
		));
	notech_mux2 i_19710(.S(n_61128), .A(\wrD[6] ), .B(data_miss[6]), .Z(n_14816
		));
	notech_nand3 i_76649(.A(n_890), .B(n_62866), .C(n_15332), .Z(n_52592));
	notech_reg wrD_reg_7(.CP(n_62937), .D(n_14822), .CD(n_62203), .Q(\wrD[7] 
		));
	notech_mux2 i_19718(.S(n_61128), .A(\wrD[7] ), .B(data_miss[7]), .Z(n_14822
		));
	notech_nand3 i_76653(.A(n_890), .B(n_62866), .C(n_15330), .Z(n_52604));
	notech_reg req_miss_reg(.CP(n_62937), .D(n_14828), .CD(n_62203), .Q(req_miss
		));
	notech_mux2 i_19726(.S(n_15263), .A(req_miss), .B(n_52519), .Z(n_14828)
		);
	notech_nand3 i_76655(.A(n_890), .B(n_62866), .C(n_15329), .Z(n_52610));
	notech_reg cr2_reg_0(.CP(n_62937), .D(n_14834), .CD(n_62203), .Q(cr2[0])
		);
	notech_mux2 i_19734(.S(n_808), .A(iDaddr_f[0]), .B(cr2[0]), .Z(n_14834)
		);
	notech_nand3 i_76657(.A(n_890), .B(n_62866), .C(n_15328), .Z(n_52616));
	notech_reg cr2_reg_1(.CP(n_62937), .D(n_14840), .CD(n_62203), .Q(cr2[1])
		);
	notech_mux2 i_19742(.S(n_808), .A(iDaddr_f[1]), .B(cr2[1]), .Z(n_14840)
		);
	notech_nand3 i_76659(.A(n_890), .B(n_62871), .C(n_15327), .Z(n_52622));
	notech_reg cr2_reg_2(.CP(n_62938), .D(n_14846), .CD(n_62204), .Q(cr2[2])
		);
	notech_mux2 i_19750(.S(n_808), .A(iDaddr_f[2]), .B(cr2[2]), .Z(n_14846)
		);
	notech_nand3 i_76661(.A(n_890), .B(n_62871), .C(n_15326), .Z(n_52628));
	notech_reg cr2_reg_3(.CP(n_62943), .D(n_14852), .CD(n_62209), .Q(cr2[3])
		);
	notech_mux2 i_19758(.S(n_808), .A(iDaddr_f[3]), .B(cr2[3]), .Z(n_14852)
		);
	notech_nao3 i_76663(.A(n_890), .B(n_62871), .C(data_miss[12]), .Z(n_52634
		));
	notech_reg cr2_reg_4(.CP(n_62947), .D(n_14858), .CD(n_62213), .Q(cr2[4])
		);
	notech_mux2 i_19766(.S(n_808), .A(iDaddr_f[4]), .B(cr2[4]), .Z(n_14858)
		);
	notech_nao3 i_76665(.A(n_890), .B(n_62871), .C(data_miss[13]), .Z(n_52640
		));
	notech_reg cr2_reg_5(.CP(n_62947), .D(n_14864), .CD(n_62213), .Q(cr2[5])
		);
	notech_mux2 i_19774(.S(n_808), .A(iDaddr_f[5]), .B(cr2[5]), .Z(n_14864)
		);
	notech_nao3 i_76667(.A(n_890), .B(n_62871), .C(data_miss[14]), .Z(n_52646
		));
	notech_reg cr2_reg_6(.CP(n_62943), .D(n_14870), .CD(n_62209), .Q(cr2[6])
		);
	notech_mux2 i_19782(.S(n_808), .A(iDaddr_f[6]), .B(cr2[6]), .Z(n_14870)
		);
	notech_nao3 i_76669(.A(n_890), .B(n_62871), .C(data_miss[15]), .Z(n_52652
		));
	notech_reg cr2_reg_7(.CP(n_62943), .D(n_14876), .CD(n_62209), .Q(cr2[7])
		);
	notech_mux2 i_19790(.S(n_808), .A(iDaddr_f[7]), .B(cr2[7]), .Z(n_14876)
		);
	notech_nao3 i_76671(.A(n_62083), .B(n_62871), .C(data_miss[16]), .Z(n_52658
		));
	notech_reg cr2_reg_8(.CP(n_62943), .D(n_14882), .CD(n_62209), .Q(cr2[8])
		);
	notech_mux2 i_19798(.S(n_808), .A(iDaddr_f[8]), .B(cr2[8]), .Z(n_14882)
		);
	notech_nao3 i_76673(.A(n_62083), .B(n_62873), .C(data_miss[17]), .Z(n_52664
		));
	notech_reg cr2_reg_9(.CP(n_62943), .D(n_14888), .CD(n_62209), .Q(cr2[9])
		);
	notech_mux2 i_19806(.S(n_808), .A(iDaddr_f[9]), .B(cr2[9]), .Z(n_14888)
		);
	notech_nao3 i_76675(.A(n_62083), .B(n_62871), .C(data_miss[18]), .Z(n_52670
		));
	notech_reg cr2_reg_10(.CP(n_62947), .D(n_14894), .CD(n_62213), .Q(cr2[10
		]));
	notech_mux2 i_19814(.S(n_808), .A(iDaddr_f[10]), .B(cr2[10]), .Z(n_14894
		));
	notech_nao3 i_76677(.A(n_62083), .B(n_62871), .C(data_miss[19]), .Z(n_52676
		));
	notech_reg cr2_reg_11(.CP(n_62947), .D(n_14900), .CD(n_62213), .Q(cr2[11
		]));
	notech_mux2 i_19822(.S(n_808), .A(iDaddr_f[11]), .B(cr2[11]), .Z(n_14900
		));
	notech_nao3 i_76679(.A(n_62083), .B(n_62871), .C(data_miss[20]), .Z(n_52682
		));
	notech_reg cr2_reg_12(.CP(n_62947), .D(n_14906), .CD(n_62213), .Q(cr2[12
		]));
	notech_mux2 i_19830(.S(n_808), .A(iDaddr_f[12]), .B(cr2[12]), .Z(n_14906
		));
	notech_nao3 i_76681(.A(n_62083), .B(n_62871), .C(data_miss[21]), .Z(n_52688
		));
	notech_reg cr2_reg_13(.CP(n_62947), .D(n_14912), .CD(n_62213), .Q(cr2[13
		]));
	notech_mux2 i_19838(.S(n_808), .A(iDaddr_f[13]), .B(cr2[13]), .Z(n_14912
		));
	notech_nao3 i_76683(.A(n_62083), .B(n_62868), .C(data_miss[22]), .Z(n_52694
		));
	notech_reg cr2_reg_14(.CP(n_62947), .D(n_14918), .CD(n_62213), .Q(cr2[14
		]));
	notech_mux2 i_19846(.S(n_808), .A(iDaddr_f[14]), .B(cr2[14]), .Z(n_14918
		));
	notech_nao3 i_76685(.A(n_62083), .B(n_62868), .C(data_miss[23]), .Z(n_52700
		));
	notech_reg cr2_reg_15(.CP(n_62947), .D(n_14924), .CD(n_62213), .Q(cr2[15
		]));
	notech_mux2 i_19854(.S(n_808), .A(iDaddr_f[15]), .B(cr2[15]), .Z(n_14924
		));
	notech_nao3 i_76687(.A(n_62083), .B(n_62868), .C(data_miss[24]), .Z(n_52706
		));
	notech_reg cr2_reg_16(.CP(n_62947), .D(n_14930), .CD(n_62213), .Q(cr2[16
		]));
	notech_mux2 i_19862(.S(n_55506), .A(iDaddr_f[16]), .B(cr2[16]), .Z(n_14930
		));
	notech_nao3 i_76689(.A(n_62083), .B(n_62868), .C(data_miss[25]), .Z(n_52712
		));
	notech_reg cr2_reg_17(.CP(n_62943), .D(n_14936), .CD(n_62209), .Q(cr2[17
		]));
	notech_mux2 i_19870(.S(n_55506), .A(iDaddr_f[17]), .B(cr2[17]), .Z(n_14936
		));
	notech_nao3 i_76691(.A(n_62083), .B(n_62868), .C(data_miss[26]), .Z(n_52718
		));
	notech_reg cr2_reg_18(.CP(n_62943), .D(n_14942), .CD(n_62209), .Q(cr2[18
		]));
	notech_mux2 i_19878(.S(n_55506), .A(iDaddr_f[18]), .B(cr2[18]), .Z(n_14942
		));
	notech_nao3 i_76693(.A(n_890), .B(n_62868), .C(data_miss[27]), .Z(n_52724
		));
	notech_reg cr2_reg_19(.CP(n_62943), .D(n_14948), .CD(n_62209), .Q(cr2[19
		]));
	notech_mux2 i_19886(.S(n_55506), .A(iDaddr_f[19]), .B(cr2[19]), .Z(n_14948
		));
	notech_nao3 i_76695(.A(n_62083), .B(n_62871), .C(data_miss[28]), .Z(n_52730
		));
	notech_reg cr2_reg_20(.CP(n_62943), .D(n_14954), .CD(n_62209), .Q(cr2[20
		]));
	notech_mux2 i_19894(.S(n_55506), .A(iDaddr_f[20]), .B(cr2[20]), .Z(n_14954
		));
	notech_nao3 i_76697(.A(n_62083), .B(n_62871), .C(data_miss[29]), .Z(n_52736
		));
	notech_reg cr2_reg_21(.CP(n_62943), .D(n_14960), .CD(n_62209), .Q(cr2[21
		]));
	notech_mux2 i_19902(.S(n_55506), .A(iDaddr_f[21]), .B(cr2[21]), .Z(n_14960
		));
	notech_nao3 i_76699(.A(n_62083), .B(n_62871), .C(data_miss[30]), .Z(n_52742
		));
	notech_reg cr2_reg_22(.CP(n_62938), .D(n_14966), .CD(n_62204), .Q(cr2[22
		]));
	notech_mux2 i_19910(.S(n_55506), .A(iDaddr_f[22]), .B(cr2[22]), .Z(n_14966
		));
	notech_nao3 i_76701(.A(n_62083), .B(n_62871), .C(data_miss[31]), .Z(n_52748
		));
	notech_reg cr2_reg_23(.CP(n_62938), .D(n_14972), .CD(n_62204), .Q(cr2[23
		]));
	notech_mux2 i_19918(.S(n_55506), .A(iDaddr_f[23]), .B(cr2[23]), .Z(n_14972
		));
	notech_nand2 i_76707(.A(n_62083), .B(n_62871), .Z(n_52772));
	notech_reg cr2_reg_24(.CP(n_62943), .D(n_14978), .CD(n_62209), .Q(cr2[24
		]));
	notech_mux2 i_19926(.S(n_55506), .A(iDaddr_f[24]), .B(cr2[24]), .Z(n_14978
		));
	notech_ao4 i_76715(.A(n_912), .B(n_15193), .C(n_896), .D(\nnx_tab1[0] ),
		 .Z(n_52019));
	notech_reg cr2_reg_25(.CP(n_62943), .D(n_14984), .CD(n_62209), .Q(cr2[25
		]));
	notech_mux2 i_19934(.S(n_55506), .A(iDaddr_f[25]), .B(cr2[25]), .Z(n_14984
		));
	notech_ao4 i_76718(.A(n_912), .B(n_15195), .C(n_896), .D(n_478), .Z(n_52025
		));
	notech_reg cr2_reg_26(.CP(n_62943), .D(n_14990), .CD(n_62209), .Q(cr2[26
		]));
	notech_mux2 i_19942(.S(n_55506), .A(iDaddr_f[26]), .B(cr2[26]), .Z(n_14990
		));
	notech_ao4 i_76725(.A(n_896), .B(n_15188), .C(n_466), .D(n_926), .Z(n_52789
		));
	notech_reg cr2_reg_27(.CP(n_62943), .D(n_14996), .CD(n_62209), .Q(cr2[27
		]));
	notech_mux2 i_19950(.S(n_55506), .A(iDaddr_f[27]), .B(cr2[27]), .Z(n_14996
		));
	notech_ao4 i_76728(.A(n_896), .B(n_15190), .C(n_471), .D(n_927), .Z(n_52795
		));
	notech_reg cr2_reg_28(.CP(n_62943), .D(n_15002), .CD(n_62209), .Q(cr2[28
		]));
	notech_mux2 i_19958(.S(n_55506), .A(iDaddr_f[28]), .B(cr2[28]), .Z(n_15002
		));
	notech_nand3 i_43(.A(n_912), .B(n_935), .C(n_858), .Z(n_52553));
	notech_reg cr2_reg_29(.CP(n_62943), .D(n_15008), .CD(n_62209), .Q(cr2[29
		]));
	notech_mux2 i_19966(.S(n_55506), .A(iDaddr_f[29]), .B(cr2[29]), .Z(n_15008
		));
	notech_nand3 i_42(.A(n_938), .B(n_855), .C(n_937), .Z(n_52547));
	notech_reg cr2_reg_30(.CP(n_62943), .D(n_15014), .CD(n_62209), .Q(cr2[30
		]));
	notech_mux2 i_19974(.S(n_55506), .A(iDaddr_f[30]), .B(cr2[30]), .Z(n_15014
		));
	notech_mux2 i_41(.S(n_62882), .A(n_447), .B(n_445), .Z(n_52541));
	notech_reg cr2_reg_31(.CP(n_62943), .D(n_15020), .CD(n_62209), .Q(cr2[31
		]));
	notech_mux2 i_19982(.S(n_55506), .A(iDaddr_f[31]), .B(cr2[31]), .Z(n_15020
		));
	notech_inv i_21464(.A(n_985), .Z(n_15026));
	notech_inv i_21465(.A(n_459), .Z(n_15027));
	notech_inv i_21466(.A(n_901), .Z(n_15028));
	notech_inv i_21467(.A(n_889), .Z(n_15029));
	notech_inv i_21468(.A(n_883), .Z(n_15030));
	notech_inv i_21469(.A(\dir1[10] ), .Z(n_15031));
	notech_inv i_21470(.A(\dir1[11] ), .Z(n_15032));
	notech_inv i_21471(.A(\dir1[12] ), .Z(n_15033));
	notech_inv i_21472(.A(\dir1[13] ), .Z(n_15034));
	notech_inv i_21473(.A(\dir1[14] ), .Z(n_15035));
	notech_inv i_21474(.A(\dir1[15] ), .Z(n_15036));
	notech_inv i_21475(.A(\dir1[16] ), .Z(n_15037));
	notech_inv i_21476(.A(\dir1[17] ), .Z(n_15038));
	notech_inv i_21477(.A(\dir1[18] ), .Z(n_15039));
	notech_inv i_21478(.A(\dir1[19] ), .Z(n_15040));
	notech_inv i_21479(.A(\dir1[20] ), .Z(n_15041));
	notech_inv i_21480(.A(\dir1[21] ), .Z(n_15042));
	notech_inv i_21481(.A(\dir1[22] ), .Z(n_15043));
	notech_inv i_21482(.A(\dir1[23] ), .Z(n_15044));
	notech_inv i_21483(.A(\dir1[24] ), .Z(n_15045));
	notech_inv i_21484(.A(\dir1[25] ), .Z(n_15046));
	notech_inv i_21485(.A(\dir1[26] ), .Z(n_15047));
	notech_inv i_21486(.A(\dir1[27] ), .Z(n_15048));
	notech_inv i_21487(.A(\dir1[28] ), .Z(n_15049));
	notech_inv i_21488(.A(\dir1[29] ), .Z(n_15050));
	notech_inv i_21489(.A(\dir2[10] ), .Z(n_15051));
	notech_inv i_21490(.A(\dir2[11] ), .Z(n_15052));
	notech_inv i_21491(.A(\dir2[12] ), .Z(n_15053));
	notech_inv i_21492(.A(\dir2[13] ), .Z(n_15054));
	notech_inv i_21493(.A(\dir2[14] ), .Z(n_15055));
	notech_inv i_21494(.A(\dir2[15] ), .Z(n_15056));
	notech_inv i_21495(.A(\dir2[16] ), .Z(n_15057));
	notech_inv i_21496(.A(\dir2[17] ), .Z(n_15058));
	notech_inv i_21497(.A(\dir2[18] ), .Z(n_15059));
	notech_inv i_21498(.A(\dir2[19] ), .Z(n_15060));
	notech_inv i_21499(.A(\dir2[20] ), .Z(n_15061));
	notech_inv i_21500(.A(\dir2[21] ), .Z(n_15062));
	notech_inv i_21501(.A(\dir2[22] ), .Z(n_15063));
	notech_inv i_21502(.A(\dir2[23] ), .Z(n_15064));
	notech_inv i_21503(.A(\dir2[24] ), .Z(n_15065));
	notech_inv i_21504(.A(\dir2[25] ), .Z(n_15066));
	notech_inv i_21505(.A(\dir2[26] ), .Z(n_15067));
	notech_inv i_21506(.A(\dir2[27] ), .Z(n_15068));
	notech_inv i_21507(.A(\dir2[28] ), .Z(n_15069));
	notech_inv i_21508(.A(\dir2[29] ), .Z(n_15070));
	notech_inv i_21509(.A(n_476), .Z(n_15071));
	notech_inv i_21510(.A(\tab21[10] ), .Z(n_15072));
	notech_inv i_21511(.A(\tab21[11] ), .Z(n_15073));
	notech_inv i_21512(.A(\tab21[12] ), .Z(n_15074));
	notech_inv i_21513(.A(\tab21[13] ), .Z(n_15075));
	notech_inv i_21514(.A(\tab21[14] ), .Z(n_15076));
	notech_inv i_21515(.A(\tab21[15] ), .Z(n_15077));
	notech_inv i_21516(.A(\tab21[16] ), .Z(n_15078));
	notech_inv i_21517(.A(\tab21[17] ), .Z(n_15079));
	notech_inv i_21518(.A(\tab21[18] ), .Z(n_15080));
	notech_inv i_21519(.A(\tab21[19] ), .Z(n_15081));
	notech_inv i_21520(.A(\tab21[20] ), .Z(n_15082));
	notech_inv i_21521(.A(\tab21[21] ), .Z(n_15083));
	notech_inv i_21522(.A(\tab21[22] ), .Z(n_15084));
	notech_inv i_21523(.A(\tab21[23] ), .Z(n_15085));
	notech_inv i_21524(.A(n_497), .Z(n_15086));
	notech_inv i_21525(.A(\tab21[24] ), .Z(n_15087));
	notech_inv i_21526(.A(\tab21[25] ), .Z(n_15088));
	notech_inv i_21527(.A(\tab21[26] ), .Z(n_15089));
	notech_inv i_21528(.A(\tab21[27] ), .Z(n_15090));
	notech_inv i_21529(.A(\tab21[28] ), .Z(n_15091));
	notech_inv i_21530(.A(\tab21[29] ), .Z(n_15092));
	notech_inv i_21531(.A(\tab23[10] ), .Z(n_15093));
	notech_inv i_21532(.A(\tab23[11] ), .Z(n_15094));
	notech_inv i_21533(.A(\tab23[12] ), .Z(n_15095));
	notech_inv i_21534(.A(\tab23[13] ), .Z(n_15096));
	notech_inv i_21535(.A(\tab23[14] ), .Z(n_15097));
	notech_inv i_21536(.A(\tab23[15] ), .Z(n_15098));
	notech_inv i_21537(.A(\tab23[16] ), .Z(n_15099));
	notech_inv i_21538(.A(n_553), .Z(n_15100));
	notech_inv i_21539(.A(\tab23[17] ), .Z(n_15101));
	notech_inv i_21540(.A(\tab23[18] ), .Z(n_15102));
	notech_inv i_21541(.A(\tab23[19] ), .Z(n_15103));
	notech_inv i_21542(.A(\tab23[20] ), .Z(n_15104));
	notech_inv i_21543(.A(n_557), .Z(n_15105));
	notech_inv i_21544(.A(\tab23[21] ), .Z(n_15106));
	notech_inv i_21545(.A(\tab23[22] ), .Z(n_15107));
	notech_inv i_21546(.A(n_559), .Z(n_15108));
	notech_inv i_21547(.A(\tab23[23] ), .Z(n_15109));
	notech_inv i_21548(.A(\tab23[24] ), .Z(n_15110));
	notech_inv i_21549(.A(\tab23[25] ), .Z(n_15111));
	notech_inv i_21550(.A(\tab23[26] ), .Z(n_15112));
	notech_inv i_21551(.A(\tab23[27] ), .Z(n_15113));
	notech_inv i_21552(.A(\tab23[28] ), .Z(n_15114));
	notech_inv i_21553(.A(\tab23[29] ), .Z(n_15115));
	notech_inv i_21554(.A(hit_adr23), .Z(n_15116));
	notech_inv i_21555(.A(\tab24[10] ), .Z(n_15117));
	notech_inv i_21556(.A(\tab24[11] ), .Z(n_15118));
	notech_inv i_21557(.A(\tab24[12] ), .Z(n_15119));
	notech_inv i_21558(.A(\tab24[13] ), .Z(n_15120));
	notech_inv i_21559(.A(\tab24[14] ), .Z(n_15121));
	notech_inv i_21560(.A(\tab24[15] ), .Z(n_15122));
	notech_inv i_21561(.A(\tab24[16] ), .Z(n_15123));
	notech_inv i_21562(.A(\tab24[17] ), .Z(n_15124));
	notech_inv i_21563(.A(\tab24[18] ), .Z(n_15125));
	notech_inv i_21564(.A(\tab24[19] ), .Z(n_15126));
	notech_inv i_21565(.A(\tab24[20] ), .Z(n_15127));
	notech_inv i_21566(.A(\tab24[21] ), .Z(n_15128));
	notech_inv i_21567(.A(\tab24[22] ), .Z(n_15129));
	notech_inv i_21568(.A(\tab24[23] ), .Z(n_15130));
	notech_inv i_21569(.A(\tab24[24] ), .Z(n_15131));
	notech_inv i_21570(.A(\tab24[25] ), .Z(n_15132));
	notech_inv i_21571(.A(\tab24[26] ), .Z(n_15133));
	notech_inv i_21572(.A(\tab24[27] ), .Z(n_15134));
	notech_inv i_21573(.A(\tab24[28] ), .Z(n_15135));
	notech_inv i_21574(.A(\tab24[29] ), .Z(n_15136));
	notech_inv i_21575(.A(n_54839), .Z(n_15137));
	notech_inv i_21576(.A(\nnx_tab2[0] ), .Z(n_15138));
	notech_inv i_21577(.A(n_54845), .Z(n_15139));
	notech_inv i_21578(.A(\nnx_tab2[1] ), .Z(n_15140));
	notech_inv i_21579(.A(\nbus_14041[0] ), .Z(n_15141));
	notech_inv i_21580(.A(n_52255), .Z(n_15142));
	notech_inv i_21581(.A(\nx_tab2[0] ), .Z(n_15143));
	notech_inv i_21582(.A(n_52261), .Z(n_15144));
	notech_inv i_21583(.A(\nx_tab2[1] ), .Z(n_15145));
	notech_inv i_21584(.A(\tab12[10] ), .Z(n_15146));
	notech_inv i_21585(.A(\tab12[11] ), .Z(n_15147));
	notech_inv i_21586(.A(\tab12[12] ), .Z(n_15148));
	notech_inv i_21587(.A(\tab12[13] ), .Z(n_15149));
	notech_inv i_21588(.A(\tab12[14] ), .Z(n_15150));
	notech_inv i_21589(.A(\tab12[15] ), .Z(n_15151));
	notech_inv i_21590(.A(\tab12[16] ), .Z(n_15152));
	notech_inv i_21591(.A(\tab12[17] ), .Z(n_15153));
	notech_inv i_21592(.A(\tab12[18] ), .Z(n_15154));
	notech_inv i_21593(.A(\tab12[19] ), .Z(n_15155));
	notech_inv i_21594(.A(\tab12[20] ), .Z(n_15156));
	notech_inv i_21595(.A(\tab12[21] ), .Z(n_15157));
	notech_inv i_21596(.A(\tab12[22] ), .Z(n_15158));
	notech_inv i_21597(.A(\tab12[23] ), .Z(n_15159));
	notech_inv i_21598(.A(\tab12[24] ), .Z(n_15160));
	notech_inv i_21599(.A(\tab12[25] ), .Z(n_15161));
	notech_inv i_21600(.A(\tab12[26] ), .Z(n_15162));
	notech_inv i_21601(.A(\tab12[27] ), .Z(n_15163));
	notech_inv i_21602(.A(\tab12[28] ), .Z(n_15164));
	notech_inv i_21603(.A(\tab12[29] ), .Z(n_15165));
	notech_inv i_21604(.A(hit_adr13), .Z(n_15166));
	notech_inv i_21605(.A(\tab14[10] ), .Z(n_15167));
	notech_inv i_21606(.A(\tab14[11] ), .Z(n_15168));
	notech_inv i_21607(.A(\tab14[12] ), .Z(n_15169));
	notech_inv i_21608(.A(\tab14[13] ), .Z(n_15170));
	notech_inv i_21609(.A(\tab14[14] ), .Z(n_15171));
	notech_inv i_21610(.A(\tab14[15] ), .Z(n_15172));
	notech_inv i_21611(.A(\tab14[16] ), .Z(n_15173));
	notech_inv i_21612(.A(\tab14[17] ), .Z(n_15174));
	notech_inv i_21613(.A(\tab14[18] ), .Z(n_15175));
	notech_inv i_21614(.A(\tab14[19] ), .Z(n_15176));
	notech_inv i_21615(.A(\tab14[20] ), .Z(n_15177));
	notech_inv i_21616(.A(\tab14[21] ), .Z(n_15178));
	notech_inv i_21617(.A(\tab14[22] ), .Z(n_15179));
	notech_inv i_21618(.A(\tab14[23] ), .Z(n_15180));
	notech_inv i_21619(.A(\tab14[24] ), .Z(n_15181));
	notech_inv i_21620(.A(\tab14[25] ), .Z(n_15182));
	notech_inv i_21621(.A(\tab14[26] ), .Z(n_15183));
	notech_inv i_21622(.A(\tab14[27] ), .Z(n_15184));
	notech_inv i_21623(.A(\tab14[28] ), .Z(n_15185));
	notech_inv i_21624(.A(\tab14[29] ), .Z(n_15186));
	notech_inv i_21625(.A(n_52019), .Z(n_15187));
	notech_inv i_21626(.A(\nnx_tab1[0] ), .Z(n_15188));
	notech_inv i_21627(.A(n_52025), .Z(n_15189));
	notech_inv i_21628(.A(\nnx_tab1[1] ), .Z(n_15190));
	notech_inv i_21629(.A(\nbus_14014[0] ), .Z(n_15191));
	notech_inv i_21630(.A(n_52789), .Z(n_15192));
	notech_inv i_21631(.A(\nx_tab1[0] ), .Z(n_15193));
	notech_inv i_21632(.A(n_52795), .Z(n_15194));
	notech_inv i_21633(.A(\nx_tab1[1] ), .Z(n_15195));
	notech_inv i_21634(.A(\tab11[10] ), .Z(n_15196));
	notech_inv i_21635(.A(\tab11[11] ), .Z(n_15197));
	notech_inv i_21636(.A(\tab11[12] ), .Z(n_15198));
	notech_inv i_21637(.A(\tab11[13] ), .Z(n_15199));
	notech_inv i_21638(.A(\tab11[14] ), .Z(n_15200));
	notech_inv i_21639(.A(\tab11[15] ), .Z(n_15201));
	notech_inv i_21640(.A(\tab11[16] ), .Z(n_15202));
	notech_inv i_21641(.A(\tab11[17] ), .Z(n_15203));
	notech_inv i_21642(.A(\tab11[18] ), .Z(n_15204));
	notech_inv i_21643(.A(\tab11[19] ), .Z(n_15205));
	notech_inv i_21644(.A(\tab11[20] ), .Z(n_15206));
	notech_inv i_21645(.A(\tab11[21] ), .Z(n_15207));
	notech_inv i_21646(.A(\tab11[22] ), .Z(n_15208));
	notech_inv i_21647(.A(\tab11[23] ), .Z(n_15209));
	notech_inv i_21648(.A(\tab11[24] ), .Z(n_15210));
	notech_inv i_21649(.A(\tab11[25] ), .Z(n_15211));
	notech_inv i_21650(.A(\tab11[26] ), .Z(n_15212));
	notech_inv i_21651(.A(\tab11[27] ), .Z(n_15213));
	notech_inv i_21652(.A(\tab11[28] ), .Z(n_15214));
	notech_inv i_21653(.A(\tab11[29] ), .Z(n_15215));
	notech_inv i_21654(.A(n_52233), .Z(n_15216));
	notech_inv i_21655(.A(n_62882), .Z(n_15217));
	notech_inv i_21656(.A(fsm[3]), .Z(n_15218));
	notech_inv i_21657(.A(n_53955), .Z(n_15219));
	notech_inv i_21658(.A(n_53961), .Z(n_15220));
	notech_inv i_21659(.A(n_53967), .Z(n_15221));
	notech_inv i_21660(.A(n_53973), .Z(n_15222));
	notech_inv i_21661(.A(n_53979), .Z(n_15223));
	notech_inv i_21662(.A(n_53985), .Z(n_15224));
	notech_inv i_21663(.A(n_53991), .Z(n_15225));
	notech_inv i_21664(.A(n_53997), .Z(n_15226));
	notech_inv i_21665(.A(n_54003), .Z(n_15227));
	notech_inv i_21666(.A(n_54009), .Z(n_15228));
	notech_inv i_21667(.A(\addr_miss[2] ), .Z(n_15229));
	notech_inv i_21668(.A(\addr_miss[3] ), .Z(n_15230));
	notech_inv i_21669(.A(\addr_miss[4] ), .Z(n_15231));
	notech_inv i_21670(.A(\addr_miss[5] ), .Z(n_15232));
	notech_inv i_21671(.A(\addr_miss[6] ), .Z(n_15233));
	notech_inv i_21672(.A(\addr_miss[7] ), .Z(n_15234));
	notech_inv i_21673(.A(\addr_miss[8] ), .Z(n_15235));
	notech_inv i_21674(.A(\addr_miss[9] ), .Z(n_15236));
	notech_inv i_21675(.A(\addr_miss[10] ), .Z(n_15237));
	notech_inv i_21676(.A(\addr_miss[11] ), .Z(n_15238));
	notech_inv i_21677(.A(\wrA[12] ), .Z(n_15239));
	notech_inv i_21678(.A(\wrA[13] ), .Z(n_15240));
	notech_inv i_21679(.A(\wrA[14] ), .Z(n_15241));
	notech_inv i_21680(.A(\wrA[15] ), .Z(n_15242));
	notech_inv i_21681(.A(\wrA[16] ), .Z(n_15243));
	notech_inv i_21682(.A(\wrA[17] ), .Z(n_15244));
	notech_inv i_21683(.A(\wrA[18] ), .Z(n_15245));
	notech_inv i_21684(.A(\wrA[19] ), .Z(n_15246));
	notech_inv i_21685(.A(\wrA[20] ), .Z(n_15247));
	notech_inv i_21686(.A(\wrA[21] ), .Z(n_15248));
	notech_inv i_21687(.A(\wrA[22] ), .Z(n_15249));
	notech_inv i_21688(.A(\wrA[23] ), .Z(n_15250));
	notech_inv i_21689(.A(\wrA[24] ), .Z(n_15251));
	notech_inv i_21690(.A(\wrA[25] ), .Z(n_15252));
	notech_inv i_21691(.A(\wrA[26] ), .Z(n_15253));
	notech_inv i_21692(.A(\wrA[27] ), .Z(n_15254));
	notech_inv i_21693(.A(\wrA[28] ), .Z(n_15255));
	notech_inv i_21694(.A(\wrA[29] ), .Z(n_15256));
	notech_inv i_21695(.A(\wrA[30] ), .Z(n_15257));
	notech_inv i_21696(.A(\wrA[31] ), .Z(n_15258));
	notech_inv i_21697(.A(n_52870), .Z(n_15259));
	notech_inv i_21699(.A(n_52519), .Z(n_15261));
	notech_inv i_21700(.A(req_miss), .Z(n_15262));
	notech_inv i_21701(.A(n_52516), .Z(n_15263));
	notech_inv i_21702(.A(addr_phys_31101029), .Z(addr_phys[31]));
	notech_inv i_21703(.A(addr_phys_30101028), .Z(addr_phys[30]));
	notech_inv i_21704(.A(addr_phys_29101027), .Z(addr_phys[29]));
	notech_inv i_21705(.A(addr_phys_28101026), .Z(addr_phys[28]));
	notech_inv i_21706(.A(addr_phys_27101025), .Z(addr_phys[27]));
	notech_inv i_21707(.A(addr_phys_26101024), .Z(addr_phys[26]));
	notech_inv i_21708(.A(addr_phys_25101023), .Z(addr_phys[25]));
	notech_inv i_21709(.A(addr_phys_24101022), .Z(addr_phys[24]));
	notech_inv i_21710(.A(addr_phys_23101021), .Z(addr_phys[23]));
	notech_inv i_21711(.A(addr_phys_22101020), .Z(addr_phys[22]));
	notech_inv i_21712(.A(addr_phys_21101019), .Z(addr_phys[21]));
	notech_inv i_21713(.A(addr_phys_20101018), .Z(addr_phys[20]));
	notech_inv i_21714(.A(addr_phys_19101017), .Z(addr_phys[19]));
	notech_inv i_21715(.A(addr_phys_18101016), .Z(addr_phys[18]));
	notech_inv i_21716(.A(addr_phys_17101015), .Z(addr_phys[17]));
	notech_inv i_21717(.A(addr_phys_16101014), .Z(addr_phys[16]));
	notech_inv i_21718(.A(addr_phys_15101013), .Z(addr_phys[15]));
	notech_inv i_21719(.A(addr_phys_14101012), .Z(addr_phys[14]));
	notech_inv i_21720(.A(addr_phys_13101011), .Z(addr_phys[13]));
	notech_inv i_21721(.A(addr_phys_12101010), .Z(addr_phys[12]));
	notech_inv i_21722(.A(n_61576), .Z(n_15284));
	notech_inv i_21723(.A(iDaddr[2]), .Z(n_15285));
	notech_inv i_21724(.A(iDaddr[3]), .Z(n_15286));
	notech_inv i_21725(.A(iDaddr[4]), .Z(n_15287));
	notech_inv i_21726(.A(iDaddr[5]), .Z(n_15288));
	notech_inv i_21727(.A(iDaddr[6]), .Z(n_15289));
	notech_inv i_21728(.A(iDaddr[7]), .Z(n_15290));
	notech_inv i_21729(.A(iDaddr[8]), .Z(n_15291));
	notech_inv i_21730(.A(iDaddr[9]), .Z(n_15292));
	notech_inv i_21731(.A(iDaddr[10]), .Z(n_15293));
	notech_inv i_21732(.A(iDaddr[11]), .Z(n_15294));
	notech_inv i_21733(.A(iDaddr[12]), .Z(n_15295));
	notech_inv i_21734(.A(iDaddr[13]), .Z(n_15296));
	notech_inv i_21735(.A(iDaddr[14]), .Z(n_15297));
	notech_inv i_21736(.A(iDaddr[15]), .Z(n_15298));
	notech_inv i_21737(.A(iDaddr[16]), .Z(n_15299));
	notech_inv i_21738(.A(iDaddr[17]), .Z(n_15300));
	notech_inv i_21739(.A(iDaddr[18]), .Z(n_15301));
	notech_inv i_21740(.A(iDaddr[19]), .Z(n_15302));
	notech_inv i_21741(.A(iDaddr[20]), .Z(n_15303));
	notech_inv i_21742(.A(iDaddr[21]), .Z(n_15304));
	notech_inv i_21743(.A(iDaddr[22]), .Z(n_15305));
	notech_inv i_21744(.A(iDaddr[23]), .Z(n_15306));
	notech_inv i_21745(.A(iDaddr[24]), .Z(n_15307));
	notech_inv i_21746(.A(iDaddr[25]), .Z(n_15308));
	notech_inv i_21747(.A(iDaddr[26]), .Z(n_15309));
	notech_inv i_21748(.A(iDaddr[27]), .Z(n_15310));
	notech_inv i_21749(.A(iDaddr[28]), .Z(n_15311));
	notech_inv i_21750(.A(iDaddr[29]), .Z(n_15312));
	notech_inv i_21751(.A(iDaddr[30]), .Z(n_15313));
	notech_inv i_21752(.A(iDaddr[31]), .Z(n_15314));
	notech_inv i_21753(.A(n_62831), .Z(owrite_req));
	notech_inv i_21754(.A(\dir1_0[9] ), .Z(n_15316));
	notech_inv i_21755(.A(\dir1_0[8] ), .Z(n_15317));
	notech_inv i_21756(.A(\dir1_0[7] ), .Z(n_15318));
	notech_inv i_21757(.A(\dir1_0[6] ), .Z(n_15319));
	notech_inv i_21758(.A(\dir1_0[5] ), .Z(n_15320));
	notech_inv i_21759(.A(\dir1_0[4] ), .Z(n_15321));
	notech_inv i_21760(.A(\dir1_0[3] ), .Z(n_15322));
	notech_inv i_21761(.A(\dir1_0[2] ), .Z(n_15323));
	notech_inv i_21762(.A(\dir1_0[1] ), .Z(n_15324));
	notech_inv i_21763(.A(\dir1_0[0] ), .Z(n_15325));
	notech_inv i_21764(.A(\tab11_0[9] ), .Z(n_15326));
	notech_inv i_21765(.A(\tab11_0[8] ), .Z(n_15327));
	notech_inv i_21766(.A(\tab11_0[7] ), .Z(n_15328));
	notech_inv i_21767(.A(\tab11_0[6] ), .Z(n_15329));
	notech_inv i_21768(.A(\tab11_0[5] ), .Z(n_15330));
	notech_inv i_21769(.A(\tab11_0[4] ), .Z(n_15331));
	notech_inv i_21770(.A(\tab11_0[3] ), .Z(n_15332));
	notech_inv i_21771(.A(\tab11_0[2] ), .Z(n_15333));
	notech_inv i_21772(.A(\tab11_0[1] ), .Z(n_15334));
	notech_inv i_21773(.A(\tab11_0[0] ), .Z(n_15335));
	notech_inv i_21774(.A(oread_req101009), .Z(oread_req));
	notech_inv i_21775(.A(hit_tab21), .Z(n_15337));
	notech_inv i_21776(.A(hit_tab23), .Z(n_15338));
	notech_inv i_21777(.A(hit_tab12), .Z(n_15339));
	notech_inv i_21778(.A(\hit_dir1[7] ), .Z(n_15340));
	notech_inv i_21779(.A(n_62908), .Z(n_15341));
	notech_inv i_21780(.A(iread_req), .Z(n_15342));
	notech_inv i_21781(.A(hit_dir2), .Z(n_15343));
	notech_inv i_21782(.A(pg_fault), .Z(n_15344));
	cmp14_19 t11(.ina({\tab11[33] , UNCONNECTED_000, UNCONNECTED_001, 
		UNCONNECTED_002, \tab11[9] , \tab11[8] , \tab11[7] , \tab11[6] ,
		 \tab11[5] , \tab11[4] , \tab11[3] , \tab11[2] , \tab11[1] , \tab11[0] 
		}), .inb({UNCONNECTED_003, UNCONNECTED_004, UNCONNECTED_005, 
		UNCONNECTED_006, \tab11_0[9] , \tab11_0[8] , \tab11_0[7] , \tab11_0[6] 
		, \tab11_0[5] , \tab11_0[4] , \tab11_0[3] , \tab11_0[2] , \tab11_0[1] 
		, \tab11_0[0] }), .out(hit_tab11), .out2(hit_add11));
	cmp14_18 t14(.ina({\tab14[33] , UNCONNECTED_007, UNCONNECTED_008, 
		UNCONNECTED_009, \tab14[9] , \tab14[8] , \tab14[7] , \tab14[6] ,
		 \tab14[5] , \tab14[4] , \tab14[3] , \tab14[2] , \tab14[1] , \tab14[0] 
		}), .inb({UNCONNECTED_010, UNCONNECTED_011, UNCONNECTED_012, 
		UNCONNECTED_013, \tab11_0[9] , \tab11_0[8] , \tab11_0[7] , \tab11_0[6] 
		, \tab11_0[5] , \tab11_0[4] , \tab11_0[3] , \tab11_0[2] , \tab11_0[1] 
		, \tab11_0[0] }), .out(hit_tab14), .out2(hit_add14));
	cmp14_17 t13(.ina({\tab13[33] , UNCONNECTED_014, UNCONNECTED_015, 
		UNCONNECTED_016, \tab13[9] , \tab13[8] , \tab13[7] , \tab13[6] ,
		 \tab13[5] , \tab13[4] , \tab13[3] , \tab13[2] , \tab13[1] , \tab13[0] 
		}), .inb({UNCONNECTED_017, UNCONNECTED_018, UNCONNECTED_019, 
		UNCONNECTED_020, \tab11_0[9] , \tab11_0[8] , \tab11_0[7] , \tab11_0[6] 
		, \tab11_0[5] , \tab11_0[4] , \tab11_0[3] , \tab11_0[2] , \tab11_0[1] 
		, \tab11_0[0] }), .out(hit_tab13), .out2(hit_add13));
	cmp14_16 t12(.ina({\tab12[33] , UNCONNECTED_021, UNCONNECTED_022, 
		UNCONNECTED_023, \tab12[9] , \tab12[8] , \tab12[7] , \tab12[6] ,
		 \tab12[5] , \tab12[4] , \tab12[3] , \tab12[2] , \tab12[1] , \tab12[0] 
		}), .inb({UNCONNECTED_024, UNCONNECTED_025, UNCONNECTED_026, 
		UNCONNECTED_027, \tab11_0[9] , \tab11_0[8] , \tab11_0[7] , \tab11_0[6] 
		, \tab11_0[5] , \tab11_0[4] , \tab11_0[3] , \tab11_0[2] , \tab11_0[1] 
		, \tab11_0[0] }), .out(hit_tab12), .out2(hit_add12));
	cmp14_15 t24(.ina({\tab24[33] , UNCONNECTED_028, UNCONNECTED_029, 
		UNCONNECTED_030, \tab24[9] , \tab24[8] , \tab24[7] , \tab24[6] ,
		 \tab24[5] , \tab24[4] , \tab24[3] , \tab24[2] , \tab24[1] , \tab24[0] 
		}), .inb({UNCONNECTED_031, UNCONNECTED_032, UNCONNECTED_033, 
		UNCONNECTED_034, \tab11_0[9] , \tab11_0[8] , \tab11_0[7] , \tab11_0[6] 
		, \tab11_0[5] , \tab11_0[4] , \tab11_0[3] , \tab11_0[2] , \tab11_0[1] 
		, \tab11_0[0] }), .out(hit_tab24), .out2(hit_add24));
	cmp14_14 t23(.ina({\tab23[33] , UNCONNECTED_035, UNCONNECTED_036, 
		UNCONNECTED_037, \tab23[9] , \tab23[8] , \tab23[7] , \tab23[6] ,
		 \tab23[5] , \tab23[4] , \tab23[3] , \tab23[2] , \tab23[1] , \tab23[0] 
		}), .inb({UNCONNECTED_038, UNCONNECTED_039, UNCONNECTED_040, 
		UNCONNECTED_041, \tab11_0[9] , \tab11_0[8] , \tab11_0[7] , \tab11_0[6] 
		, \tab11_0[5] , \tab11_0[4] , \tab11_0[3] , \tab11_0[2] , \tab11_0[1] 
		, \tab11_0[0] }), .out(hit_tab23), .out2(hit_add23));
	cmp14_13 t22(.ina({\tab22[33] , UNCONNECTED_042, UNCONNECTED_043, 
		UNCONNECTED_044, \tab22[9] , \tab22[8] , \tab22[7] , \tab22[6] ,
		 \tab22[5] , \tab22[4] , \tab22[3] , \tab22[2] , \tab22[1] , \tab22[0] 
		}), .inb({UNCONNECTED_045, UNCONNECTED_046, UNCONNECTED_047, 
		UNCONNECTED_048, \tab11_0[9] , \tab11_0[8] , \tab11_0[7] , \tab11_0[6] 
		, \tab11_0[5] , \tab11_0[4] , \tab11_0[3] , \tab11_0[2] , \tab11_0[1] 
		, \tab11_0[0] }), .out(hit_tab22), .out2(hit_add22));
	cmp14_12 t21(.ina({\tab21[33] , UNCONNECTED_049, UNCONNECTED_050, 
		UNCONNECTED_051, \tab21[9] , \tab21[8] , \tab21[7] , \tab21[6] ,
		 \tab21[5] , \tab21[4] , \tab21[3] , \tab21[2] , \tab21[1] , \tab21[0] 
		}), .inb({UNCONNECTED_052, UNCONNECTED_053, UNCONNECTED_054, 
		UNCONNECTED_055, \tab11_0[9] , \tab11_0[8] , \tab11_0[7] , \tab11_0[6] 
		, \tab11_0[5] , \tab11_0[4] , \tab11_0[3] , \tab11_0[2] , \tab11_0[1] 
		, \tab11_0[0] }), .out(hit_tab21), .out2(hit_add21));
	cmp14_11 d2(.ina({\dir2[33] , UNCONNECTED_056, UNCONNECTED_057, 
		UNCONNECTED_058, \dir2[9] , \dir2[8] , \dir2[7] , \dir2[6] , \dir2[5] 
		, \dir2[4] , \dir2[3] , \dir2[2] , \dir2[1] , \dir2[0] }), .inb(
		{UNCONNECTED_059, UNCONNECTED_060, UNCONNECTED_061, 
		UNCONNECTED_062, \dir1_0[9] , \dir1_0[8] , \dir1_0[7] , \dir1_0[6] 
		, \dir1_0[5] , \dir1_0[4] , \dir1_0[3] , \dir1_0[2] , \dir1_0[1] 
		, \dir1_0[0] }), .out(hit_dir2));
	cmp14_10 d1(.ina({\dir1[33] , UNCONNECTED_063, UNCONNECTED_064, 
		UNCONNECTED_065, \dir1[9] , \dir1[8] , \dir1[7] , \dir1[6] , \dir1[5] 
		, \dir1[4] , \dir1[3] , \dir1[2] , \dir1[1] , \dir1[0] }), .inb(
		{UNCONNECTED_066, UNCONNECTED_067, UNCONNECTED_068, 
		UNCONNECTED_069, \dir1_0[9] , \dir1_0[8] , \dir1_0[7] , \dir1_0[6] 
		, \dir1_0[5] , \dir1_0[4] , \dir1_0[3] , \dir1_0[2] , \dir1_0[1] 
		, \dir1_0[0] }), .out(\hit_dir1[7] ));
	AWDP_INC_422889 i_75574(.O0(fsm5_cnt_0), .fsm5_cnt(fsm5_cnt));
endmodule
module AWDP_partition_5(O0, pfx_sz, twobyte, fpu, sib_dec, displc, mod_dec, imm_sz);
    output [5:0] O0;
    input [4:0] pfx_sz;
    input  twobyte;
    input  fpu;
    input  sib_dec;
    input [2:0] displc;
    input  mod_dec;
    input [2:0] imm_sz;
    // Line 404
    wire [5:0] N18;
    // Line 211
    wire [5:0] O0;
    // Line 406
    wire [6:0] N21;
    // Line 406
    wire [5:0] N28;
    // Line 404
    wire [7:0] N26;

    // Line 404
    assign N18 = pfx_sz + fpu + twobyte;
    // Line 211
    assign O0 = N28;
    // Line 406
    assign N21 = N18 + mod_dec + 7'h1;
    // Line 406
    assign N28 = N26 + imm_sz;
    // Line 404
    assign N26 = N21 + displc + sib_dec;
endmodule

module deco8(in8, indic);

	input [7:0] in8;
	output [72:0] indic;

	wire \indic[10] ;
	wire \indic[14] ;
	wire \indic[15] ;
	wire \indic[22] ;
	wire \indic[0] ;
	wire \indic[1] ;
	wire \indic[2] ;
	wire \indic[3] ;
	wire \indic[4] ;
	wire \indic[5] ;
	wire \indic[6] ;
	wire \indic[7] ;
	wire \indic[8] ;
	wire \indic[9] ;
	wire \indic[11] ;
	wire \indic[12] ;
	wire \indic[13] ;
	wire \indic[16] ;
	wire \indic[17] ;
	wire \indic[18] ;
	wire \indic[19] ;
	wire \indic[20] ;
	wire \indic[21] ;
	wire \indic[23] ;
	wire \indic[24] ;
	wire \indic[25] ;
	wire \indic[26] ;
	wire \indic[27] ;
	wire \indic[28] ;
	wire \indic[29] ;
	wire \indic[30] ;
	wire \indic[32] ;
	wire \indic[33] ;
	wire \indic[34] ;
	wire \indic[35] ;
	wire \indic[36] ;
	wire \indic[37] ;
	wire \indic[38] ;
	wire \indic[39] ;
	wire \indic[40] ;
	wire \indic[41] ;
	wire \indic[42] ;
	wire \indic[43] ;
	wire \indic[44] ;
	wire \indic[45] ;
	wire \indic[46] ;
	wire \indic[47] ;
	wire \indic[48] ;
	wire \indic[49] ;
	wire \indic[50] ;
	wire \indic[51] ;
	wire \indic[53] ;
	wire \indic[54] ;
	wire \indic[55] ;
	wire \indic[56] ;
	wire \indic[57] ;
	wire \indic[58] ;
	wire \indic[59] ;
	wire \indic[60] ;
	wire \indic[61] ;
	wire \indic[62] ;
	wire \indic[63] ;
	wire \indic[64] ;
	wire \indic[67] ;
	wire \indic[68] ;
	wire \indic[69] ;
	wire \indic[70] ;
	wire \indic[71] ;
	wire \indic[72] ;


	assign indic[10] = \indic[10] ;
	assign indic[14] = \indic[14] ;
	assign indic[15] = \indic[15] ;
	assign indic[22] = \indic[22] ;
	assign indic[0] = \indic[0] ;
	assign indic[1] = \indic[1] ;
	assign indic[2] = \indic[2] ;
	assign indic[3] = \indic[3] ;
	assign indic[4] = \indic[4] ;
	assign indic[5] = \indic[5] ;
	assign indic[6] = \indic[6] ;
	assign indic[7] = \indic[7] ;
	assign indic[8] = \indic[8] ;
	assign indic[9] = \indic[9] ;
	assign indic[11] = \indic[11] ;
	assign indic[12] = \indic[12] ;
	assign indic[13] = \indic[13] ;
	assign indic[16] = \indic[16] ;
	assign indic[17] = \indic[17] ;
	assign indic[18] = \indic[18] ;
	assign indic[19] = \indic[19] ;
	assign indic[20] = \indic[20] ;
	assign indic[21] = \indic[21] ;
	assign indic[23] = \indic[23] ;
	assign indic[24] = \indic[24] ;
	assign indic[25] = \indic[25] ;
	assign indic[26] = \indic[26] ;
	assign indic[27] = \indic[27] ;
	assign indic[28] = \indic[28] ;
	assign indic[29] = \indic[29] ;
	assign indic[30] = \indic[30] ;
	assign indic[32] = \indic[32] ;
	assign indic[33] = \indic[33] ;
	assign indic[34] = \indic[34] ;
	assign indic[66] = \indic[35] ;
	assign indic[35] = \indic[35] ;
	assign indic[36] = \indic[36] ;
	assign indic[37] = \indic[37] ;
	assign indic[38] = \indic[38] ;
	assign indic[39] = \indic[39] ;
	assign indic[40] = \indic[40] ;
	assign indic[52] = \indic[41] ;
	assign indic[41] = \indic[41] ;
	assign indic[42] = \indic[42] ;
	assign indic[43] = \indic[43] ;
	assign indic[44] = \indic[44] ;
	assign indic[45] = \indic[45] ;
	assign indic[46] = \indic[46] ;
	assign indic[47] = \indic[47] ;
	assign indic[48] = \indic[48] ;
	assign indic[49] = \indic[49] ;
	assign indic[65] = \indic[50] ;
	assign indic[50] = \indic[50] ;
	assign indic[51] = \indic[51] ;
	assign indic[53] = \indic[53] ;
	assign indic[54] = \indic[54] ;
	assign indic[55] = \indic[55] ;
	assign indic[56] = \indic[56] ;
	assign indic[57] = \indic[57] ;
	assign indic[58] = \indic[58] ;
	assign indic[59] = \indic[59] ;
	assign indic[60] = \indic[60] ;
	assign indic[61] = \indic[61] ;
	assign indic[62] = \indic[62] ;
	assign indic[63] = \indic[63] ;
	assign indic[64] = \indic[64] ;
	assign indic[67] = \indic[67] ;
	assign indic[68] = \indic[68] ;
	assign indic[69] = \indic[69] ;
	assign indic[70] = \indic[70] ;
	assign indic[71] = \indic[71] ;
	assign indic[72] = \indic[72] ;

	notech_and3 i_79(.A(in8[6]), .B(in8[7]), .C(n_75), .Z(n_102));
	notech_and3 i_77(.A(n_33992), .B(n_33993), .C(in8[3]), .Z(n_96));
	notech_and2 i_80(.A(n_33992), .B(n_33991), .Z(n_93));
	notech_and2 i_97(.A(n_33993), .B(n_33991), .Z(n_92));
	notech_and2 i_96(.A(in8[0]), .B(in8[2]), .Z(n_90));
	notech_and4 i_72(.A(in8[6]), .B(in8[7]), .C(in8[4]), .D(n_33995), .Z(n_88
		));
	notech_and3 i_69(.A(in8[6]), .B(in8[7]), .C(n_85), .Z(n_86));
	notech_nor2 i_78(.A(in8[4]), .B(in8[5]), .Z(n_85));
	notech_and2 i_86(.A(n_33991), .B(in8[2]), .Z(n_80));
	notech_and2 i_88(.A(n_78), .B(in8[1]), .Z(n_79));
	notech_nor2 i_71(.A(in8[7]), .B(in8[6]), .Z(n_78));
	notech_nor2 i_70(.A(in8[4]), .B(n_33995), .Z(n_75));
	notech_and3 i_15(.A(in8[0]), .B(in8[3]), .C(in8[2]), .Z(n_73));
	notech_and3 i_10(.A(n_33994), .B(in8[1]), .C(n_33993), .Z(n_72));
	notech_and2 i_23(.A(in8[6]), .B(in8[7]), .Z(n_71));
	notech_and2 i_14(.A(n_33994), .B(n_33993), .Z(n_70));
	notech_and4 i_116(.A(n_92), .B(in8[1]), .C(n_33995), .D(in8[3]), .Z(n_113
		));
	notech_nand3 i_119(.A(\indic[4] ), .B(n_33994), .C(in8[0]), .Z(n_116));
	notech_and4 i_075889(.A(n_71), .B(\indic[41] ), .C(n_33994), .D(n_33993)
		, .Z(\indic[0] ));
	notech_and4 i_1(.A(n_75), .B(\indic[24] ), .C(n_33994), .D(in8[2]), .Z(\indic[1] 
		));
	notech_and4 i_2(.A(n_80), .B(in8[3]), .C(in8[5]), .D(n_79), .Z(\indic[2] 
		));
	notech_and4 i_3(.A(\indic[6] ), .B(n_80), .C(n_78), .D(in8[5]), .Z(\indic[3] 
		));
	notech_and2 i_4(.A(n_78), .B(n_33993), .Z(\indic[4] ));
	notech_and3 i_5(.A(n_75), .B(\indic[24] ), .C(n_33993), .Z(\indic[5] )
		);
	notech_and2 i_6(.A(n_33994), .B(in8[1]), .Z(\indic[6] ));
	notech_and2 i_7(.A(in8[0]), .B(in8[3]), .Z(\indic[7] ));
	notech_ao3 i_8(.A(in8[7]), .B(n_85), .C(in8[6]), .Z(\indic[8] ));
	notech_and4 i_9(.A(in8[6]), .B(in8[7]), .C(n_85), .D(n_33994), .Z(\indic[9] 
		));
	notech_and4 i_11(.A(in8[4]), .B(n_71), .C(n_70), .D(n_33995), .Z(\indic[11] 
		));
	notech_and4 i_12(.A(n_71), .B(\indic[41] ), .C(in8[2]), .D(in8[1]), .Z(\indic[12] 
		));
	notech_ao3 i_13(.A(n_78), .B(n_33995), .C(in8[4]), .Z(\indic[13] ));
	notech_and3 i_16(.A(in8[4]), .B(n_78), .C(in8[5]), .Z(\indic[16] ));
	notech_and4 i_17(.A(n_90), .B(\indic[28] ), .C(n_33994), .D(in8[1]), .Z(\indic[17] 
		));
	notech_ao3 i_18(.A(in8[7]), .B(n_75), .C(in8[6]), .Z(\indic[18] ));
	notech_and2 i_19(.A(n_33992), .B(n_33993), .Z(\indic[19] ));
	notech_and3 i_20(.A(n_33993), .B(n_33991), .C(in8[1]), .Z(\indic[60] )
		);
	notech_and4 i_21(.A(in8[6]), .B(in8[7]), .C(n_85), .D(in8[3]), .Z(\indic[20] 
		));
	notech_and3 i_22(.A(n_33992), .B(n_33991), .C(in8[2]), .Z(\indic[21] )
		);
	notech_and3 i_24(.A(n_78), .B(in8[0]), .C(in8[2]), .Z(\indic[23] ));
	notech_and2 i_25(.A(in8[6]), .B(n_33996), .Z(\indic[24] ));
	notech_nor2 i_26(.A(in8[6]), .B(n_33996), .Z(\indic[25] ));
	notech_and4 i_27(.A(n_78), .B(n_33992), .C(n_33991), .D(in8[2]), .Z(\indic[26] 
		));
	notech_and3 i_28(.A(in8[3]), .B(\indic[5] ), .C(in8[1]), .Z(\indic[27] )
		);
	notech_and3 i_29(.A(in8[4]), .B(\indic[24] ), .C(in8[5]), .Z(\indic[28] 
		));
	notech_ao3 i_30(.A(\indic[43] ), .B(n_33992), .C(in8[0]), .Z(\indic[29] 
		));
	notech_and4 i_31(.A(n_85), .B(in8[0]), .C(\indic[25] ), .D(n_72), .Z(\indic[30] 
		));
	notech_ao3 i_32(.A(\indic[18] ), .B(n_96), .C(in8[0]), .Z(\indic[32] )
		);
	notech_and4 i_33(.A(in8[4]), .B(\indic[25] ), .C(in8[5]), .D(n_33994), .Z
		(\indic[33] ));
	notech_and4 i_34(.A(n_71), .B(n_85), .C(n_70), .D(n_33992), .Z(\indic[34] 
		));
	notech_and3 i_35(.A(n_73), .B(n_86), .C(n_33992), .Z(\indic[36] ));
	notech_and4 i_36(.A(in8[2]), .B(n_33992), .C(n_88), .D(n_33994), .Z(\indic[37] 
		));
	notech_ao3 i_37(.A(n_71), .B(n_75), .C(in8[3]), .Z(\indic[38] ));
	notech_and4 i_38(.A(n_102), .B(in8[1]), .C(\indic[7] ), .D(n_33993), .Z(\indic[39] 
		));
	notech_and4 i_39(.A(\indic[6] ), .B(n_71), .C(\indic[41] ), .D(n_80), .Z
		(\indic[40] ));
	notech_and4 i_40(.A(n_86), .B(n_33993), .C(n_33991), .D(in8[1]), .Z(\indic[42] 
		));
	notech_and4 i_41(.A(\indic[25] ), .B(n_85), .C(n_33994), .D(n_33993), .Z
		(\indic[43] ));
	notech_and4 i_42(.A(n_78), .B(in8[0]), .C(in8[2]), .D(n_33992), .Z(\indic[44] 
		));
	notech_and4 i_43(.A(in8[4]), .B(\indic[25] ), .C(in8[5]), .D(in8[3]), .Z
		(\indic[45] ));
	notech_and4 i_44(.A(in8[6]), .B(in8[7]), .C(n_75), .D(n_96), .Z(\indic[46] 
		));
	notech_and3 i_45(.A(n_75), .B(\indic[24] ), .C(n_96), .Z(\indic[47] ));
	notech_and4 i_46(.A(\indic[25] ), .B(n_75), .C(n_33994), .D(n_33993), .Z
		(\indic[48] ));
	notech_and3 i_47(.A(\indic[25] ), .B(n_96), .C(in8[5]), .Z(\indic[49] )
		);
	notech_and4 i_48(.A(\indic[6] ), .B(n_71), .C(\indic[41] ), .D(n_90), .Z
		(\indic[51] ));
	notech_and2 i_49(.A(in8[4]), .B(in8[5]), .Z(\indic[41] ));
	notech_and3 i_50(.A(\indic[45] ), .B(in8[1]), .C(n_92), .Z(\indic[53] )
		);
	notech_and4 i_51(.A(n_85), .B(n_78), .C(in8[1]), .D(n_73), .Z(\indic[54] 
		));
	notech_and4 i_52(.A(n_93), .B(\indic[41] ), .C(\indic[24] ), .D(n_70), .Z
		(\indic[55] ));
	notech_ao3 i_53(.A(\indic[18] ), .B(\indic[21] ), .C(in8[3]), .Z(\indic[56] 
		));
	notech_ao3 i_54(.A(n_72), .B(n_86), .C(in8[0]), .Z(\indic[57] ));
	notech_and3 i_55(.A(in8[2]), .B(\indic[9] ), .C(n_93), .Z(\indic[58] )
		);
	notech_and4 i_56(.A(in8[0]), .B(in8[2]), .C(\indic[9] ), .D(n_33992), .Z
		(\indic[59] ));
	notech_and4 i_57(.A(in8[4]), .B(n_71), .C(in8[3]), .D(n_33995), .Z(\indic[61] 
		));
	notech_and4 i_58(.A(n_75), .B(\indic[24] ), .C(\indic[6] ), .D(n_80), .Z
		(\indic[62] ));
	notech_and4 i_59(.A(\indic[6] ), .B(n_71), .C(\indic[41] ), .D(n_33993),
		 .Z(\indic[63] ));
	notech_and4 i_60(.A(n_92), .B(in8[3]), .C(n_102), .D(in8[1]), .Z(\indic[64] 
		));
	notech_and4 i_61(.A(\indic[6] ), .B(n_86), .C(in8[0]), .D(in8[2]), .Z(\indic[50] 
		));
	notech_and4 i_62(.A(n_86), .B(n_33991), .C(in8[2]), .D(\indic[6] ), .Z(\indic[35] 
		));
	notech_and4 i_63(.A(\indic[6] ), .B(n_90), .C(n_75), .D(\indic[24] ), .Z
		(\indic[67] ));
	notech_and3 i_64(.A(in8[4]), .B(\indic[25] ), .C(n_113), .Z(\indic[68] )
		);
	notech_ao3 i_65(.A(n_85), .B(n_33992), .C(n_116), .Z(\indic[69] ));
	notech_and4 i_66(.A(\indic[18] ), .B(n_33992), .C(n_33991), .D(in8[2]), 
		.Z(\indic[70] ));
	notech_and4 i_67(.A(n_72), .B(\indic[25] ), .C(n_85), .D(n_33991), .Z(\indic[71] 
		));
	notech_and4 i_68(.A(n_72), .B(\indic[41] ), .C(\indic[25] ), .D(n_33991)
		, .Z(\indic[72] ));
	notech_inv i_34033(.A(in8[0]), .Z(n_33991));
	notech_inv i_34034(.A(in8[1]), .Z(n_33992));
	notech_inv i_34035(.A(in8[2]), .Z(n_33993));
	notech_inv i_34036(.A(in8[3]), .Z(n_33994));
	notech_inv i_34037(.A(in8[5]), .Z(n_33995));
	notech_inv i_34038(.A(in8[7]), .Z(n_33996));
	notech_inv i_34039(.A(n_70), .Z(\indic[14] ));
	notech_inv i_34040(.A(n_71), .Z(\indic[22] ));
	notech_inv i_34041(.A(n_72), .Z(\indic[10] ));
	notech_inv i_34042(.A(n_73), .Z(\indic[15] ));
endmodule
module deco_rm(in8, indic);

	input [7:0] in8;
	output [7:0] indic;




	notech_nand2 i_1(.A(in8[7]), .B(in8[6]), .Z(indic[1]));
	notech_and3 i_077940(.A(in8[2]), .B(n_34229), .C(n_34228), .Z(indic[0])
		);
	notech_and4 i_2(.A(in8[2]), .B(in8[0]), .C(indic[7]), .D(n_34228), .Z(indic
		[2]));
	notech_and2 i_3(.A(in8[7]), .B(n_34227), .Z(indic[3]));
	notech_nor2 i_4(.A(in8[7]), .B(n_34227), .Z(indic[4]));
	notech_nor2 i_5(.A(in8[5]), .B(in8[4]), .Z(indic[5]));
	notech_and4 i_6(.A(indic[7]), .B(in8[2]), .C(in8[1]), .D(n_34229), .Z(indic
		[6]));
	notech_nor2 i_7(.A(in8[7]), .B(in8[6]), .Z(indic[7]));
	notech_inv i_36012(.A(in8[6]), .Z(n_34227));
	notech_inv i_36013(.A(in8[1]), .Z(n_34228));
	notech_inv i_36014(.A(in8[0]), .Z(n_34229));
endmodule
module udecox(op, modrm, twobyte, cpl, adz, opz, jsz, udeco, fpu, emul, ipg_fault
		);

	input [7:0] op;
	input [7:0] modrm;
	input twobyte;
	input [1:0] cpl;
	input adz;
	input [2:0] opz;
	input [3:0] jsz;
	output [127:0] udeco;
	input fpu;
	input emul;
	input ipg_fault;

	wire n_4024;
	wire \udeco[0] ;
	wire \udeco[1] ;
	wire \udeco[2] ;
	wire \udeco[3] ;
	wire \udeco[4] ;
	wire \udeco[5] ;
	wire \udeco[6] ;
	wire \udeco[8] ;
	wire \udeco[9] ;
	wire \udeco[10] ;
	wire \udeco[11] ;
	wire \udeco[12] ;
	wire \udeco[13] ;
	wire \udeco[14] ;
	wire \udeco[15] ;
	wire \udeco[16] ;
	wire \udeco[17] ;
	wire \udeco[18] ;
	wire \udeco[19] ;
	wire \udeco[20] ;
	wire \udeco[21] ;
	wire \udeco[22] ;
	wire \udeco[23] ;
	wire \udeco[24] ;
	wire \udeco[25] ;
	wire \udeco[26] ;
	wire \udeco[27] ;
	wire \udeco[28] ;
	wire \udeco[29] ;
	wire \udeco[30] ;
	wire \udeco[31] ;
	wire \udeco[32] ;
	wire \udeco[33] ;
	wire \udeco[34] ;
	wire \udeco[35] ;
	wire \udeco[36] ;
	wire \udeco[37] ;
	wire \udeco[38] ;
	wire \udeco[39] ;
	wire \udeco[40] ;
	wire \udeco[41] ;
	wire \udeco[42] ;
	wire \udeco[43] ;
	wire \udeco[44] ;
	wire \udeco[45] ;
	wire \udeco[46] ;
	wire \udeco[47] ;
	wire \udeco[48] ;
	wire \udeco[49] ;
	wire \udeco[50] ;
	wire \udeco[51] ;
	wire \udeco[52] ;
	wire \udeco[53] ;
	wire \udeco[54] ;
	wire \udeco[55] ;
	wire \udeco[56] ;
	wire \udeco[57] ;
	wire \udeco[58] ;
	wire \udeco[59] ;
	wire \udeco[60] ;
	wire \udeco[61] ;
	wire \udeco[62] ;
	wire \udeco[63] ;
	wire \udeco[64] ;
	wire \udeco[65] ;
	wire \udeco[66] ;
	wire \udeco[67] ;
	wire \udeco[68] ;
	wire \udeco[69] ;
	wire \udeco[70] ;
	wire \udeco[71] ;
	wire \udeco[72] ;
	wire \udeco[73] ;
	wire \udeco[74] ;
	wire \udeco[75] ;
	wire \udeco[77] ;
	wire \udeco[78] ;
	wire \udeco[80] ;
	wire \udeco[81] ;
	wire \udeco[82] ;
	wire \udeco[83] ;
	wire \udeco[84] ;
	wire \udeco[85] ;
	wire \udeco[86] ;
	wire \udeco[87] ;
	wire \udeco[88] ;
	wire \udeco[89] ;
	wire \udeco[90] ;
	wire \udeco[91] ;
	wire \udeco[92] ;
	wire \udeco[93] ;
	wire \udeco[95] ;
	wire \udeco[96] ;
	wire \udeco[98] ;
	wire \udeco[99] ;
	wire \udeco[100] ;
	wire \udeco[101] ;
	wire \udeco[102] ;
	wire \udeco[103] ;
	wire \udeco[104] ;
	wire \udeco[105] ;
	wire \udeco[106] ;
	wire \udeco[107] ;
	wire \udeco[108] ;
	wire \udeco[109] ;
	wire \udeco[110] ;
	wire \udeco[112] ;
	wire \udeco[113] ;
	wire \udeco[114] ;
	wire \udeco[115] ;
	wire \udeco[116] ;
	wire \udeco[117] ;
	wire \udeco[118] ;
	wire \udeco[119] ;
	wire \udeco[120] ;
	wire \udeco[121] ;
	wire \udeco[122] ;
	wire \udeco[123] ;
	wire \udeco[124] ;
	wire \udeco[125] ;
	wire \udeco[126] ;
	wire \udeco[127] ;


	assign udeco[111] = n_4024;
	assign udeco[0] = \udeco[0] ;
	assign udeco[1] = \udeco[1] ;
	assign udeco[2] = \udeco[2] ;
	assign udeco[3] = \udeco[3] ;
	assign udeco[4] = \udeco[4] ;
	assign udeco[5] = \udeco[5] ;
	assign udeco[7] = \udeco[6] ;
	assign udeco[6] = \udeco[6] ;
	assign udeco[8] = \udeco[8] ;
	assign udeco[9] = \udeco[9] ;
	assign udeco[10] = \udeco[10] ;
	assign udeco[11] = \udeco[11] ;
	assign udeco[12] = \udeco[12] ;
	assign udeco[13] = \udeco[13] ;
	assign udeco[14] = \udeco[14] ;
	assign udeco[15] = \udeco[15] ;
	assign udeco[16] = \udeco[16] ;
	assign udeco[17] = \udeco[17] ;
	assign udeco[18] = \udeco[18] ;
	assign udeco[19] = \udeco[19] ;
	assign udeco[20] = \udeco[20] ;
	assign udeco[21] = \udeco[21] ;
	assign udeco[22] = \udeco[22] ;
	assign udeco[23] = \udeco[23] ;
	assign udeco[24] = \udeco[24] ;
	assign udeco[25] = \udeco[25] ;
	assign udeco[26] = \udeco[26] ;
	assign udeco[27] = \udeco[27] ;
	assign udeco[28] = \udeco[28] ;
	assign udeco[29] = \udeco[29] ;
	assign udeco[30] = \udeco[30] ;
	assign udeco[31] = \udeco[31] ;
	assign udeco[32] = \udeco[32] ;
	assign udeco[33] = \udeco[33] ;
	assign udeco[34] = \udeco[34] ;
	assign udeco[35] = \udeco[35] ;
	assign udeco[36] = \udeco[36] ;
	assign udeco[37] = \udeco[37] ;
	assign udeco[38] = \udeco[38] ;
	assign udeco[39] = \udeco[39] ;
	assign udeco[40] = \udeco[40] ;
	assign udeco[41] = \udeco[41] ;
	assign udeco[42] = \udeco[42] ;
	assign udeco[43] = \udeco[43] ;
	assign udeco[44] = \udeco[44] ;
	assign udeco[45] = \udeco[45] ;
	assign udeco[46] = \udeco[46] ;
	assign udeco[47] = \udeco[47] ;
	assign udeco[48] = \udeco[48] ;
	assign udeco[49] = \udeco[49] ;
	assign udeco[50] = \udeco[50] ;
	assign udeco[51] = \udeco[51] ;
	assign udeco[52] = \udeco[52] ;
	assign udeco[53] = \udeco[53] ;
	assign udeco[54] = \udeco[54] ;
	assign udeco[55] = \udeco[55] ;
	assign udeco[56] = \udeco[56] ;
	assign udeco[57] = \udeco[57] ;
	assign udeco[58] = \udeco[58] ;
	assign udeco[59] = \udeco[59] ;
	assign udeco[60] = \udeco[60] ;
	assign udeco[61] = \udeco[61] ;
	assign udeco[62] = \udeco[62] ;
	assign udeco[63] = \udeco[63] ;
	assign udeco[64] = \udeco[64] ;
	assign udeco[65] = \udeco[65] ;
	assign udeco[66] = \udeco[66] ;
	assign udeco[67] = \udeco[67] ;
	assign udeco[68] = \udeco[68] ;
	assign udeco[69] = \udeco[69] ;
	assign udeco[70] = \udeco[70] ;
	assign udeco[71] = \udeco[71] ;
	assign udeco[72] = \udeco[72] ;
	assign udeco[73] = \udeco[73] ;
	assign udeco[76] = \udeco[74] ;
	assign udeco[74] = \udeco[74] ;
	assign udeco[75] = \udeco[75] ;
	assign udeco[77] = \udeco[77] ;
	assign udeco[79] = \udeco[78] ;
	assign udeco[78] = \udeco[78] ;
	assign udeco[80] = \udeco[80] ;
	assign udeco[81] = \udeco[81] ;
	assign udeco[82] = \udeco[82] ;
	assign udeco[83] = \udeco[83] ;
	assign udeco[84] = \udeco[84] ;
	assign udeco[85] = \udeco[85] ;
	assign udeco[86] = \udeco[86] ;
	assign udeco[87] = \udeco[87] ;
	assign udeco[88] = \udeco[88] ;
	assign udeco[89] = \udeco[89] ;
	assign udeco[90] = \udeco[90] ;
	assign udeco[91] = \udeco[91] ;
	assign udeco[92] = \udeco[92] ;
	assign udeco[94] = \udeco[93] ;
	assign udeco[93] = \udeco[93] ;
	assign udeco[95] = \udeco[95] ;
	assign udeco[96] = \udeco[96] ;
	assign udeco[98] = \udeco[98] ;
	assign udeco[99] = \udeco[99] ;
	assign udeco[97] = \udeco[100] ;
	assign udeco[100] = \udeco[100] ;
	assign udeco[101] = \udeco[101] ;
	assign udeco[102] = \udeco[102] ;
	assign udeco[103] = \udeco[103] ;
	assign udeco[104] = \udeco[104] ;
	assign udeco[105] = \udeco[105] ;
	assign udeco[106] = \udeco[106] ;
	assign udeco[107] = \udeco[107] ;
	assign udeco[108] = \udeco[108] ;
	assign udeco[109] = \udeco[109] ;
	assign udeco[110] = \udeco[110] ;
	assign udeco[112] = \udeco[112] ;
	assign udeco[113] = \udeco[113] ;
	assign udeco[114] = \udeco[114] ;
	assign udeco[115] = \udeco[115] ;
	assign udeco[116] = \udeco[116] ;
	assign udeco[117] = \udeco[117] ;
	assign udeco[118] = \udeco[118] ;
	assign udeco[119] = \udeco[119] ;
	assign udeco[120] = \udeco[120] ;
	assign udeco[121] = \udeco[121] ;
	assign udeco[122] = \udeco[122] ;
	assign udeco[123] = \udeco[123] ;
	assign udeco[124] = \udeco[124] ;
	assign udeco[125] = \udeco[125] ;
	assign udeco[126] = \udeco[126] ;
	assign udeco[127] = \udeco[127] ;

	notech_inv i_11647(.A(n_59638), .Z(n_59647));
	notech_inv i_11643(.A(n_59638), .Z(n_59643));
	notech_inv i_11639(.A(n_59638), .Z(n_59639));
	notech_inv i_11638(.A(op[6]), .Z(n_59638));
	notech_inv i_11635(.A(n_59629), .Z(n_59634));
	notech_inv i_11631(.A(n_59629), .Z(n_59630));
	notech_inv i_11630(.A(op[5]), .Z(n_59629));
	notech_inv i_11623(.A(n_59620), .Z(n_59621));
	notech_inv i_11622(.A(n_34196), .Z(n_59620));
	notech_inv i_11619(.A(n_59611), .Z(n_59616));
	notech_inv i_11615(.A(n_59611), .Z(n_59612));
	notech_inv i_11614(.A(op[4]), .Z(n_59611));
	notech_inv i_11607(.A(n_59602), .Z(n_59603));
	notech_inv i_11606(.A(n_34195), .Z(n_59602));
	notech_inv i_11603(.A(n_59593), .Z(n_59598));
	notech_inv i_11599(.A(n_59593), .Z(n_59594));
	notech_inv i_11598(.A(op[1]), .Z(n_59593));
	notech_inv i_11591(.A(n_59584), .Z(n_59585));
	notech_inv i_11590(.A(n_34192), .Z(n_59584));
	notech_inv i_11587(.A(n_59575), .Z(n_59580));
	notech_inv i_11583(.A(n_59575), .Z(n_59576));
	notech_inv i_11582(.A(op[2]), .Z(n_59575));
	notech_inv i_11573(.A(n_59552), .Z(n_59564));
	notech_inv i_11572(.A(n_59552), .Z(n_59563));
	notech_inv i_11567(.A(n_59552), .Z(n_59558));
	notech_inv i_11562(.A(n_59552), .Z(n_59553));
	notech_inv i_11561(.A(n_2328), .Z(n_59552));
	notech_inv i_11558(.A(n_59543), .Z(n_59548));
	notech_inv i_11554(.A(n_59543), .Z(n_59544));
	notech_inv i_11553(.A(op[0]), .Z(n_59543));
	notech_inv i_11550(.A(n_59532), .Z(n_59539));
	notech_inv i_11549(.A(n_59532), .Z(n_59538));
	notech_inv i_11544(.A(n_59532), .Z(n_59533));
	notech_inv i_11543(.A(op[3]), .Z(n_59532));
	notech_inv i_11540(.A(n_59544), .Z(n_59528));
	notech_inv i_11539(.A(n_59544), .Z(n_59527));
	notech_inv i_11534(.A(n_59544), .Z(n_59522));
	notech_inv i_11529(.A(n_59538), .Z(n_59516));
	notech_inv i_11524(.A(n_59538), .Z(n_59511));
	notech_inv i_11516(.A(n_59501), .Z(n_59502));
	notech_inv i_11515(.A(n_2360), .Z(n_59501));
	notech_inv i_11508(.A(n_59492), .Z(n_59493));
	notech_inv i_11507(.A(n_2286), .Z(n_59492));
	notech_inv i_11496(.A(n_59478), .Z(n_59479));
	notech_inv i_11495(.A(modrm[5]), .Z(n_59478));
	notech_inv i_11488(.A(n_59469), .Z(n_59470));
	notech_inv i_11487(.A(n_34193), .Z(n_59469));
	notech_inv i_11480(.A(n_59460), .Z(n_59461));
	notech_inv i_11479(.A(n_2271), .Z(n_59460));
	notech_inv i_11472(.A(n_59451), .Z(n_59452));
	notech_inv i_11471(.A(n_34010), .Z(n_59451));
	notech_inv i_11464(.A(n_59442), .Z(n_59443));
	notech_inv i_11463(.A(n_34202), .Z(n_59442));
	notech_inv i_11456(.A(n_59433), .Z(n_59434));
	notech_inv i_11455(.A(n_2325), .Z(n_59433));
	notech_inv i_11448(.A(n_59424), .Z(n_59425));
	notech_inv i_11447(.A(n_2282), .Z(n_59424));
	notech_inv i_11440(.A(n_59415), .Z(n_59416));
	notech_inv i_11439(.A(n_2410), .Z(n_59415));
	notech_and4 i_1531(.A(n_2839), .B(n_1543), .C(n_2931), .D(n_2924), .Z(n_2934
		));
	notech_ao3 i_1534(.A(n_2934), .B(n_2904), .C(n_34110), .Z(n_2936));
	notech_and2 i_793(.A(n_2179), .B(n_1603), .Z(n_2937));
	notech_and4 i_1535(.A(n_2663), .B(n_2352), .C(n_2937), .D(n_2567), .Z(n_2939
		));
	notech_and4 i_1546(.A(n_3993), .B(n_4040), .C(n_3733), .D(n_1907), .Z(n_2942
		));
	notech_and4 i_306(.A(n_2137), .B(n_2942), .C(n_2026), .D(n_3984), .Z(n_2945
		));
	notech_and3 i_770(.A(n_2638), .B(n_2014), .C(n_1896), .Z(n_2946));
	notech_and4 i_1552(.A(n_4019), .B(n_2080), .C(n_2945), .D(n_2946), .Z(n_2949
		));
	notech_and4 i_1557(.A(n_2189), .B(n_2206), .C(n_2028), .D(n_2457), .Z(n_2953
		));
	notech_and4 i_245(.A(n_2611), .B(n_2949), .C(n_2953), .D(n_2484), .Z(n_2955
		));
	notech_and4 i_1561(.A(n_2435), .B(n_2631), .C(n_1953), .D(n_2030), .Z(n_2958
		));
	notech_and4 i_303(.A(n_2141), .B(n_4013), .C(n_2058), .D(n_2958), .Z(n_2959
		));
	notech_and3 i_1569(.A(n_2033), .B(n_2032), .C(n_4020), .Z(n_2961));
	notech_and4 i_1572(.A(n_2176), .B(n_1837), .C(n_2034), .D(n_2961), .Z(n_2964
		));
	notech_and4 i_724(.A(n_2332), .B(n_2964), .C(n_2091), .D(n_3972), .Z(n_2967
		));
	notech_and4 i_521(.A(n_34077), .B(n_34042), .C(n_34076), .D(n_2031), .Z(n_2969
		));
	notech_ao4 i_1576(.A(n_3963), .B(n_2574), .C(n_2362), .D(n_2331), .Z(n_2970
		));
	notech_and4 i_1578(.A(n_3992), .B(n_1895), .C(n_2970), .D(n_3672), .Z(n_2972
		));
	notech_and4 i_1581(.A(n_2972), .B(n_2406), .C(n_2969), .D(n_2967), .Z(n_2975
		));
	notech_ao3 i_653(.A(n_2668), .B(n_3777), .C(n_34014), .Z(n_2978));
	notech_and4 i_1607(.A(n_843), .B(n_1332), .C(n_2494), .D(n_2046), .Z(n_2983
		));
	notech_and3 i_1611(.A(n_3994), .B(n_2983), .C(n_1340), .Z(n_2985));
	notech_and4 i_1615(.A(n_1329), .B(n_2021), .C(n_2562), .D(n_2985), .Z(n_2987
		));
	notech_ao4 i_510(.A(n_2098), .B(n_2101), .C(n_4065), .D(n_2027), .Z(n_2988
		));
	notech_ao4 i_1598(.A(n_34080), .B(n_34127), .C(adz), .D(n_2305), .Z(n_2989
		));
	notech_and4 i_1596(.A(n_2040), .B(n_2219), .C(n_34064), .D(n_2041), .Z(n_2992
		));
	notech_and4 i_1600(.A(n_2042), .B(n_2045), .C(n_2989), .D(n_2992), .Z(n_2995
		));
	notech_and4 i_1603(.A(n_2195), .B(n_4022), .C(n_2995), .D(n_1346), .Z(n_2999
		));
	notech_and4 i_1610(.A(n_2050), .B(n_2999), .C(n_2051), .D(n_2053), .Z(n_3002
		));
	notech_and4 i_1616(.A(n_3002), .B(n_1728), .C(n_2665), .D(n_2246), .Z(n_3005
		));
	notech_ao4 i_1633(.A(n_34080), .B(n_2574), .C(n_34138), .D(n_2355), .Z(n_3008
		));
	notech_ao3 i_1635(.A(n_2829), .B(n_3008), .C(n_3820), .Z(n_3010));
	notech_and4 i_244(.A(n_2392), .B(n_2967), .C(n_3955), .D(n_3010), .Z(n_3013
		));
	notech_and4 i_1640(.A(n_2435), .B(n_2631), .C(n_1526), .D(n_4025), .Z(n_3015
		));
	notech_and4 i_1643(.A(n_3015), .B(n_2379), .C(n_2852), .D(n_1905), .Z(n_3018
		));
	notech_and2 i_726(.A(n_3890), .B(n_2238), .Z(n_3021));
	notech_and4 i_1656(.A(n_1855), .B(n_1854), .C(n_4028), .D(n_2071), .Z(n_3023
		));
	notech_and4 i_1662(.A(n_2073), .B(n_3023), .C(n_1656), .D(n_2076), .Z(n_3026
		));
	notech_ao3 i_1669(.A(n_3026), .B(n_3021), .C(n_2077), .Z(n_3028));
	notech_and3 i_176(.A(n_4026), .B(n_1284), .C(n_4027), .Z(n_3030));
	notech_and4 i_1672(.A(n_3977), .B(n_1306), .C(n_3030), .D(n_3028), .Z(n_3033
		));
	notech_and4 i_1653(.A(n_2252), .B(n_222298895), .C(n_2188), .D(n_2070), 
		.Z(n_3039));
	notech_and4 i_1659(.A(n_2190), .B(n_3039), .C(n_2709), .D(n_2072), .Z(n_3042
		));
	notech_and4 i_1668(.A(n_3042), .B(n_4029), .C(n_2074), .D(n_1290), .Z(n_3045
		));
	notech_and4 i_1671(.A(n_3045), .B(n_2075), .C(n_2598), .D(n_4005), .Z(n_3046
		));
	notech_and4 i_1675(.A(n_4055), .B(n_1857), .C(n_3046), .D(n_3033), .Z(n_3048
		));
	notech_and2 i_549(.A(n_2264), .B(n_1911), .Z(n_3049));
	notech_and4 i_1677(.A(n_3049), .B(n_3048), .C(n_2789), .D(n_34015), .Z(n_3052
		));
	notech_and4 i_1679(.A(n_1329), .B(n_2021), .C(n_2826), .D(n_3052), .Z(n_3054
		));
	notech_and3 i_210(.A(n_4027), .B(n_4036), .C(n_4076), .Z(n_3056));
	notech_and4 i_1720(.A(n_2151), .B(n_3992), .C(n_3977), .D(n_34050), .Z(n_3059
		));
	notech_and2 i_624(.A(n_4017), .B(n_4019), .Z(n_3061));
	notech_and3 i_556(.A(n_2192), .B(n_4017), .C(n_3981), .Z(n_3062));
	notech_and4 i_1527(.A(n_1434), .B(n_2928), .C(n_34044), .D(n_4016), .Z(n_2931
		));
	notech_and3 i_206(.A(n_34063), .B(n_1958), .C(n_2377), .Z(n_3064));
	notech_ao4 i_1780(.A(n_34143), .B(n_59528), .C(n_34185), .D(n_34200), .Z
		(n_3067));
	notech_and3 i_1782(.A(n_3067), .B(n_2086), .C(n_3980), .Z(n_3069));
	notech_and4 i_1787(.A(n_4047), .B(n_223496909), .C(n_3069), .D(n_2305), 
		.Z(n_3072));
	notech_ao4 i_1788(.A(n_2124), .B(n_59516), .C(n_2333), .D(n_2359), .Z(n_3073
		));
	notech_and4 i_1792(.A(n_4017), .B(n_3073), .C(n_3072), .D(n_4019), .Z(n_3075
		));
	notech_and4 i_1799(.A(n_3075), .B(n_3967), .C(n_2090), .D(n_3064), .Z(n_3078
		));
	notech_and2 i_4702(.A(n_34046), .B(n_4082), .Z(n_3079));
	notech_and4 i_1789(.A(n_3079), .B(n_2087), .C(n_2089), .D(n_1624), .Z(n_3083
		));
	notech_and4 i_1795(.A(n_3083), .B(n_2579), .C(n_2609), .D(n_3981), .Z(n_3086
		));
	notech_and4 i_1800(.A(n_2663), .B(n_3086), .C(n_2978), .D(n_2091), .Z(n_3089
		));
	notech_and4 i_1803(.A(n_3089), .B(n_3078), .C(n_5254), .D(n_34071), .Z(n_3091
		));
	notech_and2 i_1808(.A(n_4040), .B(n_733), .Z(n_3095));
	notech_and4 i_258(.A(n_4002), .B(n_1332), .C(n_1329), .D(n_3095), .Z(n_3098
		));
	notech_ao3 i_809(.A(n_4055), .B(n_2097), .C(n_2100), .Z(n_3102));
	notech_ao4 i_560(.A(n_2499), .B(n_2485), .C(n_2596), .D(n_2302), .Z(n_3103
		));
	notech_and4 i_1821(.A(n_1984), .B(n_1801), .C(n_2159), .D(n_2104), .Z(n_3105
		));
	notech_and3 i_20377856(.A(n_2206), .B(n_4028), .C(n_2790), .Z(n_3107));
	notech_and3 i_296(.A(n_3965), .B(n_2579), .C(n_34074), .Z(n_2928));
	notech_and3 i_64777826(.A(n_2238), .B(n_4053), .C(n_2159), .Z(n_3109));
	notech_and4 i_1864(.A(n_3109), .B(n_222198894), .C(n_3107), .D(n_34079),
		 .Z(n_3111));
	notech_and4 i_1869(.A(n_3111), .B(n_2327), .C(n_2103), .D(n_34046), .Z(n_3114
		));
	notech_and4 i_1874(.A(n_34063), .B(n_4044), .C(n_3114), .D(n_4027), .Z(n_3117
		));
	notech_and4 i_1877(.A(n_2057), .B(n_1794), .C(n_2105), .D(n_3117), .Z(n_3119
		));
	notech_and4 i_1884(.A(n_3119), .B(n_2480), .C(n_2108), .D(n_2572), .Z(n_3122
		));
	notech_and2 i_719(.A(n_2218), .B(n_3970), .Z(n_3124));
	notech_and4 i_1887(.A(n_3970), .B(n_3122), .C(n_2218), .D(n_2116), .Z(n_3126
		));
	notech_ao3 i_317(.A(n_2609), .B(n_1792), .C(n_1795), .Z(n_3128));
	notech_and4 i_1871(.A(n_1932), .B(n_2123), .C(n_4041), .D(n_4043), .Z(n_3131
		));
	notech_and4 i_1879(.A(n_3131), .B(n_2107), .C(n_2104), .D(n_2106), .Z(n_3134
		));
	notech_and4 i_1883(.A(n_2176), .B(n_2195), .C(n_1970), .D(n_3134), .Z(n_3136
		));
	notech_and4 i_1888(.A(n_34148), .B(n_3128), .C(n_3136), .D(n_34044), .Z(n_3138
		));
	notech_and4 i_1891(.A(n_3098), .B(n_3126), .C(n_2109), .D(n_3138), .Z(n_3141
		));
	notech_and2 i_4754(.A(n_2688), .B(n_3739), .Z(n_3143));
	notech_and4 i_1924(.A(n_2579), .B(n_1970), .C(n_222898901), .D(n_2125), 
		.Z(n_3145));
	notech_and4 i_1917(.A(n_3061), .B(n_4032), .C(n_3981), .D(n_2122), .Z(n_3150
		));
	notech_and4 i_1919(.A(n_574), .B(n_4046), .C(n_2121), .D(n_3150), .Z(n_3151
		));
	notech_ao4 i_746(.A(n_2297), .B(n_2118), .C(n_2382), .D(n_2325), .Z(n_3152
		));
	notech_and4 i_444(.A(n_1855), .B(n_1854), .C(n_2111), .D(n_2255), .Z(n_3154
		));
	notech_and3 i_1904(.A(n_2119), .B(n_223496909), .C(n_34185), .Z(n_3157)
		);
	notech_and4 i_1908(.A(n_2627), .B(n_34046), .C(n_2364), .D(n_3157), .Z(n_3160
		));
	notech_and4 i_1910(.A(n_3154), .B(n_3160), .C(n_3992), .D(n_2120), .Z(n_3162
		));
	notech_and4 i_1918(.A(n_3152), .B(n_709), .C(n_3162), .D(n_2465), .Z(n_3165
		));
	notech_and4 i_1923(.A(n_673), .B(n_3165), .C(n_3151), .D(n_960), .Z(n_3168
		));
	notech_and4 i_1927(.A(n_3168), .B(n_703), .C(n_2126), .D(n_3145), .Z(n_3171
		));
	notech_nand2 i_441(.A(n_2625), .B(n_3779), .Z(n_3174));
	notech_and4 i_817(.A(n_2631), .B(n_1780), .C(n_2137), .D(n_34016), .Z(n_3177
		));
	notech_and3 i_811(.A(n_4058), .B(n_2049), .C(n_2129), .Z(n_3178));
	notech_and2 i_234(.A(n_3178), .B(n_2130), .Z(n_3179));
	notech_and3 i_1937(.A(n_2141), .B(n_2131), .C(n_34057), .Z(n_3181));
	notech_and4 i_1940(.A(n_2258), .B(n_3975), .C(n_3181), .D(n_34031), .Z(n_3184
		));
	notech_and3 i_1988(.A(n_3982), .B(n_34043), .C(n_455), .Z(n_3187));
	notech_and4 i_1981(.A(n_3977), .B(n_2377), .C(n_2134), .D(n_2978), .Z(n_3193
		));
	notech_and4 i_1986(.A(n_2218), .B(n_3970), .C(n_3193), .D(n_444), .Z(n_3195
		));
	notech_and3 i_37477842(.A(n_2104), .B(n_3154), .C(n_4046), .Z(n_3197));
	notech_ao4 i_1972(.A(n_2400), .B(n_2497), .C(n_2278), .D(n_2339), .Z(n_3200
		));
	notech_and4 i_1974(.A(n_3197), .B(n_2216), .C(n_4051), .D(n_3200), .Z(n_3201
		));
	notech_and4 i_1976(.A(n_34063), .B(n_4019), .C(n_3201), .D(n_1923), .Z(n_3204
		));
	notech_and4 i_1983(.A(n_3204), .B(n_2579), .C(n_2395), .D(n_3021), .Z(n_3207
		));
	notech_and4 i_1985(.A(n_4002), .B(n_1526), .C(n_3207), .D(n_2166), .Z(n_3208
		));
	notech_and4 i_1991(.A(n_2522), .B(n_3208), .C(n_3195), .D(n_2352), .Z(n_3211
		));
	notech_and4 i_1993(.A(n_3177), .B(n_3187), .C(n_3211), .D(n_2893), .Z(n_3213
		));
	notech_and4 i_2032(.A(n_2555), .B(n_1873), .C(n_3102), .D(n_3178), .Z(n_3217
		));
	notech_and4 i_2039(.A(n_3217), .B(n_2352), .C(n_2308), .D(n_2294), .Z(n_3219
		));
	notech_and4 i_2030(.A(n_3021), .B(n_2513), .C(n_3972), .D(n_2144), .Z(n_3223
		));
	notech_ao3 i_2013(.A(n_4028), .B(n_1829), .C(n_2142), .Z(n_3225));
	notech_and4 i_2007(.A(n_2433), .B(n_4048), .C(n_1263), .D(n_696), .Z(n_3227
		));
	notech_and4 i_2010(.A(n_2140), .B(n_4014), .C(n_2141), .D(n_3227), .Z(n_3230
		));
	notech_and4 i_2015(.A(n_3230), .B(n_4051), .C(n_3225), .D(n_34057), .Z(n_3233
		));
	notech_and4 i_2019(.A(n_1656), .B(n_4007), .C(n_3233), .D(n_34040), .Z(n_3236
		));
	notech_and3 i_2020(.A(n_1958), .B(n_4022), .C(n_34031), .Z(n_3240));
	notech_and4 i_2026(.A(n_3103), .B(n_3240), .C(n_2143), .D(n_34047), .Z(n_3243
		));
	notech_and4 i_2028(.A(n_3236), .B(n_3243), .C(n_3697), .D(n_2614), .Z(n_3244
		));
	notech_and4 i_2037(.A(n_3244), .B(n_466), .C(n_2854), .D(n_3223), .Z(n_3247
		));
	notech_and4 i_259(.A(n_3970), .B(n_2136), .C(n_2137), .D(n_1332), .Z(n_3250
		));
	notech_ao4 i_571(.A(n_2139), .B(n_34142), .C(n_2458), .D(n_2275), .Z(n_3252
		));
	notech_and4 i_2038(.A(n_3252), .B(n_3250), .C(n_2145), .D(n_455), .Z(n_3254
		));
	notech_and4 i_2042(.A(n_3254), .B(n_3247), .C(n_3219), .D(n_2834), .Z(n_3257
		));
	notech_ao4 i_171(.A(n_2278), .B(n_2154), .C(n_2318), .D(n_2161), .Z(n_3261
		));
	notech_and3 i_2073(.A(n_3970), .B(n_2166), .C(n_2168), .Z(n_3263));
	notech_and4 i_2082(.A(n_2065), .B(n_3261), .C(n_3263), .D(n_1623), .Z(n_3266
		));
	notech_and4 i_2091(.A(n_2538), .B(n_2663), .C(n_2173), .D(n_3266), .Z(n_3269
		));
	notech_and4 i_2097(.A(n_3979), .B(n_3269), .C(n_4032), .D(n_3984), .Z(n_3271
		));
	notech_and4 i_2105(.A(n_3271), .B(n_2526), .C(n_3179), .D(n_2175), .Z(n_3273
		));
	notech_and4 i_764(.A(n_2234), .B(n_4005), .C(n_2159), .D(n_4004), .Z(n_3275
		));
	notech_ao4 i_627(.A(n_34136), .B(n_2517), .C(n_3963), .D(n_2407), .Z(n_3276
		));
	notech_or4 i_98(.A(n_2403), .B(n_2311), .C(n_59580), .D(n_34192), .Z(n_3277
		));
	notech_and2 i_360477875(.A(n_1797), .B(n_2106), .Z(n_3279));
	notech_ao4 i_1502(.A(n_2140), .B(n_59548), .C(n_2433), .D(n_59539), .Z(n_2925
		));
	notech_and3 i_38277841(.A(n_1993), .B(n_2665), .C(n_3143), .Z(n_3280));
	notech_ao3 i_2067(.A(n_3280), .B(n_3279), .C(n_34176), .Z(n_3282));
	notech_and3 i_2068(.A(n_1925), .B(n_3107), .C(n_3282), .Z(n_3283));
	notech_and4 i_2072(.A(n_2516), .B(n_3283), .C(n_2163), .D(n_1828), .Z(n_3286
		));
	notech_and4 i_2079(.A(n_3286), .B(n_2170), .C(n_3276), .D(n_2169), .Z(n_3289
		));
	notech_ao4 i_777(.A(n_2495), .B(n_2376), .C(n_2337), .D(n_34053), .Z(n_3290
		));
	notech_and4 i_2083(.A(n_3290), .B(n_2076), .C(n_3289), .D(n_3890), .Z(n_3293
		));
	notech_and4 i_2087(.A(n_3975), .B(n_4037), .C(n_2172), .D(n_2174), .Z(n_3297
		));
	notech_and4 i_2092(.A(n_3293), .B(n_1526), .C(n_2639), .D(n_3297), .Z(n_3299
		));
	notech_and4 i_2103(.A(n_673), .B(n_3299), .C(n_3275), .D(n_3177), .Z(n_3302
		));
	notech_and4 i_2096(.A(n_3987), .B(n_2029), .C(n_3128), .D(n_1712), .Z(n_3307
		));
	notech_and4 i_2104(.A(n_3252), .B(n_3307), .C(n_2563), .D(n_497), .Z(n_3309
		));
	notech_ao4 i_2112(.A(n_2329), .B(n_2448), .C(n_2407), .D(n_2408), .Z(n_3312
		));
	notech_and2 i_2127(.A(n_2188), .B(n_4013), .Z(n_3316));
	notech_and4 i_2130(.A(n_2189), .B(n_2234), .C(n_2190), .D(n_3316), .Z(n_3319
		));
	notech_and4 i_2139(.A(n_2192), .B(n_3319), .C(n_4051), .D(n_3290), .Z(n_3322
		));
	notech_ao4 i_2131(.A(n_2278), .B(n_34151), .C(n_34128), .D(n_2531), .Z(n_3323
		));
	notech_and4 i_2140(.A(n_3323), .B(n_2631), .C(n_3276), .D(n_34037), .Z(n_3326
		));
	notech_and4 i_2150(.A(n_3326), .B(n_3322), .C(n_2196), .D(n_34074), .Z(n_3329
		));
	notech_and4 i_2138(.A(n_2193), .B(n_223496909), .C(n_2327), .D(n_34039),
		 .Z(n_3333));
	notech_and4 i_2147(.A(n_3333), .B(n_1892), .C(n_3672), .D(n_1806), .Z(n_3336
		));
	notech_and4 i_2154(.A(n_3329), .B(n_2380), .C(n_2377), .D(n_3336), .Z(n_3338
		));
	notech_and4 i_2162(.A(n_2198), .B(n_3056), .C(n_1970), .D(n_3338), .Z(n_3340
		));
	notech_and4 i_2172(.A(n_3340), .B(n_3728), .C(n_493), .D(n_2200), .Z(n_3343
		));
	notech_ao4 i_2144(.A(n_2186), .B(n_59516), .C(n_1819), .D(n_2285), .Z(n_3347
		));
	notech_and4 i_2152(.A(n_3347), .B(n_2195), .C(n_2639), .D(n_2565), .Z(n_3349
		));
	notech_and4 i_2160(.A(n_2723), .B(n_3349), .C(n_2533), .D(n_2197), .Z(n_3351
		));
	notech_and4 i_2167(.A(n_2663), .B(n_3351), .C(n_2945), .D(n_2183), .Z(n_3353
		));
	notech_and3 i_453(.A(n_4032), .B(n_2365), .C(n_2181), .Z(n_3355));
	notech_and4 i_2161(.A(n_4034), .B(n_2465), .C(n_4053), .D(n_1924), .Z(n_3358
		));
	notech_and4 i_1529(.A(n_2921), .B(n_2534), .C(n_2620), .D(n_2656), .Z(n_2924
		));
	notech_and3 i_3668(.A(n_4031), .B(n_4056), .C(n_34071), .Z(n_3360));
	notech_and4 i_2168(.A(n_497), .B(n_3358), .C(n_3360), .D(n_2199), .Z(n_3362
		));
	notech_and4 i_2173(.A(n_3362), .B(n_533), .C(n_3353), .D(n_3355), .Z(n_3364
		));
	notech_and3 i_2177(.A(n_2258), .B(n_3739), .C(n_2202), .Z(n_3367));
	notech_and4 i_375(.A(n_3049), .B(n_2790), .C(n_3367), .D(n_1905), .Z(n_3370
		));
	notech_and4 i_2203(.A(n_4005), .B(n_2532), .C(n_2218), .D(n_3779), .Z(n_3373
		));
	notech_ao4 i_488(.A(n_2412), .B(n_34152), .C(n_2455), .D(n_2297), .Z(n_3374
		));
	notech_and4 i_2195(.A(n_2637), .B(n_3374), .C(n_3965), .D(n_2207), .Z(n_3377
		));
	notech_and4 i_2186(.A(n_4048), .B(n_3109), .C(n_2516), .D(n_2206), .Z(n_3381
		));
	notech_and4 i_2189(.A(n_1855), .B(n_3381), .C(n_1854), .D(n_34039), .Z(n_3383
		));
	notech_and4 i_2192(.A(n_2668), .B(n_3383), .C(n_3973), .D(n_34036), .Z(n_3385
		));
	notech_and4 i_2199(.A(n_3385), .B(n_3377), .C(n_2305), .D(n_4056), .Z(n_3388
		));
	notech_ao4 i_815(.A(n_2205), .B(n_2285), .C(n_2331), .D(n_2586), .Z(n_3389
		));
	notech_and4 i_2202(.A(n_3777), .B(n_4055), .C(n_3389), .D(n_3388), .Z(n_3392
		));
	notech_and4 i_2205(.A(n_1796), .B(n_3392), .C(n_3373), .D(n_4029), .Z(n_3394
		));
	notech_and4 i_2208(.A(n_3250), .B(n_3394), .C(n_960), .D(n_3370), .Z(n_3397
		));
	notech_and2 i_408977874(.A(n_4079), .B(n_1984), .Z(n_3402));
	notech_and4 i_59977833(.A(n_2192), .B(n_2305), .C(n_34057), .D(n_34036),
		 .Z(n_3403));
	notech_and4 i_2219(.A(n_3403), .B(n_3402), .C(n_4048), .D(n_2668), .Z(n_3406
		));
	notech_and4 i_2222(.A(n_4058), .B(n_3406), .C(n_3838), .D(n_2216), .Z(n_3408
		));
	notech_and4 i_2225(.A(n_3408), .B(n_4029), .C(n_2217), .D(n_730), .Z(n_3411
		));
	notech_and4 i_2228(.A(n_2218), .B(n_3411), .C(n_3030), .D(n_3981), .Z(n_3413
		));
	notech_and4 i_2232(.A(n_3413), .B(n_2538), .C(n_2111), .D(n_34044), .Z(n_3415
		));
	notech_and4 i_2233(.A(n_2395), .B(n_218), .C(n_4049), .D(n_2411), .Z(n_3419
		));
	notech_and4 i_2236(.A(n_2534), .B(n_3415), .C(n_3250), .D(n_3419), .Z(n_3421
		));
	notech_ao4 i_2214(.A(n_34136), .B(n_2594), .C(n_2391), .D(n_34053), .Z(n_3422
		));
	notech_and4 i_2239(.A(n_204), .B(n_3421), .C(n_3370), .D(n_2379), .Z(n_3425
		));
	notech_and4 i_2281(.A(n_3994), .B(n_204), .C(n_3370), .D(n_4085), .Z(n_3429
		));
	notech_ao4 i_2258(.A(n_2678), .B(n_34196), .C(n_2485), .D(n_2689), .Z(n_3430
		));
	notech_and4 i_2261(.A(n_2631), .B(n_3374), .C(n_3430), .D(n_2222), .Z(n_3433
		));
	notech_and4 i_2253(.A(n_3998), .B(n_2220), .C(n_3402), .D(n_34075), .Z(n_3437
		));
	notech_and4 i_2257(.A(n_2221), .B(n_2130), .C(n_2223), .D(n_3437), .Z(n_3440
		));
	notech_and4 i_2264(.A(n_3975), .B(n_3103), .C(n_3389), .D(n_3440), .Z(n_3443
		));
	notech_and4 i_2268(.A(n_3433), .B(n_3443), .C(n_2116), .D(n_34050), .Z(n_3445
		));
	notech_and4 i_2269(.A(n_3030), .B(n_1130), .C(n_2695), .D(n_2854), .Z(n_3449
		));
	notech_and4 i_2274(.A(n_2675), .B(n_3449), .C(n_3445), .D(n_34045), .Z(n_3451
		));
	notech_and4 i_2272(.A(n_2076), .B(n_2080), .C(n_3275), .D(n_34031), .Z(n_3452
		));
	notech_and4 i_2278(.A(n_444), .B(n_960), .C(n_2722), .D(n_2226), .Z(n_3457
		));
	notech_and4 i_2280(.A(n_2534), .B(n_3452), .C(n_3451), .D(n_3457), .Z(n_3458
		));
	notech_and4 i_2326(.A(n_2294), .B(n_2587), .C(n_1340), .D(n_2228), .Z(n_3463
		));
	notech_and4 i_2330(.A(n_3994), .B(n_3463), .C(n_34045), .D(n_2850), .Z(n_3465
		));
	notech_ao4 i_2300(.A(n_2363), .B(n_2412), .C(n_2065), .D(n_34192), .Z(n_3466
		));
	notech_and4 i_2308(.A(n_3466), .B(n_3154), .C(n_2598), .D(n_4037), .Z(n_3469
		));
	notech_and4 i_2318(.A(n_3469), .B(n_2614), .C(n_1332), .D(n_34029), .Z(n_3472
		));
	notech_and4 i_2312(.A(n_2238), .B(n_4031), .C(n_2239), .D(n_2099), .Z(n_3475
		));
	notech_and4 i_2321(.A(n_4034), .B(n_3475), .C(n_3062), .D(n_3472), .Z(n_3478
		));
	notech_and2 i_631(.A(n_2229), .B(n_3965), .Z(n_3481));
	notech_and4 i_2297(.A(n_2231), .B(n_3279), .C(n_2232), .D(n_2233), .Z(n_3485
		));
	notech_and4 i_2301(.A(n_4028), .B(n_3485), .C(n_223496909), .D(n_4044), 
		.Z(n_3488));
	notech_and4 i_2307(.A(n_3488), .B(n_2394), .C(n_2237), .D(n_4084), .Z(n_3490
		));
	notech_and4 i_2310(.A(n_4007), .B(n_34036), .C(n_1936), .D(n_3490), .Z(n_3491
		));
	notech_and4 i_2317(.A(n_2572), .B(n_34043), .C(n_3481), .D(n_3491), .Z(n_3494
		));
	notech_and4 i_2322(.A(n_4076), .B(n_3494), .C(n_2615), .D(n_3128), .Z(n_3496
		));
	notech_and4 i_2327(.A(n_3496), .B(n_3252), .C(n_2240), .D(n_3478), .Z(n_3498
		));
	notech_and4 i_2331(.A(n_1329), .B(n_2021), .C(n_3498), .D(n_2898), .Z(n_3500
		));
	notech_and2 i_2381(.A(n_2723), .B(n_2946), .Z(n_3507));
	notech_ao4 i_2368(.A(n_59528), .B(n_2250), .C(n_2285), .D(n_2245), .Z(n_3508
		));
	notech_and2 i_21977855(.A(n_4007), .B(n_4047), .Z(n_3510));
	notech_and4 i_2356(.A(n_1193), .B(n_1833), .C(n_3510), .D(n_34032), .Z(n_3513
		));
	notech_and4 i_2359(.A(n_2252), .B(n_3513), .C(n_2253), .D(n_2254), .Z(n_3516
		));
	notech_ao3 i_2361(.A(n_3516), .B(n_2255), .C(n_1807), .Z(n_3518));
	notech_and4 i_2364(.A(n_4058), .B(n_2256), .C(n_2257), .D(n_3518), .Z(n_3521
		));
	notech_and4 i_2367(.A(n_2233), .B(n_1938), .C(n_3521), .D(n_2571), .Z(n_3523
		));
	notech_and4 i_2374(.A(n_2263), .B(n_3523), .C(n_3508), .D(n_2262), .Z(n_3525
		));
	notech_and4 i_2375(.A(n_4017), .B(n_4019), .C(n_4022), .D(n_2264), .Z(n_3528
		));
	notech_and4 i_2379(.A(n_2206), .B(n_733), .C(n_2265), .D(n_3528), .Z(n_3530
		));
	notech_and4 i_2384(.A(n_3525), .B(n_3530), .C(n_3507), .D(n_2266), .Z(n_3532
		));
	notech_ao4 i_2366(.A(n_34136), .B(n_34127), .C(n_2285), .D(n_2288), .Z(n_3534
		));
	notech_and4 i_2377(.A(n_3534), .B(n_3261), .C(n_2532), .D(n_3481), .Z(n_3537
		));
	notech_and4 i_2385(.A(n_4046), .B(n_3537), .C(n_3967), .D(n_34071), .Z(n_3540
		));
	notech_and4 i_2390(.A(n_3540), .B(n_3532), .C(n_466), .D(n_2790), .Z(n_3542
		));
	notech_and4 i_2391(.A(n_2304), .B(n_960), .C(n_3542), .D(n_2267), .Z(n_3543
		));
	notech_and3 i_3610(.A(n_223496909), .B(n_1792), .C(n_3355), .Z(n_3545)
		);
	notech_and4 i_2394(.A(n_68), .B(n_901), .C(n_3543), .D(n_3545), .Z(n_3548
		));
	notech_ao3 i_2425(.A(n_894), .B(n_2620), .C(n_34105), .Z(n_3552));
	notech_and4 i_2431(.A(n_2826), .B(n_3452), .C(n_2157), .D(n_3552), .Z(n_3553
		));
	notech_and4 i_2432(.A(n_2884), .B(n_1728), .C(n_2379), .D(n_2850), .Z(n_3556
		));
	notech_and3 i_2433(.A(n_4016), .B(n_2498), .C(n_3972), .Z(n_3558));
	notech_and4 i_2440(.A(n_3556), .B(n_3553), .C(n_3558), .D(n_2937), .Z(n_3560
		));
	notech_and4 i_2416(.A(n_3062), .B(n_2560), .C(n_2610), .D(n_2829), .Z(n_3564
		));
	notech_and4 i_2400(.A(n_3107), .B(n_2614), .C(n_2269), .D(n_34075), .Z(n_3567
		));
	notech_and4 i_2404(.A(n_2516), .B(n_2638), .C(n_3567), .D(n_1985), .Z(n_3570
		));
	notech_and4 i_2407(.A(n_3570), .B(n_2709), .C(n_2631), .D(n_3834), .Z(n_3572
		));
	notech_and4 i_2411(.A(n_4058), .B(n_2049), .C(n_2457), .D(n_3572), .Z(n_3574
		));
	notech_and4 i_2408(.A(n_2678), .B(n_2791), .C(n_730), .D(n_1958), .Z(n_3576
		));
	notech_and4 i_2415(.A(n_3576), .B(n_3779), .C(n_3574), .D(n_2099), .Z(n_3579
		));
	notech_and4 i_2420(.A(n_2555), .B(n_3579), .C(n_3564), .D(n_2557), .Z(n_3581
		));
	notech_and4 i_2423(.A(n_2686), .B(n_2675), .C(n_2526), .D(n_3581), .Z(n_3584
		));
	notech_and4 i_2434(.A(n_2903), .B(n_3584), .C(n_2654), .D(n_2702), .Z(n_3586
		));
	notech_and4 i_2435(.A(n_2572), .B(n_2415), .C(n_2309), .D(n_1969), .Z(n_3588
		));
	notech_and4 i_2441(.A(n_2904), .B(n_3588), .C(n_3586), .D(n_2664), .Z(n_3591
		));
	notech_and4 i_1522(.A(n_2572), .B(n_2906), .C(n_2513), .D(n_2918), .Z(n_2921
		));
	notech_or2 i_104577882(.A(n_3957), .B(n_2401), .Z(n_208153600));
	notech_and2 i_186(.A(n_2689), .B(n_2501), .Z(n_3957));
	notech_ao3 i_117077881(.A(n_34009), .B(n_34006), .C(n_3277), .Z(n_207953599
		));
	notech_nao3 i_23111370(.A(n_59539), .B(n_2397), .C(n_2282), .Z(n_1984)
		);
	notech_or4 i_860(.A(n_2282), .B(n_2407), .C(n_59580), .D(n_34192), .Z(n_4079
		));
	notech_and2 i_5677869(.A(n_34047), .B(n_34207), .Z(n_1960));
	notech_and4 i_62490(.A(n_2688), .B(n_2684), .C(n_2662), .D(n_1996), .Z(n_4024
		));
	notech_nor2 i_14(.A(n_2182), .B(n_2185), .Z(n_3971));
	notech_nao3 i_448(.A(modrm[5]), .B(n_34007), .C(n_2325), .Z(n_4027));
	notech_or4 i_23110599(.A(n_2311), .B(n_59539), .C(n_59528), .D(n_34136),
		 .Z(n_4047));
	notech_or2 i_462(.A(n_3957), .B(n_2355), .Z(n_4007));
	notech_or4 i_23111055(.A(n_2383), .B(n_2486), .C(n_2290), .D(n_2292), .Z
		(n_4055));
	notech_and2 i_28477850(.A(n_4022), .B(n_34072), .Z(n_1114));
	notech_or4 i_409(.A(n_2292), .B(n_59548), .C(n_59539), .D(n_34151), .Z(n_4022
		));
	notech_nor2 i_23111358(.A(n_2299), .B(n_2339), .Z(n_4088));
	notech_nor2 i_67177848(.A(n_2101), .B(n_2485), .Z(n_204853574));
	notech_or4 i_359(.A(n_59563), .B(n_2313), .C(n_2389), .D(n_2303), .Z(n_4046
		));
	notech_ao4 i_45777839(.A(n_2118), .B(n_2363), .C(n_2278), .D(n_2339), .Z
		(n_1193));
	notech_or4 i_23111355(.A(n_2339), .B(n_59539), .C(n_59528), .D(n_2271), 
		.Z(n_4044));
	notech_or4 i_8(.A(n_2360), .B(n_2280), .C(n_2282), .D(n_2363), .Z(n_4056
		));
	notech_and4 i_1518(.A(n_4017), .B(n_2915), .C(n_2628), .D(n_3996), .Z(n_2918
		));
	notech_and3 i_55877835(.A(n_4031), .B(n_4036), .C(n_1637), .Z(n_696));
	notech_ao3 i_188(.A(n_34009), .B(n_34041), .C(n_2297), .Z(n_4050));
	notech_nand2 i_63977828(.A(n_3107), .B(n_2614), .Z(n_1086));
	notech_and2 i_68877823(.A(n_4048), .B(n_2195), .Z(n_1925));
	notech_or4 i_23110836(.A(n_59563), .B(n_34195), .C(n_34157), .D(n_59539)
		, .Z(n_4048));
	notech_or4 i_853(.A(n_2311), .B(n_59548), .C(n_59516), .D(n_34080), .Z(n_2305
		));
	notech_or4 i_23110824(.A(n_2286), .B(n_2383), .C(n_34195), .D(n_34157), 
		.Z(n_3993));
	notech_ao3 i_23110716(.A(n_59528), .B(n_59516), .C(n_2464), .Z(n_3969)
		);
	notech_and3 i_79577812(.A(n_4064), .B(n_2377), .C(n_4040), .Z(n_1263));
	notech_or4 i_23110830(.A(n_59563), .B(n_2428), .C(n_59580), .D(n_59598),
		 .Z(n_4040));
	notech_and3 i_816(.A(n_2707), .B(n_2598), .C(n_2704), .Z(n_4071));
	notech_and2 i_541(.A(n_2516), .B(n_3733), .Z(n_4070));
	notech_or4 i_38(.A(n_2410), .B(n_2372), .C(n_4090), .D(n_34202), .Z(n_3984
		));
	notech_and4 i_1515(.A(n_2912), .B(n_2709), .C(n_3980), .D(n_3931), .Z(n_2915
		));
	notech_and4 i_337(.A(n_2310), .B(n_34011), .C(n_59634), .D(n_34004), .Z(n_3974
		));
	notech_or2 i_685(.A(n_2400), .B(n_4072), .Z(n_4030));
	notech_or4 i_23110569(.A(n_2286), .B(n_2311), .C(n_34136), .D(n_34206), 
		.Z(n_4093));
	notech_and4 i_1511(.A(n_2285), .B(n_4014), .C(n_3838), .D(n_2909), .Z(n_2912
		));
	notech_nand3 i_1279(.A(n_59528), .B(n_59538), .C(n_34041), .Z(n_4064));
	notech_or4 i_1053(.A(n_59647), .B(n_59634), .C(n_59616), .D(n_2355), .Z(n_4076
		));
	notech_or4 i_23110839(.A(n_59647), .B(n_2382), .C(n_59634), .D(n_59616),
		 .Z(n_4002));
	notech_or4 i_670(.A(n_2214), .B(n_2497), .C(n_34200), .D(n_34201), .Z(n_4086
		));
	notech_nor2 i_10(.A(n_3935), .B(n_2577), .Z(n_3978));
	notech_or4 i_23111052(.A(n_2360), .B(n_59563), .C(n_2333), .D(n_34053), 
		.Z(n_4026));
	notech_or4 i_11(.A(n_2360), .B(n_2280), .C(n_2282), .D(n_1818), .Z(n_4031
		));
	notech_nor2 i_19(.A(n_4090), .B(n_34142), .Z(n_3986));
	notech_ao3 i_255(.A(n_34009), .B(n_34144), .C(n_2101), .Z(n_4060));
	notech_and4 i_1508(.A(n_4013), .B(n_2255), .C(n_34058), .D(n_34033), .Z(n_2909
		));
	notech_and4 i_1519(.A(n_2162), .B(n_2623), .C(n_4082), .D(n_2019), .Z(n_2906
		));
	notech_or4 i_447(.A(n_59564), .B(n_2519), .C(n_59580), .D(n_34192), .Z(n_4014
		));
	notech_and2 i_412(.A(n_2206), .B(n_4028), .Z(n_2124));
	notech_and2 i_330(.A(n_2359), .B(n_2355), .Z(n_4072));
	notech_and4 i_155(.A(n_3967), .B(n_2171), .C(n_2479), .D(n_2014), .Z(n_2904
		));
	notech_and2 i_613(.A(n_3965), .B(n_3994), .Z(n_2903));
	notech_nao3 i_466(.A(n_34202), .B(n_34007), .C(n_2325), .Z(n_4036));
	notech_ao3 i_93(.A(n_3895), .B(adz), .C(n_2348), .Z(n_4001));
	notech_nor2 i_843(.A(n_2382), .B(n_34142), .Z(n_4080));
	notech_or4 i_139(.A(n_2360), .B(n_59564), .C(n_34089), .D(n_1802), .Z(n_4017
		));
	notech_and3 i_1429(.A(n_2516), .B(n_1890), .C(n_2264), .Z(n_2900));
	notech_or4 i_660(.A(n_2410), .B(n_2037), .C(n_3954), .D(modrm[5]), .Z(n_4053
		));
	notech_and2 i_272(.A(n_2400), .B(n_34138), .Z(n_3958));
	notech_nao3 i_526(.A(n_2397), .B(n_34010), .C(n_2276), .Z(n_4013));
	notech_and2 i_17(.A(n_4067), .B(n_34064), .Z(n_2151));
	notech_or2 i_248(.A(n_3836), .B(n_3957), .Z(n_3994));
	notech_and2 i_772(.A(n_2557), .B(n_2555), .Z(n_2899));
	notech_and4 i_177(.A(n_4008), .B(n_2894), .C(n_34031), .D(n_2895), .Z(n_2898
		));
	notech_ao4 i_239(.A(n_2410), .B(n_2403), .C(n_2325), .D(n_2282), .Z(n_2398
		));
	notech_ao3 i_243(.A(n_2380), .B(n_1951), .C(n_34132), .Z(n_1942));
	notech_and3 i_654(.A(n_2709), .B(n_2071), .C(n_2587), .Z(n_1856));
	notech_and4 i_304(.A(n_2379), .B(n_2699), .C(n_2483), .D(n_1870), .Z(n_1865
		));
	notech_and3 i_260(.A(n_34075), .B(n_1921), .C(n_34047), .Z(n_1834));
	notech_nor2 i_481(.A(n_4057), .B(n_34108), .Z(n_1950));
	notech_and2 i_4450(.A(n_3803), .B(n_3982), .Z(n_1014));
	notech_and2 i_4611(.A(n_4031), .B(n_4036), .Z(n_853));
	notech_and4 i_166(.A(n_4055), .B(n_2538), .C(n_2663), .D(n_3059), .Z(n_872
		));
	notech_and3 i_268(.A(n_2216), .B(n_4037), .C(n_4038), .Z(n_738));
	notech_ao4 i_744(.A(n_3957), .B(n_2485), .C(n_34136), .D(n_2519), .Z(n_811
		));
	notech_and2 i_1433(.A(n_2014), .B(n_2305), .Z(n_2895));
	notech_and4 i_3961(.A(n_3838), .B(n_3973), .C(n_3987), .D(n_4029), .Z(n_2894
		));
	notech_and4 i_162(.A(n_3665), .B(n_1915), .C(n_2212), .D(n_1728), .Z(n_2893
		));
	notech_ao3 i_23111247(.A(n_34200), .B(n_34201), .C(n_2113), .Z(n_4091)
		);
	notech_and4 i_384(.A(n_2654), .B(n_2887), .C(n_1951), .D(n_2619), .Z(n_2890
		));
	notech_and2 i_420(.A(n_2384), .B(n_2382), .Z(n_4090));
	notech_ao3 i_136(.A(n_59548), .B(n_59538), .C(n_2464), .Z(n_4089));
	notech_or4 i_15(.A(n_2315), .B(n_2330), .C(n_2214), .D(n_1900), .Z(n_4087
		));
	notech_or4 i_23111364(.A(n_2289), .B(n_2280), .C(n_2338), .D(n_34010), .Z
		(n_4085));
	notech_nand3 i_274(.A(n_2037), .B(n_2287), .C(n_2375), .Z(n_4084));
	notech_or4 i_33(.A(n_2360), .B(n_59563), .C(n_3935), .D(n_34206), .Z(n_4082
		));
	notech_and2 i_238(.A(n_2517), .B(n_2407), .Z(n_3935));
	notech_and4 i_1439(.A(n_2049), .B(n_2500), .C(n_2510), .D(n_34071), .Z(n_2887
		));
	notech_nao3 i_2969(.A(n_59647), .B(n_2272), .C(n_2403), .Z(n_3733));
	notech_or4 i_1256(.A(n_2282), .B(n_2300), .C(n_34195), .D(n_34157), .Z(n_4067
		));
	notech_or4 i_1265(.A(n_2346), .B(n_2302), .C(n_34202), .D(n_2374), .Z(n_4066
		));
	notech_and2 i_331(.A(n_3277), .B(n_2318), .Z(n_4065));
	notech_or4 i_1294(.A(n_2286), .B(n_2311), .C(n_34136), .D(adz), .Z(n_4062
		));
	notech_or2 i_1295(.A(n_2410), .B(n_2403), .Z(n_4061));
	notech_nor2 i_586(.A(n_3836), .B(n_2101), .Z(n_4059));
	notech_and2 i_207(.A(n_2497), .B(n_2359), .Z(n_3836));
	notech_or4 i_62(.A(n_2276), .B(n_1902), .C(n_2316), .D(n_2289), .Z(n_4058
		));
	notech_ao3 i_23110662(.A(n_59647), .B(n_2272), .C(n_2330), .Z(n_4057));
	notech_ao3 i_201(.A(n_34009), .B(n_34041), .C(n_2275), .Z(n_4054));
	notech_and3 i_355(.A(n_3777), .B(n_4046), .C(n_4034), .Z(n_2884));
	notech_and2 i_332(.A(n_2485), .B(n_2401), .Z(n_3954));
	notech_ao3 i_848(.A(n_34010), .B(n_2296), .C(n_2393), .Z(n_4052));
	notech_or4 i_235(.A(n_2289), .B(n_2338), .C(n_2271), .D(n_2280), .Z(n_4051
		));
	notech_and2 i_487(.A(n_3777), .B(n_4046), .Z(n_2883));
	notech_or2 i_368(.A(n_2285), .B(n_2128), .Z(n_4049));
	notech_ao3 i_23110827(.A(n_59616), .B(n_2324), .C(n_2368), .Z(n_4045));
	notech_or2 i_859(.A(n_2278), .B(n_2337), .Z(n_4043));
	notech_or4 i_669(.A(n_2360), .B(n_59563), .C(n_2486), .D(n_34053), .Z(n_4041
		));
	notech_or2 i_1025(.A(n_2285), .B(n_2095), .Z(n_4038));
	notech_or2 i_35(.A(n_1819), .B(n_2285), .Z(n_4037));
	notech_nor2 i_216(.A(n_2485), .B(n_2215), .Z(n_4035));
	notech_or4 i_25(.A(n_59563), .B(n_2313), .C(n_2389), .D(n_2291), .Z(n_4034
		));
	notech_ao3 i_31(.A(n_34009), .B(n_2349), .C(n_2297), .Z(n_4033));
	notech_or4 i_36(.A(n_2348), .B(n_2360), .C(n_2282), .D(n_1812), .Z(n_4032
		));
	notech_or4 i_23110623(.A(n_2292), .B(n_59548), .C(n_59538), .D(n_34054),
		 .Z(n_4029));
	notech_nand3 i_212(.A(n_34010), .B(n_2530), .C(n_34192), .Z(n_4028));
	notech_or4 i_123(.A(n_2469), .B(n_34145), .C(n_34206), .D(n_34130), .Z(n_4025
		));
	notech_ao3 i_680(.A(modrm[2]), .B(n_2271), .C(n_2564), .Z(n_4023));
	notech_or4 i_1109(.A(n_2347), .B(n_2289), .C(n_3963), .D(n_34196), .Z(n_4020
		));
	notech_and2 i_343(.A(n_34136), .B(n_34080), .Z(n_3963));
	notech_or4 i_23111382(.A(n_2289), .B(n_34089), .C(n_2284), .D(n_2271), .Z
		(n_4019));
	notech_and4 i_23011414(.A(emul), .B(fpu), .C(n_34204), .D(n_2469), .Z(n_4018
		));
	notech_nao3 i_318(.A(n_34009), .B(n_34013), .C(n_2101), .Z(n_4016));
	notech_nor2 i_388(.A(n_3958), .B(n_4072), .Z(n_4015));
	notech_and4 i_1404(.A(n_2834), .B(n_2880), .C(n_2009), .D(n_2010), .Z(n_2881
		));
	notech_and4 i_1403(.A(n_1920), .B(n_2847), .C(n_1870), .D(n_34098), .Z(n_2880
		));
	notech_and4 i_27(.A(emul), .B(fpu), .C(n_34204), .D(n_34008), .Z(n_4011)
		);
	notech_and3 i_23011426(.A(cpl[1]), .B(cpl[0]), .C(ipg_fault), .Z(n_4010)
		);
	notech_and2 i_20(.A(n_34008), .B(ipg_fault), .Z(n_4009));
	notech_or4 i_1117(.A(n_2410), .B(n_2037), .C(n_34202), .D(n_2401), .Z(n_4008
		));
	notech_ao3 i_249(.A(n_59647), .B(n_2272), .C(n_2381), .Z(n_4006));
	notech_nand3 i_133(.A(n_3895), .B(n_59616), .C(n_2324), .Z(n_4005));
	notech_nand2 i_407(.A(n_2330), .B(n_2381), .Z(n_3895));
	notech_or4 i_464(.A(n_59563), .B(n_2519), .C(n_59580), .D(n_59598), .Z(n_4004
		));
	notech_nor2 i_141(.A(n_2244), .B(n_2523), .Z(n_4003));
	notech_and2 i_411(.A(n_2485), .B(n_2497), .Z(n_3845));
	notech_or4 i_217(.A(n_2403), .B(n_2316), .C(n_2311), .D(n_2290), .Z(n_3998
		));
	notech_nao3 i_668(.A(n_34011), .B(adz), .C(n_2519), .Z(n_3996));
	notech_or4 i_1399(.A(n_34160), .B(n_34110), .C(n_2875), .D(n_34114), .Z(n_2878
		));
	notech_or4 i_23111067(.A(n_2289), .B(n_2325), .C(n_2271), .D(n_34136), .Z
		(n_3992));
	notech_or4 i_229(.A(n_2348), .B(n_2360), .C(n_2282), .D(n_2331), .Z(n_3991
		));
	notech_nor2 i_538(.A(n_2278), .B(n_2393), .Z(n_3990));
	notech_or4 i_231(.A(n_59563), .B(n_2316), .C(n_2389), .D(n_2291), .Z(n_3987
		));
	notech_ao3 i_23111121(.A(n_59516), .B(n_59548), .C(n_2318), .Z(n_3985)
		);
	notech_nao3 i_285(.A(n_34009), .B(n_34141), .C(n_2101), .Z(n_3982));
	notech_or4 i_42(.A(n_2311), .B(n_3963), .C(n_59527), .D(n_59516), .Z(n_3981
		));
	notech_or4 i_16(.A(n_59563), .B(n_3935), .C(n_2283), .D(n_34206), .Z(n_3980
		));
	notech_or4 i_125(.A(n_2360), .B(n_59563), .C(n_3935), .D(adz), .Z(n_3979
		));
	notech_or4 i_370(.A(n_2290), .B(n_2292), .C(n_2383), .D(n_2333), .Z(n_3977
		));
	notech_or4 i_498(.A(n_2360), .B(n_59563), .C(n_2325), .D(n_2299), .Z(n_3975
		));
	notech_nao3 i_2992(.A(modrm[2]), .B(n_2530), .C(n_34010), .Z(n_3973));
	notech_or4 i_51(.A(n_2410), .B(n_2373), .C(n_4090), .D(n_34202), .Z(n_3972
		));
	notech_or4 i_23110551(.A(n_2360), .B(n_59563), .C(n_2289), .D(n_2410), .Z
		(n_3970));
	notech_ao3 i_23110686(.A(n_59647), .B(n_2272), .C(n_2368), .Z(n_3968));
	notech_or4 i_338(.A(n_59563), .B(n_2316), .C(n_34089), .D(n_2303), .Z(n_3967
		));
	notech_or4 i_128(.A(n_34089), .B(n_59527), .C(n_59516), .D(n_34080), .Z(n_3965
		));
	notech_or4 i_23110554(.A(n_59564), .B(n_2621), .C(n_59598), .D(n_34193),
		 .Z(n_3964));
	notech_and2 i_147(.A(n_3867), .B(n_1875), .Z(n_2380));
	notech_or4 i_1297(.A(n_59527), .B(n_59516), .C(adz), .D(n_34145), .Z(n_3867
		));
	notech_and2 i_3098(.A(n_4062), .B(n_4093), .Z(n_2366));
	notech_ao3 i_30(.A(n_34193), .B(n_34192), .C(n_59564), .Z(n_2354));
	notech_ao3 i_37(.A(n_34193), .B(n_59598), .C(n_59564), .Z(n_2369));
	notech_nand2 i_3157(.A(n_2327), .B(n_34043), .Z(n_2307));
	notech_or4 i_1392(.A(n_34126), .B(n_34156), .C(n_2873), .D(n_34100), .Z(n_2875
		));
	notech_and2 i_415(.A(n_2286), .B(n_2290), .Z(n_3961));
	notech_ao3 i_256(.A(n_2385), .B(n_34202), .C(n_2410), .Z(n_3959));
	notech_ao3 i_89(.A(n_34200), .B(modrm[4]), .C(n_2214), .Z(n_2210));
	notech_or4 i_3282(.A(n_2386), .B(n_59548), .C(n_59516), .D(n_34195), .Z(n_2182
		));
	notech_or4 i_3297(.A(n_2386), .B(n_59527), .C(n_59516), .D(n_34195), .Z(n_2167
		));
	notech_nand2 i_3299(.A(n_34077), .B(n_34042), .Z(n_2165));
	notech_nand3 i_1388(.A(n_2538), .B(n_2111), .C(n_2872), .Z(n_2873));
	notech_or4 i_110(.A(n_2280), .B(n_2282), .C(n_59598), .D(n_34193), .Z(n_2118
		));
	notech_or4 i_3446(.A(n_59527), .B(n_59516), .C(n_2271), .D(n_34158), .Z(n_2018
		));
	notech_and4 i_1384(.A(n_1815), .B(n_4005), .C(n_2870), .D(n_2789), .Z(n_2872
		));
	notech_nor2 i_23111337(.A(n_2564), .B(n_2271), .Z(n_1987));
	notech_and2 i_12(.A(n_4025), .B(n_34074), .Z(n_1953));
	notech_and4 i_23110674(.A(adz), .B(n_2296), .C(n_2469), .D(n_2466), .Z(n_3950
		));
	notech_and4 i_1381(.A(n_2171), .B(n_2867), .C(n_2857), .D(n_2022), .Z(n_2870
		));
	notech_and3 i_3727(.A(n_3996), .B(n_2579), .C(n_4082), .Z(n_1737));
	notech_and4 i_1377(.A(n_1656), .B(n_2627), .C(n_2863), .D(n_1623), .Z(n_2867
		));
	notech_nand3 i_699(.A(n_4031), .B(n_4056), .C(n_2611), .Z(n_3956));
	notech_and2 i_3849(.A(n_3838), .B(n_4028), .Z(n_1615));
	notech_nand3 i_198(.A(n_34010), .B(n_34192), .C(n_2536), .Z(n_3838));
	notech_and4 i_3919(.A(n_2579), .B(n_1970), .C(n_3998), .D(n_34075), .Z(n_1545
		));
	notech_and2 i_72(.A(n_2063), .B(n_2969), .Z(n_3955));
	notech_or4 i_861(.A(n_59564), .B(n_2865), .C(n_59598), .D(n_34193), .Z(n_3803
		));
	notech_and2 i_4744(.A(n_3739), .B(n_2195), .Z(n_720));
	notech_or4 i_467(.A(n_59643), .B(n_59634), .C(n_59616), .D(n_2401), .Z(n_3739
		));
	notech_or2 i_273(.A(n_1858), .B(n_3963), .Z(n_3880));
	notech_and3 i_5210(.A(n_1829), .B(n_1828), .C(n_4084), .Z(n_254));
	notech_nand3 i_4(.A(n_59643), .B(n_59634), .C(n_59616), .Z(n_2410));
	notech_or4 i_1350(.A(n_2347), .B(n_2244), .C(n_34196), .D(adz), .Z(n_2865
		));
	notech_nand3 i_60(.A(n_59528), .B(n_59538), .C(n_34010), .Z(n_2302));
	notech_nand3 i_65(.A(n_59548), .B(n_59538), .C(n_34010), .Z(n_2275));
	notech_nao3 i_23(.A(n_34192), .B(n_59580), .C(n_59564), .Z(n_2383));
	notech_or4 i_18(.A(n_2372), .B(n_2214), .C(n_2330), .D(n_2504), .Z(n_3931
		));
	notech_and2 i_21(.A(n_34207), .B(n_1919), .Z(n_1951));
	notech_and2 i_22(.A(n_223496909), .B(n_1792), .Z(n_2017));
	notech_and3 i_24(.A(n_59647), .B(n_34196), .C(n_34195), .Z(n_2397));
	notech_nand3 i_61(.A(n_59516), .B(n_59548), .C(n_34010), .Z(n_2278));
	notech_and3 i_76(.A(n_59528), .B(n_59516), .C(n_34010), .Z(n_3908));
	notech_ao4 i_26(.A(n_2278), .B(n_2458), .C(n_2455), .D(n_34053), .Z(n_2123
		));
	notech_and2 i_29(.A(n_2141), .B(n_4013), .Z(n_2065));
	notech_nand2 i_74(.A(opz[1]), .B(n_2322), .Z(n_2320));
	notech_and2 i_34(.A(n_4031), .B(n_4056), .Z(n_2116));
	notech_and4 i_1374(.A(n_3964), .B(n_4004), .C(n_2860), .D(n_2676), .Z(n_2863
		));
	notech_and2 i_53(.A(n_2192), .B(n_4017), .Z(n_2176));
	notech_and2 i_57(.A(n_2071), .B(n_1835), .Z(n_2171));
	notech_and3 i_58(.A(n_2233), .B(n_1938), .C(n_4079), .Z(n_2049));
	notech_and3 i_80(.A(n_2629), .B(n_34060), .C(n_34058), .Z(n_2357));
	notech_and4 i_1371(.A(n_2435), .B(n_3998), .C(n_2008), .D(n_2630), .Z(n_2860
		));
	notech_nand3 i_97(.A(n_2062), .B(adz), .C(n_34011), .Z(n_3890));
	notech_nand3 i_122(.A(n_34077), .B(n_34042), .C(n_34076), .Z(n_2164));
	notech_or4 i_167(.A(n_59564), .B(n_2316), .C(n_34089), .D(n_2291), .Z(n_3876
		));
	notech_ao4 i_130(.A(n_2278), .B(n_2346), .C(n_2275), .D(n_2393), .Z(n_1958
		));
	notech_or4 i_131(.A(fpu), .B(twobyte), .C(ipg_fault), .D(op[7]), .Z(n_2403
		));
	notech_and4 i_135(.A(n_2623), .B(n_3964), .C(n_3965), .D(n_2380), .Z(n_2332
		));
	notech_and3 i_146(.A(n_2327), .B(n_34043), .C(n_2305), .Z(n_2304));
	notech_and2 i_160(.A(n_1918), .B(n_1794), .Z(n_1978));
	notech_ao3 i_704(.A(n_4014), .B(n_1921), .C(n_34012), .Z(n_2857));
	notech_and4 i_170(.A(n_3876), .B(n_2609), .C(n_2663), .D(n_2500), .Z(n_901
		));
	notech_and4 i_175(.A(n_1874), .B(n_2702), .C(n_2900), .D(n_34016), .Z(n_1504
		));
	notech_nand2 i_182(.A(n_34201), .B(modrm[3]), .Z(n_2315));
	notech_and4 i_191(.A(n_59647), .B(n_34196), .C(n_59616), .D(n_2369), .Z(n_3846
		));
	notech_and2 i_204(.A(n_3994), .B(n_34045), .Z(n_1999));
	notech_ao4 i_208(.A(n_2290), .B(n_2447), .C(n_34080), .D(n_2448), .Z(n_2327
		));
	notech_and2 i_211(.A(n_2308), .B(n_2294), .Z(n_2058));
	notech_or4 i_469(.A(n_2410), .B(n_2315), .C(n_2382), .D(n_34202), .Z(n_3834
		));
	notech_and2 i_214(.A(n_3996), .B(n_4082), .Z(n_1972));
	notech_and3 i_220(.A(n_4002), .B(n_1797), .C(n_4017), .Z(n_1777));
	notech_and4 i_309(.A(n_2638), .B(n_2014), .C(n_2192), .D(n_34029), .Z(n_2854
		));
	notech_ao4 i_225(.A(n_1879), .B(n_2488), .C(n_2037), .D(n_2489), .Z(n_2024
		));
	notech_and2 i_240(.A(n_4014), .B(n_2005), .Z(n_1624));
	notech_and2 i_241(.A(n_2057), .B(n_1794), .Z(n_1290));
	notech_nor2 i_862(.A(n_2400), .B(n_2098), .Z(n_3820));
	notech_and2 i_252(.A(n_1985), .B(n_34062), .Z(n_1678));
	notech_and4 i_364(.A(n_2394), .B(n_1958), .C(n_2065), .D(n_2285), .Z(n_2852
		));
	notech_and4 i_261(.A(n_2094), .B(n_4026), .C(n_2155), .D(n_1825), .Z(n_497
		));
	notech_and4 i_263(.A(n_2394), .B(n_1958), .C(n_2026), .D(n_2925), .Z(n_1434
		));
	notech_and4 i_265(.A(n_2179), .B(n_3312), .C(n_3179), .D(n_2180), .Z(n_493
		));
	notech_and4 i_267(.A(n_2398), .B(n_1545), .C(n_34057), .D(n_34036), .Z(n_68
		));
	notech_and4 i_270(.A(n_2639), .B(n_3184), .C(n_3179), .D(n_2937), .Z(n_537
		));
	notech_and2 i_271(.A(n_34040), .B(n_34039), .Z(n_2099));
	notech_ao4 i_278(.A(n_2244), .B(n_2523), .C(n_34138), .D(n_2485), .Z(n_2212
		));
	notech_and2 i_279(.A(n_4041), .B(n_1896), .Z(n_2094));
	notech_and3 i_280(.A(n_1993), .B(n_2665), .C(n_2688), .Z(n_1718));
	notech_and3 i_289(.A(n_2046), .B(n_1912), .C(n_1914), .Z(n_1993));
	notech_and2 i_295(.A(n_2136), .B(n_2978), .Z(n_1329));
	notech_and2 i_299(.A(n_3803), .B(n_34073), .Z(n_1623));
	notech_and4 i_477(.A(n_2151), .B(n_2166), .C(n_2588), .D(n_1890), .Z(n_2850
		));
	notech_and4 i_305(.A(n_2678), .B(n_2791), .C(n_1857), .D(n_533), .Z(n_530
		));
	notech_and4 i_1396(.A(n_2707), .B(n_2352), .C(n_2839), .D(n_2844), .Z(n_2847
		));
	notech_and2 i_314(.A(n_3977), .B(n_4086), .Z(n_1332));
	notech_and4 i_323(.A(n_208153600), .B(n_4049), .C(n_34040), .D(n_3981), 
		.Z(n_444));
	notech_and3 i_324(.A(n_2663), .B(n_2183), .C(n_3422), .Z(n_204));
	notech_and2 i_333(.A(n_4032), .B(n_2365), .Z(n_1905));
	notech_ao4 i_341(.A(n_2400), .B(n_3845), .C(n_3958), .D(n_2401), .Z(n_2157
		));
	notech_and4 i_357(.A(n_3996), .B(n_4014), .C(n_4082), .D(n_3980), .Z(n_1970
		));
	notech_or4 i_360(.A(n_59564), .B(n_2316), .C(n_2389), .D(n_2303), .Z(n_3779
		));
	notech_or4 i_406(.A(n_2389), .B(n_2290), .C(n_2292), .D(n_34080), .Z(n_3777
		));
	notech_and4 i_1391(.A(n_2465), .B(n_2198), .C(n_2842), .D(n_2831), .Z(n_2844
		));
	notech_or4 i_367(.A(n_3956), .B(n_34129), .C(n_34097), .D(n_34123), .Z(n_3773
		));
	notech_and3 i_371(.A(n_2157), .B(n_1930), .C(n_2625), .Z(n_1870));
	notech_and4 i_1386(.A(n_4084), .B(n_2377), .C(n_2827), .D(n_1712), .Z(n_2842
		));
	notech_and3 i_379(.A(n_2231), .B(n_1833), .C(n_1936), .Z(n_1780));
	notech_and4 i_381(.A(n_3739), .B(n_2195), .C(n_2264), .D(n_719), .Z(n_717
		));
	notech_mux2 i_391(.S(n_59598), .A(modrm[0]), .B(modrm[3]), .Z(n_3763));
	notech_nor2 i_395(.A(n_2301), .B(n_3908), .Z(n_3761));
	notech_mux2 i_397(.S(n_59598), .A(n_34200), .B(n_34198), .Z(n_3760));
	notech_nao3 i_401(.A(n_59616), .B(n_34202), .C(n_2386), .Z(n_2214));
	notech_and3 i_402(.A(n_223496909), .B(n_1792), .C(n_34050), .Z(n_2015)
		);
	notech_and2 i_413(.A(n_3838), .B(n_3973), .Z(n_2076));
	notech_and3 i_421(.A(n_4062), .B(n_4093), .C(n_34046), .Z(n_2022));
	notech_nao3 i_852(.A(n_2385), .B(n_34141), .C(n_2214), .Z(n_3751));
	notech_and2 i_425(.A(n_3751), .B(n_34074), .Z(n_1526));
	notech_and2 i_428(.A(n_4055), .B(n_1857), .Z(n_2029));
	notech_and2 i_437(.A(n_34065), .B(n_34045), .Z(n_1728));
	notech_ao4 i_440(.A(n_2501), .B(n_2382), .C(n_59564), .D(n_2646), .Z(n_733
		));
	notech_and4 i_310(.A(n_4002), .B(n_2195), .C(n_2414), .D(n_2597), .Z(n_2839
		));
	notech_and2 i_454(.A(n_2073), .B(n_2202), .Z(n_2162));
	notech_and4 i_455(.A(n_3979), .B(n_1970), .C(n_34073), .D(n_1978), .Z(n_1969
		));
	notech_and2 i_474(.A(n_3979), .B(n_3980), .Z(n_1816));
	notech_or4 i_835(.A(n_2214), .B(n_2384), .C(modrm[3]), .D(n_34201), .Z(n_3736
		));
	notech_and2 i_476(.A(n_2587), .B(n_1851), .Z(n_1603));
	notech_nand2 i_479(.A(n_3998), .B(n_34075), .Z(n_1967));
	notech_and4 i_492(.A(n_3967), .B(n_3987), .C(n_1796), .D(n_4029), .Z(n_3728
		));
	notech_or4 i_493(.A(n_59564), .B(n_2286), .C(n_59580), .D(n_34192), .Z(n_2368
		));
	notech_and3 i_501(.A(n_34057), .B(n_34036), .C(n_2305), .Z(n_1924));
	notech_and2 i_508(.A(n_2327), .B(n_4047), .Z(n_1923));
	notech_and4 i_515(.A(n_34063), .B(n_1958), .C(n_2377), .D(n_34044), .Z(n_960
		));
	notech_nao3 i_532(.A(n_34010), .B(n_2375), .C(n_2286), .Z(n_2113));
	notech_and2 i_792(.A(n_2411), .B(n_1603), .Z(n_2834));
	notech_or4 i_536(.A(n_59647), .B(n_2338), .C(n_59616), .D(n_34196), .Z(n_2234
		));
	notech_and2 i_545(.A(n_2216), .B(n_34143), .Z(n_1656));
	notech_and2 i_550(.A(n_2132), .B(n_2789), .Z(n_455));
	notech_and4 i_555(.A(n_4027), .B(n_4036), .C(n_4076), .D(n_2091), .Z(n_894
		));
	notech_and4 i_562(.A(n_2233), .B(n_1938), .C(n_4079), .D(n_4058), .Z(n_2047
		));
	notech_and3 i_567(.A(n_3838), .B(n_3973), .C(n_1798), .Z(n_3697));
	notech_and3 i_692(.A(n_4025), .B(n_34074), .C(n_2357), .Z(n_2831));
	notech_and2 i_606(.A(n_2380), .B(n_34207), .Z(n_1593));
	notech_and3 i_94(.A(n_3992), .B(n_1895), .C(n_1831), .Z(n_2829));
	notech_ao4 i_604(.A(n_2387), .B(n_34140), .C(n_2382), .D(n_34142), .Z(n_2827
		));
	notech_ao4 i_618(.A(n_34136), .B(n_2407), .C(n_2485), .D(n_34138), .Z(n_1306
		));
	notech_and2 i_625(.A(n_3982), .B(n_34043), .Z(n_1537));
	notech_and3 i_634(.A(n_3993), .B(n_4040), .C(n_2103), .Z(n_730));
	notech_and3 i_637(.A(n_3992), .B(n_2123), .C(n_34031), .Z(n_1712));
	notech_and4 i_780(.A(n_1949), .B(n_1796), .C(n_3880), .D(n_34016), .Z(n_2826
		));
	notech_or2 i_658(.A(n_3958), .B(n_2355), .Z(n_3672));
	notech_or4 i_659(.A(n_2316), .B(n_2276), .C(n_2373), .D(n_2333), .Z(n_2052
		));
	notech_or2 i_684(.A(n_2400), .B(n_2359), .Z(n_3665));
	notech_ao4 i_708(.A(n_2400), .B(n_3845), .C(n_34145), .D(n_2286), .Z(n_1543
		));
	notech_or4 i_729(.A(n_4010), .B(n_4018), .C(n_3950), .D(n_4015), .Z(n_1262
		));
	notech_and2 i_736(.A(n_3979), .B(n_4032), .Z(n_861));
	notech_and2 i_748(.A(n_2246), .B(n_1984), .Z(n_520));
	notech_and2 i_750(.A(n_2665), .B(n_2394), .Z(n_719));
	notech_and3 i_751(.A(n_2790), .B(n_1993), .C(n_3105), .Z(n_703));
	notech_ao4 i_753(.A(n_2291), .B(n_34151), .C(n_2118), .D(n_2363), .Z(n_673
		));
	notech_and2 i_755(.A(n_4002), .B(n_4048), .Z(n_2080));
	notech_ao4 i_757(.A(n_2422), .B(n_2384), .C(n_2499), .D(n_2382), .Z(n_574
		));
	notech_and2 i_768(.A(n_1936), .B(n_34036), .Z(n_215));
	notech_and3 i_769(.A(n_4041), .B(n_4036), .C(n_2056), .Z(n_1284));
	notech_and3 i_779(.A(n_3880), .B(n_3374), .C(n_2213), .Z(n_218));
	notech_and2 i_781(.A(n_2206), .B(n_733), .Z(n_709));
	notech_and3 i_782(.A(n_2625), .B(n_3779), .C(n_2073), .Z(n_533));
	notech_and3 i_791(.A(n_3979), .B(n_3980), .C(n_4082), .Z(n_1815));
	notech_or4 i_1318(.A(n_34164), .B(n_2817), .C(n_1998), .D(n_2000), .Z(n_2820
		));
	notech_and3 i_804(.A(n_4055), .B(n_2538), .C(n_3834), .Z(n_1340));
	notech_and3 i_810(.A(n_2166), .B(n_2108), .C(n_2380), .Z(n_466));
	notech_and3 i_812(.A(n_1886), .B(n_2686), .C(n_1887), .Z(n_2246));
	notech_and4 i_813(.A(n_3834), .B(n_2036), .C(n_1924), .D(n_3984), .Z(n_1920
		));
	notech_and3 i_818(.A(n_2025), .B(n_2103), .C(n_4027), .Z(n_1346));
	notech_and4 i_2932(.A(n_4047), .B(n_2091), .C(n_1999), .D(n_34065), .Z(n_1996
		));
	notech_or4 i_1315(.A(n_34105), .B(n_34122), .C(n_34159), .D(n_2814), .Z(n_2817
		));
	notech_nao3 i_1313(.A(n_1678), .B(n_2588), .C(n_2812), .Z(n_2814));
	notech_or4 i_1311(.A(n_1997), .B(n_34134), .C(n_2809), .D(n_2078), .Z(n_2812
		));
	notech_nao3 i_1308(.A(n_3777), .B(n_2808), .C(n_222398896), .Z(n_2809)
		);
	notech_and4 i_1307(.A(n_3665), .B(n_1923), .C(n_2804), .D(n_34070), .Z(n_2808
		));
	notech_and4 i_1304(.A(n_2627), .B(n_1995), .C(n_3965), .D(n_2801), .Z(n_2804
		));
	notech_ao3 i_1300(.A(n_2799), .B(n_2216), .C(n_1933), .Z(n_2801));
	notech_and4 i_1298(.A(n_2516), .B(n_2797), .C(n_3998), .D(n_2794), .Z(n_2799
		));
	notech_and4 i_1292(.A(n_34060), .B(n_34058), .C(n_1990), .D(n_1994), .Z(n_2797
		));
	notech_ao4 i_1290(.A(n_59528), .B(n_2734), .C(n_2140), .D(n_59516), .Z(n_2794
		));
	notech_and2 i_237(.A(n_2791), .B(n_2790), .Z(n_2792));
	notech_ao4 i_486(.A(n_2384), .B(n_34138), .C(n_2403), .D(n_34089), .Z(n_2791
		));
	notech_and2 i_43(.A(n_2789), .B(n_1982), .Z(n_2790));
	notech_and3 i_349(.A(n_1901), .B(n_4087), .C(n_3931), .Z(n_2789));
	notech_or4 i_1262(.A(n_222998902), .B(n_1975), .C(n_1976), .D(n_2782), .Z
		(n_2785));
	notech_nand3 i_1259(.A(n_2780), .B(n_2729), .C(n_222798900), .Z(n_2782)
		);
	notech_and4 i_1257(.A(n_2778), .B(n_2212), .C(n_34031), .D(n_2532), .Z(n_2780
		));
	notech_and4 i_1254(.A(n_2765), .B(n_1978), .C(n_2136), .D(n_2777), .Z(n_2778
		));
	notech_and4 i_1253(.A(n_2192), .B(n_2775), .C(n_2744), .D(n_2305), .Z(n_2777
		));
	notech_and4 i_1248(.A(n_1877), .B(n_2772), .C(n_3996), .D(n_34042), .Z(n_2775
		));
	notech_and4 i_1245(.A(n_2768), .B(n_3993), .C(n_2771), .D(n_34075), .Z(n_2772
		));
	notech_ao4 i_1244(.A(n_2458), .B(n_2299), .C(n_2383), .D(n_2621), .Z(n_2771
		));
	notech_ao4 i_1240(.A(n_2734), .B(n_34192), .C(n_2140), .D(n_34195), .Z(n_2768
		));
	notech_and3 i_173(.A(n_2216), .B(n_2733), .C(n_2730), .Z(n_2765));
	notech_and4 i_3740(.A(n_223496909), .B(n_1792), .C(n_2151), .D(n_34050),
		 .Z(n_2760));
	notech_and4 i_226(.A(n_34065), .B(n_34045), .C(n_2091), .D(n_3994), .Z(n_2759
		));
	notech_and2 i_478(.A(n_1993), .B(n_2665), .Z(n_2757));
	notech_and4 i_1213(.A(n_2751), .B(n_222798900), .C(n_2729), .D(n_1955), 
		.Z(n_2754));
	notech_and4 i_1210(.A(n_34148), .B(n_2749), .C(n_34075), .D(n_1954), .Z(n_2751
		));
	notech_and4 i_1208(.A(n_1930), .B(n_2741), .C(n_2747), .D(n_1737), .Z(n_2749
		));
	notech_and4 i_1206(.A(n_1949), .B(n_2744), .C(n_1952), .D(n_2743), .Z(n_2747
		));
	notech_and2 i_251(.A(n_1932), .B(n_34106), .Z(n_2744));
	notech_and2 i_138(.A(n_2192), .B(n_2305), .Z(n_2743));
	notech_and4 i_1203(.A(n_2730), .B(n_2731), .C(n_3965), .D(n_2739), .Z(n_2741
		));
	notech_and4 i_1200(.A(n_3993), .B(n_3992), .C(n_2736), .D(n_3980), .Z(n_2739
		));
	notech_and3 i_1194(.A(n_2733), .B(n_2234), .C(n_1947), .Z(n_2736));
	notech_ao4 i_218(.A(n_2403), .B(n_2389), .C(n_59564), .D(n_2646), .Z(n_2734
		));
	notech_ao4 i_543(.A(n_34080), .B(n_2446), .C(n_2325), .D(n_2282), .Z(n_2733
		));
	notech_ao4 i_1196(.A(n_2166), .B(n_34175), .C(n_2290), .D(n_2464), .Z(n_2731
		));
	notech_ao4 i_696(.A(n_2318), .B(n_2286), .C(n_34080), .D(n_2519), .Z(n_2730
		));
	notech_and4 i_157(.A(n_4084), .B(n_2377), .C(n_3751), .D(n_2727), .Z(n_2729
		));
	notech_ao4 i_1154(.A(n_2118), .B(n_2027), .C(n_2362), .D(n_2331), .Z(n_2727
		));
	notech_and4 i_1173(.A(n_34063), .B(n_1780), .C(n_2395), .D(n_2414), .Z(n_2726
		));
	notech_and2 i_485(.A(n_4002), .B(n_1797), .Z(n_2723));
	notech_and3 i_300(.A(n_3967), .B(n_2171), .C(n_2479), .Z(n_2722));
	notech_and4 i_1182(.A(n_2141), .B(n_4013), .C(n_2015), .D(n_1941), .Z(n_2719
		));
	notech_and4 i_348(.A(n_2195), .B(n_2714), .C(n_2611), .D(n_2713), .Z(n_2717
		));
	notech_ao4 i_1177(.A(n_2384), .B(n_1937), .C(n_2052), .D(n_2331), .Z(n_2714
		));
	notech_and2 i_701(.A(n_4016), .B(n_3972), .Z(n_2713));
	notech_and2 i_452(.A(n_1798), .B(n_2111), .Z(n_2709));
	notech_and4 i_387(.A(n_2190), .B(n_3973), .C(n_2463), .D(n_2675), .Z(n_2707
		));
	notech_and2 i_646(.A(n_2703), .B(n_2543), .Z(n_2704));
	notech_and4 i_473(.A(n_1873), .B(n_2555), .C(n_1874), .D(n_2702), .Z(n_2703
		));
	notech_and2 i_233(.A(n_1800), .B(n_2563), .Z(n_2702));
	notech_and4 i_1127(.A(n_2417), .B(n_2695), .C(n_2198), .D(n_2696), .Z(n_2699
		));
	notech_and4 i_1124(.A(n_2073), .B(n_4067), .C(n_2202), .D(n_34064), .Z(n_2696
		));
	notech_and2 i_399(.A(n_1796), .B(n_4029), .Z(n_2695));
	notech_and2 i_566(.A(n_2157), .B(n_1930), .Z(n_2694));
	notech_and3 i_3466(.A(n_3994), .B(n_34045), .C(n_34065), .Z(n_2690));
	notech_or4 i_101(.A(n_2386), .B(n_2037), .C(n_34195), .D(n_34202), .Z(n_2689
		));
	notech_and2 i_288(.A(n_2246), .B(n_2264), .Z(n_2688));
	notech_ao4 i_376(.A(n_2553), .B(n_2685), .C(n_2557), .D(n_2037), .Z(n_2686
		));
	notech_nand2 i_936(.A(n_1885), .B(modrm[1]), .Z(n_2685));
	notech_and4 i_711(.A(n_2681), .B(n_2675), .C(n_2665), .D(n_2664), .Z(n_2684
		));
	notech_and4 i_1021(.A(n_2179), .B(n_2678), .C(n_2457), .D(n_2022), .Z(n_2681
		));
	notech_and3 i_193(.A(n_2676), .B(n_2189), .C(n_2190), .Z(n_2678));
	notech_and2 i_54(.A(n_2188), .B(n_1907), .Z(n_2676));
	notech_and4 i_358(.A(n_4055), .B(n_1857), .C(n_3977), .D(n_2673), .Z(n_2675
		));
	notech_and4 i_877(.A(n_1855), .B(n_1854), .C(n_2668), .D(n_2238), .Z(n_2673
		));
	notech_ao4 i_137(.A(n_2667), .B(n_2300), .C(n_2666), .D(n_2292), .Z(n_2668
		));
	notech_nand2 i_868(.A(n_2530), .B(n_59598), .Z(n_2667));
	notech_nand2 i_867(.A(n_34192), .B(n_2536), .Z(n_2666));
	notech_and2 i_758(.A(n_2024), .B(n_1911), .Z(n_2665));
	notech_and2 i_614(.A(n_2663), .B(n_2352), .Z(n_2664));
	notech_ao4 i_52(.A(n_2291), .B(n_2052), .C(n_2278), .D(n_2337), .Z(n_2663
		));
	notech_and4 i_1111(.A(n_2484), .B(n_2549), .C(n_2483), .D(n_2661), .Z(n_2662
		));
	notech_and4 i_1108(.A(n_2658), .B(n_2619), .C(n_2607), .D(n_2567), .Z(n_2661
		));
	notech_and4 i_1100(.A(n_2654), .B(n_2157), .C(n_2650), .D(n_2656), .Z(n_2658
		));
	notech_and2 i_602(.A(n_2655), .B(n_4025), .Z(n_2656));
	notech_ao4 i_356(.A(n_2391), .B(n_2303), .C(n_2291), .D(n_34054), .Z(n_2655
		));
	notech_and2 i_293(.A(n_2030), .B(n_3991), .Z(n_2654));
	notech_and4 i_1093(.A(n_2648), .B(n_2643), .C(n_2304), .D(n_2620), .Z(n_2650
		));
	notech_and4 i_383(.A(n_4002), .B(n_4048), .C(n_2076), .D(n_34031), .Z(n_2648
		));
	notech_or4 i_997(.A(n_59647), .B(n_59634), .C(n_34195), .D(n_59538), .Z(n_2646
		));
	notech_and4 i_1087(.A(n_2625), .B(n_2634), .C(n_2332), .D(n_2641), .Z(n_2643
		));
	notech_and4 i_1084(.A(n_4058), .B(n_2049), .C(n_2639), .D(n_3981), .Z(n_2641
		));
	notech_and2 i_242(.A(n_2638), .B(n_2014), .Z(n_2639));
	notech_ao4 i_215(.A(n_2325), .B(n_2384), .C(n_2383), .D(n_2428), .Z(n_2638
		));
	notech_and2 i_616(.A(n_2233), .B(n_1938), .Z(n_2637));
	notech_and4 i_1081(.A(n_2631), .B(n_2628), .C(n_2357), .D(n_34074), .Z(n_2634
		));
	notech_and3 i_302(.A(n_2433), .B(n_2140), .C(n_4064), .Z(n_2631));
	notech_and2 i_569(.A(n_2433), .B(n_2140), .Z(n_2630));
	notech_nor2 i_426(.A(n_4010), .B(n_4018), .Z(n_2629));
	notech_and3 i_774(.A(n_3993), .B(n_4040), .C(n_3733), .Z(n_2628));
	notech_and2 i_410(.A(n_3993), .B(n_4040), .Z(n_2627));
	notech_and2 i_134(.A(n_1877), .B(n_1831), .Z(n_2625));
	notech_and2 i_45(.A(n_34057), .B(n_34036), .Z(n_2623));
	notech_or4 i_923(.A(n_2386), .B(n_34195), .C(n_59548), .D(n_59539), .Z(n_2621
		));
	notech_and2 i_509(.A(n_3987), .B(n_4029), .Z(n_2620));
	notech_and4 i_36696642(.A(n_2611), .B(n_2379), .C(n_2614), .D(n_2616), .Z
		(n_2619));
	notech_and4 i_978(.A(n_4027), .B(n_4036), .C(n_34040), .D(n_34039), .Z(n_2616
		));
	notech_and2 i_783(.A(n_4027), .B(n_4036), .Z(n_2615));
	notech_and3 i_430(.A(n_4041), .B(n_1896), .C(n_4026), .Z(n_2614));
	notech_and4 i_196(.A(n_4044), .B(n_2609), .C(n_2108), .D(n_34072), .Z(n_2611
		));
	notech_and4 i_802(.A(n_4044), .B(n_4051), .C(n_34072), .D(n_4085), .Z(n_2610
		));
	notech_and2 i_458(.A(n_4051), .B(n_4085), .Z(n_2609));
	notech_and4 i_1102(.A(n_2572), .B(n_1969), .C(n_2605), .D(n_2309), .Z(n_2607
		));
	notech_and4 i_63(.A(n_2591), .B(n_2602), .C(n_2588), .D(n_2587), .Z(n_2605
		));
	notech_and4 i_1076(.A(n_3931), .B(n_2598), .C(n_2171), .D(n_2601), .Z(n_2602
		));
	notech_and3 i_1075(.A(n_2192), .B(n_4017), .C(n_2195), .Z(n_2601));
	notech_and3 i_199(.A(n_2103), .B(n_2159), .C(n_1851), .Z(n_2598));
	notech_and2 i_830(.A(n_2103), .B(n_2159), .Z(n_2597));
	notech_or4 i_823(.A(n_59564), .B(n_2486), .C(n_59580), .D(n_34192), .Z(n_2596
		));
	notech_or4 i_863(.A(n_2302), .B(n_59616), .C(n_34157), .D(modrm[5]), .Z(n_2594
		));
	notech_and4 i_787(.A(n_2162), .B(n_34077), .C(n_34042), .D(n_34076), .Z(n_2591
		));
	notech_and3 i_598(.A(n_3970), .B(n_1806), .C(n_34047), .Z(n_2588));
	notech_and2 i_152(.A(n_1825), .B(n_2070), .Z(n_2587));
	notech_or4 i_1069(.A(n_59564), .B(n_2283), .C(n_34089), .D(n_34202), .Z(n_2586
		));
	notech_and3 i_223(.A(n_3979), .B(n_34073), .C(n_1978), .Z(n_2579));
	notech_or4 i_910(.A(n_59564), .B(n_34193), .C(n_34192), .D(adz), .Z(n_2577
		));
	notech_or4 i_663(.A(n_59647), .B(n_59616), .C(n_34196), .D(n_34130), .Z(n_2574
		));
	notech_and4 i_378(.A(n_1984), .B(n_1801), .C(n_4019), .D(n_34143), .Z(n_2572
		));
	notech_and2 i_517(.A(n_1984), .B(n_1801), .Z(n_2571));
	notech_and2 i_3478(.A(n_4019), .B(n_34143), .Z(n_2569));
	notech_and3 i_377(.A(n_2565), .B(n_2563), .C(n_2562), .Z(n_2567));
	notech_and3 i_759(.A(n_4067), .B(n_2166), .C(n_34064), .Z(n_2565));
	notech_or4 i_499(.A(n_59647), .B(n_2282), .C(n_59634), .D(n_34195), .Z(n_2564
		));
	notech_ao4 i_442(.A(n_2494), .B(n_2315), .C(n_2489), .D(n_2373), .Z(n_2563
		));
	notech_and4 i_723(.A(n_1873), .B(n_2555), .C(n_1874), .D(n_1800), .Z(n_2562
		));
	notech_or4 i_108(.A(n_2497), .B(n_2333), .C(modrm[1]), .D(modrm[0]), .Z(n_2560
		));
	notech_or4 i_109(.A(n_2497), .B(n_2333), .C(modrm[1]), .D(n_34198), .Z(n_2557
		));
	notech_and2 i_291(.A(n_1869), .B(n_1871), .Z(n_2555));
	notech_or2 i_496(.A(n_2497), .B(n_2333), .Z(n_2553));
	notech_and4 i_1101(.A(n_2510), .B(n_2500), .C(n_2547), .D(n_2498), .Z(n_2549
		));
	notech_and4 i_1095(.A(n_2534), .B(n_2522), .C(n_2526), .D(n_2545), .Z(n_2547
		));
	notech_and4 i_1088(.A(n_2538), .B(n_2111), .C(n_3982), .D(n_2543), .Z(n_2545
		));
	notech_and2 i_433(.A(n_3880), .B(n_34016), .Z(n_2543));
	notech_nor2 i_832(.A(n_2486), .B(n_2288), .Z(n_2542));
	notech_ao3 i_829(.A(modrm[2]), .B(n_2287), .C(n_2333), .Z(n_2541));
	notech_and3 i_608(.A(n_1798), .B(n_1796), .C(n_2111), .Z(n_2539));
	notech_and2 i_190(.A(n_1798), .B(n_1796), .Z(n_2538));
	notech_and4 i_84(.A(n_59528), .B(n_2431), .C(n_34193), .D(n_34202), .Z(n_2536
		));
	notech_and4 i_362(.A(n_2206), .B(n_4028), .C(n_2532), .D(n_3777), .Z(n_2534
		));
	notech_and4 i_638(.A(n_2206), .B(n_4028), .C(n_3992), .D(n_2123), .Z(n_2533
		));
	notech_and2 i_423(.A(n_3992), .B(n_2123), .Z(n_2532));
	notech_nand2 i_963(.A(n_34192), .B(n_34010), .Z(n_2531));
	notech_and4 i_83(.A(n_2431), .B(n_59528), .C(n_34193), .D(modrm[5]), .Z(n_2530
		));
	notech_and4 i_315(.A(n_3665), .B(n_2216), .C(n_3672), .D(n_2212), .Z(n_2526
		));
	notech_nand3 i_833(.A(n_2310), .B(n_34011), .C(n_59634), .Z(n_2523));
	notech_and4 i_298(.A(n_4004), .B(n_2398), .C(n_2513), .D(n_2518), .Z(n_2522
		));
	notech_or4 i_187(.A(n_59647), .B(n_2244), .C(n_59616), .D(n_34196), .Z(n_2519
		));
	notech_and2 i_713(.A(n_2516), .B(n_1890), .Z(n_2518));
	notech_or4 i_495(.A(n_59647), .B(n_2289), .C(n_59616), .D(n_34196), .Z(n_2517
		));
	notech_and2 i_903(.A(n_2515), .B(n_2032), .Z(n_2516));
	notech_or4 i_580(.A(n_2279), .B(n_59564), .C(n_34195), .D(n_59539), .Z(n_2515
		));
	notech_and2 i_703(.A(n_2234), .B(n_4005), .Z(n_2513));
	notech_and2 i_392(.A(n_2289), .B(n_34130), .Z(n_2512));
	notech_and4 i_380(.A(n_1901), .B(n_4087), .C(n_2198), .D(n_3972), .Z(n_2510
		));
	notech_or4 i_991(.A(n_2410), .B(modrm[3]), .C(modrm[4]), .D(modrm[5]), .Z
		(n_2505));
	notech_xor2 i_432(.A(n_34203), .B(modrm[7]), .Z(n_2504));
	notech_or4 i_90(.A(n_2410), .B(modrm[3]), .C(n_34201), .D(n_34202), .Z(n_2501
		));
	notech_and2 i_213(.A(n_3834), .B(n_3984), .Z(n_2500));
	notech_or4 i_87(.A(n_2386), .B(n_2315), .C(n_34195), .D(n_34202), .Z(n_2499
		));
	notech_and2 i_771(.A(n_1993), .B(n_1915), .Z(n_2498));
	notech_or4 i_48(.A(n_2329), .B(n_2292), .C(n_59548), .D(n_59539), .Z(n_2497
		));
	notech_and2 i_418(.A(n_2373), .B(n_2372), .Z(n_2495));
	notech_or4 i_578(.A(n_2486), .B(n_2485), .C(modrm[1]), .D(n_34198), .Z(n_2494
		));
	notech_and2 i_403(.A(n_34200), .B(n_34201), .Z(n_2492));
	notech_or4 i_885(.A(n_59616), .B(n_34157), .C(n_34202), .D(modrm[1]), .Z
		(n_2490));
	notech_or2 i_106(.A(n_2488), .B(modrm[0]), .Z(n_2489));
	notech_or4 i_836(.A(n_2325), .B(n_2485), .C(n_34202), .D(n_34199), .Z(n_2488
		));
	notech_or4 i_40(.A(n_59647), .B(n_59634), .C(n_59616), .D(n_34202), .Z(n_2486
		));
	notech_or4 i_49(.A(n_2329), .B(n_2300), .C(n_59548), .D(n_59539), .Z(n_2485
		));
	notech_and4 i_799(.A(n_1919), .B(n_3998), .C(n_34071), .D(n_34075), .Z(n_2484
		));
	notech_and4 i_319(.A(n_3967), .B(n_2480), .C(n_2479), .D(n_2415), .Z(n_2483
		));
	notech_ao4 i_129(.A(n_2027), .B(n_2393), .C(n_2346), .D(n_2387), .Z(n_2480
		));
	notech_and2 i_611(.A(n_3876), .B(n_4022), .Z(n_2479));
	notech_nand3 i_803(.A(n_2450), .B(n_2036), .C(n_2474), .Z(n_2475));
	notech_and3 i_795(.A(n_247296910), .B(n_2465), .C(n_1848), .Z(n_2474));
	notech_and3 i_800(.A(n_4025), .B(n_34060), .C(n_34058), .Z(n_247296910)
		);
	notech_and2 i_831(.A(cpl[1]), .B(cpl[0]), .Z(n_2469));
	notech_ao3 i_408(.A(n_59647), .B(n_2272), .C(n_2383), .Z(n_2466));
	notech_and4 i_504(.A(n_3965), .B(n_34077), .C(n_34042), .D(n_34076), .Z(n_2465
		));
	notech_or4 i_530(.A(n_59564), .B(n_34089), .C(n_59580), .D(n_34192), .Z(n_2464
		));
	notech_and4 i_119(.A(n_2189), .B(n_2206), .C(n_2179), .D(n_2457), .Z(n_2463
		));
	notech_or4 i_528(.A(n_59647), .B(n_59634), .C(n_59616), .D(n_34080), .Z(n_2458
		));
	notech_and3 i_316(.A(n_2255), .B(n_1805), .C(n_3975), .Z(n_2457));
	notech_or4 i_99(.A(n_59564), .B(n_59616), .C(n_34157), .D(n_59580), .Z(n_2455
		));
	notech_ao3 i_470(.A(n_3970), .B(n_1806), .C(n_1807), .Z(n_2450));
	notech_nand3 i_150(.A(n_2310), .B(n_59634), .C(n_34004), .Z(n_2448));
	notech_or4 i_849(.A(n_59563), .B(n_2311), .C(n_59580), .D(n_59585), .Z(n_2447
		));
	notech_nao3 i_457(.A(n_59548), .B(n_59539), .C(n_2311), .Z(n_2446));
	notech_or4 i_801(.A(n_34051), .B(n_34134), .C(n_2442), .D(n_3986), .Z(n_2445
		));
	notech_nao3 i_784(.A(n_2440), .B(n_2430), .C(n_1846), .Z(n_2442));
	notech_and4 i_775(.A(n_1843), .B(n_2437), .C(n_2140), .D(n_34075), .Z(n_2440
		));
	notech_and4 i_761(.A(n_2435), .B(n_1960), .C(n_3993), .D(n_2305), .Z(n_2437
		));
	notech_and2 i_44977840(.A(n_2234), .B(n_2398), .Z(n_2435));
	notech_and2 i_69077822(.A(n_3993), .B(n_2305), .Z(n_2434));
	notech_or2 i_250(.A(n_2403), .B(n_2389), .Z(n_2433));
	notech_nor2 i_579(.A(n_59647), .B(n_2403), .Z(n_2431));
	notech_ao4 i_773(.A(n_34193), .B(n_1842), .C(n_2383), .D(n_2428), .Z(n_2430
		));
	notech_or4 i_527(.A(n_59528), .B(n_59516), .C(n_34195), .D(n_34157), .Z(n_2428
		));
	notech_and3 i_674(.A(n_34195), .B(n_2324), .C(n_2369), .Z(n_2427));
	notech_and4 i_636(.A(n_4062), .B(n_4093), .C(n_34046), .D(n_34057), .Z(n_2426
		));
	notech_or4 i_352(.A(n_2386), .B(n_2372), .C(n_59603), .D(n_34202), .Z(n_2422
		));
	notech_and4 i_127(.A(n_59647), .B(n_34196), .C(n_59603), .D(n_2354), .Z(n_2418
		));
	notech_and2 i_594(.A(n_1938), .B(n_1835), .Z(n_2417));
	notech_and3 i_450(.A(n_2137), .B(n_2045), .C(n_2411), .Z(n_2415));
	notech_and2 i_307(.A(n_2137), .B(n_2045), .Z(n_2414));
	notech_and2 i_398(.A(n_2302), .B(n_34152), .Z(n_2413));
	notech_or4 i_194(.A(n_59558), .B(n_2325), .C(n_59598), .D(n_34193), .Z(n_2412
		));
	notech_and3 i_142(.A(n_2231), .B(n_1833), .C(n_2026), .Z(n_2411));
	notech_nao3 i_730(.A(n_34193), .B(n_59598), .C(n_2276), .Z(n_2408));
	notech_or4 i_77(.A(n_59647), .B(n_2290), .C(n_59616), .D(n_34196), .Z(n_2407
		));
	notech_and4 i_246(.A(n_2395), .B(n_2402), .C(n_2392), .D(n_2379), .Z(n_2406
		));
	notech_ao4 i_725(.A(n_2401), .B(n_3958), .C(n_3963), .D(n_2396), .Z(n_2402
		));
	notech_or4 i_67(.A(n_2329), .B(n_59539), .C(n_59528), .D(n_34010), .Z(n_2401
		));
	notech_and2 i_390(.A(n_34142), .B(n_2399), .Z(n_2400));
	notech_or4 i_96(.A(n_2410), .B(n_34200), .C(n_34201), .D(modrm[5]), .Z(n_2399
		));
	notech_or4 i_691(.A(n_59643), .B(n_2299), .C(n_59634), .D(n_59612), .Z(n_2396
		));
	notech_and3 i_434(.A(n_1829), .B(n_1828), .C(n_1958), .Z(n_2395));
	notech_ao4 i_132(.A(n_2297), .B(n_2393), .C(n_2346), .D(n_2299), .Z(n_2394
		));
	notech_or4 i_107(.A(n_2347), .B(n_2313), .C(n_2282), .D(n_34196), .Z(n_2393
		));
	notech_ao4 i_778(.A(n_2391), .B(n_2387), .C(n_34138), .D(n_4090), .Z(n_2392
		));
	notech_and2 i_429(.A(n_34054), .B(n_34140), .Z(n_2391));
	notech_and4 i_100(.A(n_59643), .B(n_34196), .C(n_59612), .D(n_2354), .Z(n_2390
		));
	notech_nand3 i_664(.A(n_59643), .B(n_34196), .C(n_59612), .Z(n_2389));
	notech_and2 i_185(.A(n_2278), .B(n_2299), .Z(n_2387));
	notech_nand2 i_369(.A(n_59643), .B(n_59634), .Z(n_2386));
	notech_nand2 i_419(.A(n_2372), .B(n_2315), .Z(n_2385));
	notech_nao3 i_95(.A(modrm[6]), .B(modrm[7]), .C(n_2381), .Z(n_2384));
	notech_or4 i_85(.A(n_2329), .B(n_59528), .C(n_59516), .D(n_2271), .Z(n_2382
		));
	notech_or4 i_661(.A(n_59558), .B(n_2283), .C(n_59528), .D(n_59516), .Z(n_2381
		));
	notech_and4 i_325(.A(n_4031), .B(n_4056), .C(n_4084), .D(n_2377), .Z(n_2379
		));
	notech_and2 i_339(.A(n_4066), .B(n_34038), .Z(n_2377));
	notech_or4 i_344(.A(n_2286), .B(n_34010), .C(n_2346), .D(n_34202), .Z(n_2376
		));
	notech_nor2 i_705(.A(n_2346), .B(n_59443), .Z(n_2375));
	notech_xor2 i_389(.A(n_34201), .B(modrm[3]), .Z(n_2374));
	notech_nand2 i_46(.A(n_34200), .B(modrm[4]), .Z(n_2373));
	notech_nand2 i_183(.A(n_34200), .B(n_34201), .Z(n_2372));
	notech_or4 i_693(.A(n_2279), .B(n_59598), .C(n_34193), .D(n_59603), .Z(n_2371
		));
	notech_and2 i_168(.A(n_1817), .B(n_2364), .Z(n_2365));
	notech_and2 i_756(.A(n_3991), .B(n_1813), .Z(n_2364));
	notech_and2 i_459(.A(n_2275), .B(n_2302), .Z(n_2363));
	notech_or4 i_86(.A(n_2347), .B(n_2360), .C(n_2282), .D(n_34196), .Z(n_2362
		));
	notech_nand2 i_535(.A(n_59585), .B(n_59580), .Z(n_2360));
	notech_or4 i_71(.A(n_2329), .B(n_59548), .C(n_59539), .D(n_2271), .Z(n_2359
		));
	notech_or4 i_66(.A(n_2329), .B(n_59539), .C(n_59528), .D(n_2271), .Z(n_2355
		));
	notech_and4 i_64(.A(n_223496909), .B(n_1792), .C(n_34050), .D(n_1797), .Z
		(n_2352));
	notech_or4 i_577(.A(n_2348), .B(n_2284), .C(n_34130), .D(n_34010), .Z(n_2350
		));
	notech_nor2 i_111(.A(n_2348), .B(n_2284), .Z(n_2349));
	notech_nao3 i_13(.A(n_59603), .B(n_59630), .C(n_59643), .Z(n_2348));
	notech_or2 i_600(.A(n_59643), .B(n_59612), .Z(n_2347));
	notech_or4 i_79(.A(n_2282), .B(n_2280), .C(n_59580), .D(n_59585), .Z(n_2346
		));
	notech_and4 i_351(.A(n_2141), .B(n_4013), .C(n_2058), .D(n_2343), .Z(n_2344
		));
	notech_and4 i_683(.A(n_2340), .B(n_2233), .C(n_2195), .D(n_2099), .Z(n_2343
		));
	notech_and2 i_513(.A(n_4044), .B(n_34072), .Z(n_2340));
	notech_nao3 i_671(.A(n_59639), .B(n_2272), .C(n_2338), .Z(n_2339));
	notech_nao3 i_151(.A(n_34193), .B(n_59585), .C(n_2282), .Z(n_2338));
	notech_or4 i_585(.A(n_2316), .B(n_2276), .C(n_2037), .D(n_2333), .Z(n_2337
		));
	notech_or4 i_32(.A(n_59639), .B(n_59630), .C(n_59612), .D(modrm[5]), .Z(n_2333
		));
	notech_nao3 i_574(.A(modrm[7]), .B(modrm[6]), .C(n_2290), .Z(n_2331));
	notech_or4 i_121(.A(n_59553), .B(n_2283), .C(n_59548), .D(n_59516), .Z(n_2330
		));
	notech_nao3 i_1(.A(n_59580), .B(n_59598), .C(n_59553), .Z(n_2329));
	notech_or4 i_0(.A(twobyte), .B(fpu), .C(ipg_fault), .D(n_34197), .Z(n_2328
		));
	notech_nao3 i_3(.A(n_59621), .B(n_59603), .C(n_59639), .Z(n_2325));
	notech_nor2 i_449(.A(n_59643), .B(n_59630), .Z(n_2324));
	notech_nor2 i_599(.A(opz[0]), .B(opz[2]), .Z(n_2322));
	notech_and2 i_73(.A(opz[2]), .B(n_2319), .Z(n_2321));
	notech_nor2 i_597(.A(opz[0]), .B(opz[1]), .Z(n_2319));
	notech_or4 i_92(.A(n_2403), .B(n_2311), .C(n_59580), .D(n_59598), .Z(n_2318
		));
	notech_nand2 i_584(.A(n_34193), .B(n_59585), .Z(n_2316));
	notech_nand2 i_446(.A(n_59470), .B(n_59598), .Z(n_2313));
	notech_nand3 i_41(.A(n_59639), .B(n_59603), .C(n_59630), .Z(n_2311));
	notech_and2 i_382(.A(n_59643), .B(n_59603), .Z(n_2310));
	notech_and4 i_436(.A(n_2141), .B(n_4013), .C(n_2308), .D(n_2294), .Z(n_2309
		));
	notech_and3 i_657(.A(n_4037), .B(n_1820), .C(n_1824), .Z(n_2308));
	notech_ao4 i_405(.A(n_2290), .B(n_2300), .C(n_2289), .D(n_34010), .Z(n_2303
		));
	notech_ao3 i_91(.A(n_59528), .B(n_59516), .C(n_2300), .Z(n_2301));
	notech_nao3 i_282(.A(modrm[7]), .B(modrm[6]), .C(modrm[2]), .Z(n_2300)
		);
	notech_nand3 i_68(.A(n_59511), .B(n_59548), .C(n_2271), .Z(n_2299));
	notech_nand3 i_59(.A(n_59548), .B(n_59539), .C(n_2271), .Z(n_2297));
	notech_and2 i_5(.A(n_59544), .B(n_59539), .Z(n_2296));
	notech_nao3 i_468(.A(modrm[2]), .B(n_2271), .C(n_2286), .Z(n_2295));
	notech_and2 i_790(.A(n_2258), .B(n_1821), .Z(n_2294));
	notech_nao3 i_88(.A(n_59528), .B(n_59511), .C(n_2292), .Z(n_2293));
	notech_nand3 i_276(.A(modrm[7]), .B(modrm[2]), .C(modrm[6]), .Z(n_2292)
		);
	notech_and2 i_393(.A(n_2278), .B(n_34053), .Z(n_2291));
	notech_nand2 i_2(.A(n_59527), .B(n_59511), .Z(n_2290));
	notech_nand2 i_6(.A(n_59511), .B(n_59544), .Z(n_2289));
	notech_or4 i_590(.A(modrm[2]), .B(n_59544), .C(n_59511), .D(n_34010), .Z
		(n_2288));
	notech_and4 i_120(.A(modrm[7]), .B(n_59522), .C(n_59539), .D(modrm[6]), 
		.Z(n_2287));
	notech_nand2 i_777939(.A(n_59522), .B(n_59539), .Z(n_2286));
	notech_or4 i_75(.A(n_59425), .B(n_2280), .C(n_59470), .D(n_59585), .Z(n_2285
		));
	notech_nao3 i_856(.A(n_59576), .B(n_59598), .C(n_59425), .Z(n_2284));
	notech_nand2 i_589(.A(n_59576), .B(n_59598), .Z(n_2283));
	notech_or4 i_9(.A(fpu), .B(ipg_fault), .C(n_34197), .D(n_34205), .Z(n_2282
		));
	notech_nao3 i_44(.A(n_59630), .B(n_59612), .C(n_59643), .Z(n_2280));
	notech_or2 i_593(.A(n_59643), .B(n_59621), .Z(n_2279));
	notech_or4 i_857(.A(fpu), .B(ipg_fault), .C(op[7]), .D(n_34205), .Z(n_2276
		));
	notech_and2 i_537(.A(n_59621), .B(n_59603), .Z(n_2272));
	notech_and2 i_230(.A(modrm[7]), .B(modrm[6]), .Z(n_2271));
	notech_and4 i_281(.A(n_3591), .B(n_3560), .C(n_717), .D(n_1593), .Z(n_2270
		));
	notech_or2 i_2397(.A(n_2398), .B(n_59522), .Z(n_2269));
	notech_nand3 i_308(.A(n_2757), .B(n_3548), .C(n_1951), .Z(\udeco[8] ));
	notech_nand2 i_2345(.A(modrm[3]), .B(n_3174), .Z(n_2267));
	notech_nao3 i_2349(.A(opz[1]), .B(n_2322), .C(n_2247), .Z(n_2266));
	notech_or4 i_2341(.A(n_2410), .B(n_2373), .C(n_3954), .D(n_59443), .Z(n_2265
		));
	notech_or2 i_335(.A(n_2485), .B(n_2333), .Z(n_2264));
	notech_or4 i_2350(.A(n_59558), .B(n_2248), .C(n_59576), .D(n_59598), .Z(n_2263
		));
	notech_nand2 i_2353(.A(n_59533), .B(n_2251), .Z(n_2262));
	notech_or4 i_144(.A(n_2286), .B(modrm[2]), .C(n_2285), .D(n_59452), .Z(n_2258
		));
	notech_or4 i_2344(.A(n_2412), .B(n_59522), .C(n_59511), .D(n_2271), .Z(n_2257
		));
	notech_or4 i_2342(.A(n_59558), .B(n_2316), .C(n_2389), .D(n_2278), .Z(n_2256
		));
	notech_or4 i_23111154(.A(n_2313), .B(n_59522), .C(n_2271), .D(n_34150), 
		.Z(n_2255));
	notech_or4 i_2351(.A(n_59558), .B(n_59594), .C(n_59470), .D(n_2249), .Z(n_2254
		));
	notech_or4 i_2346(.A(n_2347), .B(n_2338), .C(n_2512), .D(n_59621), .Z(n_2253
		));
	notech_or4 i_822(.A(n_2280), .B(n_59558), .C(n_59533), .D(n_59576), .Z(n_2252
		));
	notech_nand2 i_202(.A(n_2433), .B(n_2678), .Z(n_2251));
	notech_and3 i_203(.A(n_2141), .B(n_4013), .C(n_2140), .Z(n_2250));
	notech_and2 i_205(.A(n_2448), .B(n_2243), .Z(n_2249));
	notech_ao4 i_209(.A(n_2486), .B(n_2288), .C(n_2348), .D(n_2289), .Z(n_2248
		));
	notech_ao4 i_219(.A(n_2318), .B(n_2297), .C(n_2401), .D(n_2101), .Z(n_2247
		));
	notech_ao3 i_222(.A(n_2275), .B(n_2302), .C(n_2301), .Z(n_2245));
	notech_and2 i_404(.A(n_59493), .B(n_34130), .Z(n_2244));
	notech_nao3 i_2339(.A(n_2310), .B(n_59630), .C(n_2244), .Z(n_2243));
	notech_and4 i_320(.A(n_2484), .B(n_2703), .C(n_3500), .D(n_3465), .Z(n_2241
		));
	notech_nand2 i_2293(.A(n_3174), .B(modrm[4]), .Z(n_2240));
	notech_or4 i_2294(.A(n_2410), .B(n_2373), .C(n_2230), .D(n_59443), .Z(n_2239
		));
	notech_or4 i_287(.A(n_2383), .B(n_2486), .C(n_2290), .D(n_2300), .Z(n_2238
		));
	notech_nand2 i_2291(.A(n_59612), .B(n_34117), .Z(n_2237));
	notech_or4 i_23111283(.A(n_2348), .B(n_2320), .C(n_2275), .D(n_2284), .Z
		(n_223496909));
	notech_or4 i_23111397(.A(n_59452), .B(n_2337), .C(n_59544), .D(n_59533),
		 .Z(n_2233));
	notech_or4 i_2290(.A(n_2285), .B(n_59522), .C(n_59511), .D(n_2271), .Z(n_2232
		));
	notech_or4 i_23111349(.A(n_2347), .B(n_2290), .C(n_2408), .D(n_59621), .Z
		(n_2231));
	notech_and2 i_200(.A(n_2382), .B(n_2485), .Z(n_2230));
	notech_or4 i_2286(.A(n_59493), .B(n_2329), .C(n_2325), .D(n_59461), .Z(n_2229
		));
	notech_or4 i_2285(.A(n_2285), .B(n_59533), .C(n_59522), .D(n_59452), .Z(n_2228
		));
	notech_and4 i_334(.A(n_2694), .B(n_3458), .C(n_3429), .D(n_2704), .Z(n_2227
		));
	notech_nand2 i_2248(.A(n_3174), .B(modrm[5]), .Z(n_2226));
	notech_nao3 i_2249(.A(n_34009), .B(n_34141), .C(n_2499), .Z(n_2223));
	notech_or2 i_2243(.A(n_2065), .B(n_59470), .Z(n_2222));
	notech_or4 i_2247(.A(n_2360), .B(n_59553), .C(n_59434), .D(n_2297), .Z(n_2221
		));
	notech_or4 i_2250(.A(n_2316), .B(n_2276), .C(n_2289), .D(n_2280), .Z(n_2220
		));
	notech_and4 i_345(.A(n_2904), .B(n_2703), .C(n_2484), .D(n_3425), .Z(n_221996908
		));
	notech_or4 i_149(.A(n_2244), .B(n_2185), .C(n_59603), .D(n_2386), .Z(n_2218
		));
	notech_or2 i_2216(.A(n_2065), .B(n_59511), .Z(n_2217));
	notech_or4 i_23110611(.A(n_2329), .B(n_59533), .C(n_59522), .D(n_2389), 
		.Z(n_2216));
	notech_and4 i_431(.A(n_2689), .B(n_2501), .C(n_2499), .D(n_2422), .Z(n_2215
		));
	notech_or2 i_2215(.A(n_2215), .B(n_2359), .Z(n_2213));
	notech_and4 i_363(.A(n_2484), .B(n_3397), .C(n_2904), .D(n_2704), .Z(n_2208
		));
	notech_or2 i_2183(.A(n_2215), .B(n_2497), .Z(n_2207));
	notech_or4 i_23111151(.A(n_2316), .B(n_59522), .C(n_34150), .D(n_59461),
		 .Z(n_2206));
	notech_and2 i_353(.A(n_2295), .B(n_2293), .Z(n_2205));
	notech_or4 i_361(.A(n_59493), .B(n_2292), .C(n_2329), .D(n_34138), .Z(n_2202
		));
	notech_nand3 i_385(.A(n_3364), .B(n_3343), .C(n_1951), .Z(\udeco[16] )
		);
	notech_nao3 i_2126(.A(opz[1]), .B(n_2322), .C(n_2187), .Z(n_2200));
	notech_or2 i_2123(.A(n_2883), .B(n_34200), .Z(n_2199));
	notech_or2 i_297(.A(n_4090), .B(n_34138), .Z(n_2198));
	notech_or4 i_2125(.A(n_2373), .B(n_59443), .C(n_2410), .D(n_2115), .Z(n_2197
		));
	notech_or4 i_2120(.A(n_59416), .B(n_2037), .C(n_3954), .D(n_59443), .Z(n_2196
		));
	notech_or4 i_153(.A(n_59643), .B(n_2330), .C(n_59634), .D(n_59612), .Z(n_2195
		));
	notech_or4 i_2119(.A(n_2292), .B(n_2285), .C(n_59544), .D(n_59533), .Z(n_2193
		));
	notech_or4 i_677(.A(n_34089), .B(n_59533), .C(n_59522), .D(n_34136), .Z(n_2192
		));
	notech_or2 i_2982(.A(n_2300), .B(n_34128), .Z(n_2190));
	notech_or4 i_1241(.A(n_59522), .B(n_34150), .C(n_59576), .D(n_59452), .Z
		(n_2189));
	notech_or4 i_179(.A(n_59643), .B(n_2403), .C(n_2360), .D(n_59544), .Z(n_2188
		));
	notech_ao4 i_181(.A(n_4065), .B(n_2297), .C(n_2098), .D(n_2101), .Z(n_2187
		));
	notech_and2 i_524(.A(n_2668), .B(n_3154), .Z(n_2186));
	notech_and3 i_394(.A(n_2383), .B(n_34136), .C(n_34080), .Z(n_2185));
	notech_or4 i_2116(.A(n_2285), .B(n_59544), .C(n_59533), .D(n_59461), .Z(n_2183
		));
	notech_nao3 i_2115(.A(opz[1]), .B(n_2322), .C(n_2350), .Z(n_2181));
	notech_nand3 i_2110(.A(n_3895), .B(n_59634), .C(n_2310), .Z(n_2180));
	notech_or4 i_39(.A(n_2458), .B(n_59527), .C(n_59511), .D(n_59461), .Z(n_2179
		));
	notech_and4 i_400(.A(n_3309), .B(n_3302), .C(n_3273), .D(n_2562), .Z(n_2177
		));
	notech_or2 i_2061(.A(n_2883), .B(n_34201), .Z(n_2175));
	notech_or4 i_2060(.A(n_59416), .B(n_2373), .C(n_3836), .D(n_59443), .Z(n_2174
		));
	notech_nand2 i_2064(.A(n_59612), .B(n_34163), .Z(n_2173));
	notech_nao3 i_2062(.A(n_2321), .B(n_34144), .C(n_2101), .Z(n_2172));
	notech_or4 i_2063(.A(n_2403), .B(n_2161), .C(n_2313), .D(n_2311), .Z(n_2170
		));
	notech_or4 i_2058(.A(n_59416), .B(n_2037), .C(n_59443), .D(n_2355), .Z(n_2169
		));
	notech_nao3 i_2056(.A(n_2385), .B(n_34007), .C(n_2214), .Z(n_2168));
	notech_or4 i_227(.A(n_59434), .B(n_59461), .C(n_34130), .D(n_34136), .Z(n_2166
		));
	notech_or4 i_2059(.A(n_59544), .B(n_59533), .C(n_59461), .D(n_34054), .Z
		(n_2163));
	notech_ao4 i_518(.A(n_2297), .B(n_34158), .C(n_2275), .D(n_2149), .Z(n_2161
		));
	notech_or4 i_224(.A(n_59493), .B(n_2486), .C(n_59461), .D(n_34080), .Z(n_2159
		));
	notech_or4 i_2050(.A(n_59553), .B(n_2594), .C(n_59576), .D(n_59594), .Z(n_2155
		));
	notech_and2 i_290(.A(n_2285), .B(n_34054), .Z(n_2154));
	notech_and2 i_328(.A(n_2320), .B(n_34158), .Z(n_2149));
	notech_and4 i_414(.A(n_2757), .B(n_3257), .C(n_1504), .D(n_520), .Z(n_2146
		));
	notech_or2 i_2004(.A(n_2883), .B(n_59443), .Z(n_2145));
	notech_or4 i_2002(.A(n_59416), .B(n_2037), .C(n_3836), .D(n_59443), .Z(n_2144
		));
	notech_nand2 i_2005(.A(n_59634), .B(n_34163), .Z(n_2143));
	notech_and3 i_2003(.A(n_2287), .B(n_2375), .C(n_2385), .Z(n_2142));
	notech_nao3 i_1250(.A(n_2397), .B(n_59461), .C(n_2276), .Z(n_2141));
	notech_or4 i_180(.A(n_59643), .B(n_2403), .C(n_2283), .D(n_59630), .Z(n_2140
		));
	notech_and3 i_326(.A(n_2485), .B(n_2401), .C(n_2497), .Z(n_2139));
	notech_or4 i_675(.A(n_59502), .B(n_59553), .C(n_59434), .D(n_2027), .Z(n_2137
		));
	notech_or2 i_591(.A(n_2497), .B(n_34138), .Z(n_2136));
	notech_and4 i_438(.A(n_530), .B(n_2703), .C(n_3213), .D(n_537), .Z(n_2135
		));
	notech_or4 i_1968(.A(n_59416), .B(n_2373), .C(n_3954), .D(modrm[5]), .Z(n_2134
		));
	notech_or4 i_1967(.A(n_59544), .B(n_59533), .C(n_59461), .D(n_34151), .Z
		(n_2132));
	notech_nao3 i_1935(.A(n_34200), .B(n_34201), .C(n_2376), .Z(n_2131));
	notech_or4 i_1934(.A(n_59416), .B(n_2373), .C(n_2384), .D(n_59443), .Z(n_2130
		));
	notech_or4 i_1933(.A(n_59502), .B(n_59553), .C(n_59434), .D(n_2302), .Z(n_2129
		));
	notech_ao3 i_1931(.A(n_2299), .B(n_2297), .C(n_2301), .Z(n_2128));
	notech_and4 i_48310302(.A(n_719), .B(n_3171), .C(n_3143), .D(n_1950), .Z
		(n_2127));
	notech_nand3 i_1902(.A(opz[1]), .B(n_2322), .C(n_2117), .Z(n_2126));
	notech_or2 i_1898(.A(n_3728), .B(n_34200), .Z(n_2125));
	notech_or4 i_1901(.A(n_59416), .B(n_2037), .C(n_2115), .D(n_59443), .Z(n_2122
		));
	notech_or2 i_1899(.A(n_3697), .B(n_59511), .Z(n_2121));
	notech_or2 i_1897(.A(n_2151), .B(n_59527), .Z(n_2120));
	notech_or2 i_1900(.A(n_2052), .B(n_34053), .Z(n_2119));
	notech_nand2 i_169(.A(n_2988), .B(n_2350), .Z(n_2117));
	notech_and3 i_174(.A(n_2497), .B(n_2359), .C(n_2355), .Z(n_2115));
	notech_nand3 i_124(.A(n_59452), .B(n_59594), .C(n_2536), .Z(n_2111));
	notech_nao3 i_472(.A(n_1718), .B(n_3141), .C(n_4024), .Z(\udeco[25] ));
	notech_nand2 i_1860(.A(modrm[4]), .B(n_34066), .Z(n_2109));
	notech_or4 i_838(.A(n_59643), .B(n_59630), .C(n_59612), .D(n_2098), .Z(n_2108
		));
	notech_nand2 i_1861(.A(n_59612), .B(n_34067), .Z(n_2107));
	notech_nao3 i_1197(.A(opz[2]), .B(n_2319), .C(n_2350), .Z(n_2106));
	notech_or2 i_1858(.A(n_2151), .B(n_59585), .Z(n_2105));
	notech_nao3 i_827(.A(n_2287), .B(n_2375), .C(n_2374), .Z(n_2104));
	notech_or4 i_47(.A(n_2596), .B(n_59544), .C(n_59511), .D(n_59461), .Z(n_2103
		));
	notech_ao3 i_16377884(.A(opz[2]), .B(n_2319), .C(n_2083), .Z(n_2102));
	notech_and2 i_633(.A(n_2499), .B(n_2422), .Z(n_2101));
	notech_ao3 i_1824(.A(n_34009), .B(n_34013), .C(n_2499), .Z(n_2100));
	notech_and2 i_329(.A(n_2401), .B(n_2355), .Z(n_2098));
	notech_or4 i_1823(.A(n_59416), .B(n_2315), .C(n_3836), .D(n_59443), .Z(n_2097
		));
	notech_and4 i_1811(.A(n_2278), .B(n_2275), .C(n_34053), .D(n_2293), .Z(n_2095
		));
	notech_and4 i_546(.A(n_3091), .B(n_2903), .C(n_34189), .D(n_34149), .Z(n_2092
		));
	notech_or2 i_416(.A(n_3957), .B(n_2098), .Z(n_2091));
	notech_nao3 i_1775(.A(opz[1]), .B(n_2322), .C(n_2083), .Z(n_2090));
	notech_or4 i_1776(.A(n_2348), .B(n_59502), .C(n_59425), .D(n_2291), .Z(n_2089
		));
	notech_or4 i_1778(.A(n_2311), .B(n_3963), .C(n_59544), .D(n_59533), .Z(n_2087
		));
	notech_or4 i_1777(.A(n_59502), .B(n_2280), .C(n_59425), .D(n_34152), .Z(n_2086
		));
	notech_ao4 i_516(.A(n_2101), .B(n_2355), .C(n_4065), .D(n_2027), .Z(n_2083
		));
	notech_nand3 i_745(.A(n_3054), .B(n_2079), .C(n_34207), .Z(\udeco[108] )
		);
	notech_nand2 i_1646(.A(opz[0]), .B(n_2067), .Z(n_2079));
	notech_nor2 i_192(.A(n_2400), .B(n_3845), .Z(n_2078));
	notech_ao4 i_1647(.A(n_2418), .B(n_34154), .C(n_2301), .D(n_3908), .Z(n_2077
		));
	notech_or2 i_1648(.A(n_2359), .B(n_2069), .Z(n_2075));
	notech_or2 i_1645(.A(n_2523), .B(n_3961), .Z(n_2074));
	notech_or4 i_55(.A(modrm[2]), .B(n_2330), .C(n_59452), .D(n_34138), .Z(n_2073
		));
	notech_or4 i_1649(.A(n_2347), .B(n_59493), .C(n_3963), .D(n_59621), .Z(n_2072
		));
	notech_or4 i_23110701(.A(n_34089), .B(n_2329), .C(n_2331), .D(modrm[5]),
		 .Z(n_2071));
	notech_or4 i_23110704(.A(n_2586), .B(n_59548), .C(n_59533), .D(n_59452),
		 .Z(n_2070));
	notech_and3 i_163(.A(n_2400), .B(n_34089), .C(n_34138), .Z(n_2069));
	notech_nand3 i_165(.A(n_3018), .B(n_3013), .C(n_2955), .Z(n_2067));
	notech_or4 i_1629(.A(n_59553), .B(n_2574), .C(n_59576), .D(n_59585), .Z(n_2063
		));
	notech_nand2 i_1627(.A(n_2407), .B(n_2061), .Z(n_2062));
	notech_or4 i_254(.A(n_59643), .B(n_59493), .C(n_59612), .D(n_59621), .Z(n_2061
		));
	notech_and2 i_294(.A(n_2383), .B(n_2329), .Z(n_2059));
	notech_nao3 i_1622(.A(n_34011), .B(n_34206), .C(n_2407), .Z(n_2057));
	notech_or4 i_1620(.A(n_59553), .B(n_2407), .C(n_59576), .D(n_59594), .Z(n_2056
		));
	notech_and4 i_762(.A(n_3005), .B(n_2987), .C(n_2054), .D(n_34207), .Z(n_2055
		));
	notech_nand2 i_1590(.A(opz[1]), .B(n_34168), .Z(n_2054));
	notech_nao3 i_1586(.A(opz[1]), .B(n_2322), .C(n_2988), .Z(n_2053));
	notech_or2 i_1584(.A(adz), .B(n_2036), .Z(n_2051));
	notech_nao3 i_1585(.A(n_34198), .B(n_2037), .C(n_2488), .Z(n_2050));
	notech_or4 i_1228(.A(n_2485), .B(n_2490), .C(n_2492), .D(modrm[0]), .Z(n_2046
		));
	notech_or4 i_854(.A(n_59502), .B(n_59553), .C(n_59434), .D(n_2413), .Z(n_2045
		));
	notech_or4 i_1589(.A(n_59553), .B(n_2313), .C(n_2486), .D(n_2288), .Z(n_2042
		));
	notech_or4 i_1592(.A(n_59434), .B(n_3963), .C(n_59443), .D(n_2295), .Z(n_2041
		));
	notech_or4 i_1587(.A(n_59558), .B(n_2428), .C(n_59470), .D(n_59585), .Z(n_2040
		));
	notech_and4 i_158(.A(n_2309), .B(n_2958), .C(n_2975), .D(n_2955), .Z(n_2038
		));
	notech_nand2 i_564(.A(modrm[3]), .B(modrm[4]), .Z(n_2037));
	notech_and3 i_197(.A(n_2327), .B(n_4047), .C(n_3981), .Z(n_2036));
	notech_nand3 i_1566(.A(n_59643), .B(n_2272), .C(n_34013), .Z(n_2034));
	notech_or2 i_1567(.A(n_2523), .B(n_2512), .Z(n_2033));
	notech_or4 i_826(.A(n_2279), .B(n_59558), .C(n_59603), .D(n_59511), .Z(n_2032
		));
	notech_or4 i_1562(.A(n_2347), .B(n_2512), .C(n_59621), .D(n_2059), .Z(n_2031
		));
	notech_or4 i_1282(.A(n_2348), .B(n_59425), .C(n_1888), .D(n_59502), .Z(n_2030
		));
	notech_or4 i_1553(.A(n_3963), .B(n_2027), .C(n_59612), .D(n_34157), .Z(n_2028
		));
	notech_and2 i_301(.A(n_2275), .B(n_2297), .Z(n_2027));
	notech_or4 i_845(.A(n_2313), .B(n_59425), .C(n_2348), .D(n_2387), .Z(n_2026
		));
	notech_or4 i_1543(.A(n_2214), .B(n_2497), .C(modrm[3]), .D(n_34201), .Z(n_2025
		));
	notech_or4 i_1541(.A(n_2280), .B(n_59558), .C(n_59538), .D(n_59470), .Z(n_2021
		));
	notech_and4 i_796(.A(n_2939), .B(n_2936), .C(n_1718), .D(n_2890), .Z(n_2020
		));
	notech_or2 i_1174(.A(n_2400), .B(n_2401), .Z(n_2019));
	notech_or4 i_834(.A(n_59493), .B(n_59603), .C(n_34157), .D(n_34080), .Z(n_2014
		));
	notech_ao4 i_178(.A(n_2542), .B(n_2541), .C(n_2369), .D(n_2354), .Z(n_2013
		));
	notech_nand3 i_873(.A(n_2881), .B(n_1593), .C(n_2011), .Z(\udeco[117] )
		);
	notech_nand2 i_1366(.A(n_34119), .B(n_34170), .Z(n_2011));
	notech_nand2 i_1367(.A(modrm[4]), .B(n_3773), .Z(n_2010));
	notech_nand2 i_1368(.A(modrm[1]), .B(n_2007), .Z(n_2009));
	notech_or4 i_1365(.A(n_59425), .B(n_34089), .C(n_59516), .D(n_59585), .Z
		(n_2008));
	notech_nand3 i_140(.A(n_2099), .B(n_3736), .C(n_2654), .Z(n_2007));
	notech_mux2 i_396(.S(n_59594), .A(n_34201), .B(n_34199), .Z(n_2006));
	notech_or4 i_1361(.A(n_59502), .B(n_59558), .C(n_2519), .D(n_34206), .Z(n_2005
		));
	notech_or4 i_90810224(.A(n_2002), .B(n_2001), .C(n_2820), .D(n_1180), .Z
		(\udeco[120] ));
	notech_and2 i_1287(.A(n_3763), .B(n_1968), .Z(n_2002));
	notech_and2 i_1281(.A(n_34056), .B(n_34055), .Z(n_2001));
	notech_and2 i_1285(.A(modrm[0]), .B(n_34171), .Z(n_2000));
	notech_and2 i_1286(.A(modrm[3]), .B(n_1988), .Z(n_1998));
	notech_nor2 i_1288(.A(n_2362), .B(n_1989), .Z(n_1997));
	notech_or4 i_1141(.A(n_59502), .B(n_2280), .C(n_59425), .D(n_2413), .Z(n_1995
		));
	notech_or4 i_1280(.A(n_59563), .B(n_2517), .C(n_59580), .D(n_59594), .Z(n_1994
		));
	notech_or4 i_1284(.A(n_2347), .B(n_2338), .C(n_2244), .D(n_59621), .Z(n_1990
		));
	notech_and4 i_116(.A(n_2275), .B(n_2297), .C(n_2278), .D(n_2299), .Z(n_1989
		));
	notech_nand3 i_118(.A(n_2480), .B(n_1777), .C(n_2415), .Z(n_1988));
	notech_and4 i_655(.A(n_2309), .B(n_2760), .C(n_2717), .D(n_2759), .Z(n_1986
		));
	notech_or4 i_1275(.A(n_2315), .B(n_2214), .C(n_2330), .D(n_59452), .Z(n_1985
		));
	notech_or2 i_1273(.A(n_2382), .B(n_34138), .Z(n_1982));
	notech_or4 i_1272(.A(n_2372), .B(n_2214), .C(n_2330), .D(n_59452), .Z(n_1981
		));
	notech_or4 i_908(.A(n_1979), .B(n_1321), .C(n_1977), .D(n_2785), .Z(\udeco[121] 
		));
	notech_and2 i_1239(.A(n_1968), .B(n_34172), .Z(n_1979));
	notech_and2 i_1231(.A(n_34055), .B(n_34170), .Z(n_1977));
	notech_and2 i_1237(.A(modrm[1]), .B(n_34171), .Z(n_1976));
	notech_and2 i_1238(.A(modrm[4]), .B(n_1964), .Z(n_1975));
	notech_nand3 i_114(.A(n_2688), .B(n_2757), .C(n_2166), .Z(n_1968));
	notech_mux2 i_422(.S(n_59594), .A(n_34199), .B(n_34201), .Z(n_1965));
	notech_nand3 i_115(.A(n_2395), .B(n_1777), .C(n_2415), .Z(n_1964));
	notech_or4 i_483(.A(n_1326), .B(n_222998902), .C(n_1956), .D(n_34111), .Z
		(\udeco[122] ));
	notech_and2 i_1192(.A(modrm[2]), .B(n_1946), .Z(n_1956));
	notech_nand2 i_1191(.A(modrm[5]), .B(n_1945), .Z(n_1955));
	notech_nand2 i_1189(.A(n_1944), .B(n_34146), .Z(n_1954));
	notech_or4 i_1190(.A(n_2387), .B(n_59612), .C(n_34157), .D(n_34080), .Z(n_1952
		));
	notech_or4 i_1187(.A(n_59563), .B(n_59434), .C(n_59580), .D(n_3761), .Z(n_1949
		));
	notech_or2 i_1186(.A(n_2734), .B(n_59470), .Z(n_1947));
	notech_nand3 i_104(.A(n_2719), .B(n_2717), .C(n_2091), .Z(n_1946));
	notech_nand3 i_112(.A(n_2723), .B(n_4017), .C(n_2726), .Z(n_1945));
	notech_mux2 i_506(.S(n_59594), .A(n_59479), .B(modrm[2]), .Z(n_1944));
	notech_mux2 i_505(.S(n_59594), .A(modrm[2]), .B(n_59479), .Z(n_1943));
	notech_or2 i_1180(.A(n_1940), .B(n_2285), .Z(n_1941));
	notech_and4 i_113(.A(n_2027), .B(n_2387), .C(n_2302), .D(n_34053), .Z(n_1940
		));
	notech_or4 i_23111403(.A(n_59452), .B(n_2052), .C(n_59544), .D(n_59538),
		 .Z(n_1938));
	notech_and2 i_313(.A(n_2422), .B(n_2325), .Z(n_1937));
	notech_or4 i_1170(.A(n_2393), .B(n_59538), .C(n_59527), .D(n_34010), .Z(n_1936
		));
	notech_and4 i_1157(.A(n_59612), .B(n_2324), .C(n_2296), .D(n_34011), .Z(n_1933
		));
	notech_or2 i_1156(.A(n_2101), .B(n_2382), .Z(n_1932));
	notech_or2 i_1123(.A(n_3845), .B(n_34138), .Z(n_1930));
	notech_or4 i_1116(.A(n_59502), .B(n_59558), .C(n_34089), .D(n_2289), .Z(n_1921
		));
	notech_or4 i_1057(.A(n_2214), .B(n_2382), .C(n_34200), .D(n_34201), .Z(n_1919
		));
	notech_or4 i_1044(.A(n_2348), .B(n_34130), .C(adz), .D(n_2059), .Z(n_1918
		));
	notech_or4 i_284(.A(n_59558), .B(n_2286), .C(n_59594), .D(n_59470), .Z(n_1917
		));
	notech_and2 i_1042(.A(n_2330), .B(n_1917), .Z(n_1916));
	notech_or2 i_1030(.A(n_3836), .B(n_34138), .Z(n_1915));
	notech_or2 i_1028(.A(n_2494), .B(n_1913), .Z(n_1914));
	notech_and3 i_311(.A(n_2373), .B(n_2372), .C(n_2037), .Z(n_1913));
	notech_nao3 i_1027(.A(n_34198), .B(n_2385), .C(n_2488), .Z(n_1912));
	notech_or2 i_1018(.A(n_2497), .B(n_2486), .Z(n_1911));
	notech_or4 i_1011(.A(n_59594), .B(n_59470), .C(n_59527), .D(n_34150), .Z
		(n_1907));
	notech_ao4 i_1003(.A(n_2037), .B(n_2486), .C(n_59603), .D(n_2279), .Z(n_1902
		));
	notech_or4 i_992(.A(n_2330), .B(modrm[6]), .C(modrm[7]), .D(n_2505), .Z(n_1901
		));
	notech_and2 i_989(.A(modrm[6]), .B(modrm[7]), .Z(n_1900));
	notech_or4 i_975(.A(n_2412), .B(n_59538), .C(n_59527), .D(n_59461), .Z(n_1896
		));
	notech_or4 i_968(.A(n_2458), .B(n_59538), .C(n_59527), .D(n_59461), .Z(n_1895
		));
	notech_or4 i_956(.A(n_2313), .B(n_59425), .C(n_2280), .D(n_2387), .Z(n_1892
		));
	notech_or2 i_946(.A(n_3935), .B(n_3963), .Z(n_1890));
	notech_and4 i_940(.A(n_2027), .B(n_2387), .C(n_34053), .D(n_2413), .Z(n_1888
		));
	notech_or4 i_938(.A(modrm[1]), .B(n_2553), .C(n_34198), .D(n_2495), .Z(n_1887
		));
	notech_or4 i_937(.A(modrm[1]), .B(n_2553), .C(modrm[0]), .D(n_2492), .Z(n_1886
		));
	notech_mux2 i_321(.S(modrm[0]), .A(n_1882), .B(n_2037), .Z(n_1885));
	notech_nand3 i_322(.A(n_2372), .B(n_2315), .C(n_2037), .Z(n_1882));
	notech_nand2 i_932(.A(n_2037), .B(modrm[0]), .Z(n_1879));
	notech_or4 i_922(.A(n_2300), .B(n_2455), .C(n_59544), .D(n_59538), .Z(n_1877
		));
	notech_or4 i_913(.A(n_2360), .B(n_59558), .C(n_34089), .D(n_59493), .Z(n_1875
		));
	notech_or4 i_898(.A(modrm[1]), .B(n_2553), .C(modrm[0]), .D(n_2372), .Z(n_1874
		));
	notech_or4 i_897(.A(modrm[1]), .B(n_2553), .C(n_2315), .D(n_34198), .Z(n_1873
		));
	notech_mux2 i_312(.S(modrm[0]), .A(n_2373), .B(n_2037), .Z(n_1872));
	notech_or4 i_894(.A(n_2497), .B(n_2333), .C(n_1872), .D(n_34199), .Z(n_1871
		));
	notech_or4 i_893(.A(n_2485), .B(n_2372), .C(n_2490), .D(modrm[0]), .Z(n_1869
		));
	notech_ao4 i_881(.A(n_2333), .B(n_2288), .C(n_2486), .D(n_2295), .Z(n_1858
		));
	notech_or4 i_875(.A(n_2383), .B(n_2333), .C(n_2290), .D(n_2300), .Z(n_1857
		));
	notech_nao3 i_870(.A(n_59585), .B(n_2530), .C(n_2300), .Z(n_1855));
	notech_nao3 i_869(.A(n_59594), .B(n_2536), .C(n_2292), .Z(n_1854));
	notech_or4 i_825(.A(n_59434), .B(n_2302), .C(n_3963), .D(n_59479), .Z(n_1851
		));
	notech_or4 i_954(.A(n_2475), .B(n_2445), .C(n_1849), .D(n_1838), .Z(\udeco[126] 
		));
	notech_and2 i_752(.A(modrm[2]), .B(n_34177), .Z(n_1849));
	notech_nand2 i_741(.A(n_1943), .B(n_34146), .Z(n_1848));
	notech_and4 i_743(.A(n_59452), .B(n_1944), .C(n_2296), .D(n_2427), .Z(n_1846
		));
	notech_or2 i_740(.A(n_2433), .B(n_59538), .Z(n_1843));
	notech_and2 i_69(.A(n_2032), .B(n_3733), .Z(n_1842));
	notech_and4 i_81(.A(n_1837), .B(n_2417), .C(n_2415), .D(n_2406), .Z(n_1841
		));
	notech_and4 i_82(.A(n_2352), .B(n_2344), .C(n_1905), .D(n_1825), .Z(n_1840
		));
	notech_and2 i_749(.A(n_59479), .B(n_34178), .Z(n_1838));
	notech_or4 i_735(.A(n_59558), .B(n_2316), .C(n_34089), .D(n_2387), .Z(n_1837
		));
	notech_nand3 i_734(.A(n_59643), .B(n_2272), .C(n_34141), .Z(n_1835));
	notech_or4 i_731(.A(n_2276), .B(n_2407), .C(n_59580), .D(n_59594), .Z(n_1833
		));
	notech_or4 i_673(.A(n_2299), .B(n_3963), .C(n_59612), .D(n_34157), .Z(n_1831
		));
	notech_or4 i_718(.A(n_2393), .B(n_59527), .C(n_59511), .D(n_59452), .Z(n_1829
		));
	notech_or4 i_717(.A(n_2313), .B(n_59425), .C(n_2280), .D(n_2299), .Z(n_1828
		));
	notech_nao3 i_851(.A(n_59643), .B(n_2272), .C(n_4072), .Z(n_1825));
	notech_or2 i_656(.A(n_2303), .B(n_2285), .Z(n_1824));
	notech_and3 i_340(.A(n_2278), .B(n_2293), .C(n_34053), .Z(n_1822));
	notech_or2 i_652(.A(n_2285), .B(n_1822), .Z(n_1821));
	notech_or2 i_651(.A(n_2285), .B(n_2027), .Z(n_1820));
	notech_and2 i_647(.A(n_2295), .B(n_2302), .Z(n_1819));
	notech_and2 i_286(.A(n_2297), .B(n_34152), .Z(n_1818));
	notech_or4 i_621(.A(n_2348), .B(n_59502), .C(n_59425), .D(n_1818), .Z(n_1817
		));
	notech_or4 i_620(.A(n_2348), .B(n_59502), .C(n_59425), .D(n_2299), .Z(n_1813
		));
	notech_and4 i_615(.A(n_2278), .B(n_2275), .C(n_2302), .D(n_34053), .Z(n_1812
		));
	notech_ao3 i_531(.A(n_59612), .B(n_2324), .C(n_2330), .Z(n_1807));
	notech_or4 i_529(.A(n_59416), .B(n_2185), .C(n_59527), .D(n_59511), .Z(n_1806
		));
	notech_or4 i_502(.A(n_59558), .B(n_59434), .C(n_2297), .D(n_59580), .Z(n_1805
		));
	notech_and2 i_463(.A(n_2289), .B(n_2290), .Z(n_1802));
	notech_or2 i_23111394(.A(n_2337), .B(n_34053), .Z(n_1801));
	notech_or4 i_184(.A(n_2488), .B(n_34200), .C(n_34201), .D(n_34198), .Z(n_1800
		));
	notech_nand3 i_145(.A(n_59452), .B(n_2530), .C(n_59594), .Z(n_1798));
	notech_or4 i_839(.A(n_2313), .B(n_59425), .C(n_2280), .D(n_2290), .Z(n_1797
		));
	notech_or4 i_855(.A(n_2292), .B(n_2455), .C(n_59544), .D(n_59538), .Z(n_1796
		));
	notech_ao3 i_1104(.A(n_34141), .B(n_2321), .C(n_2101), .Z(n_1795));
	notech_or4 i_1225(.A(adz), .B(n_59621), .C(n_2347), .D(n_1916), .Z(n_1794
		));
	notech_or4 i_1291(.A(n_59558), .B(n_2448), .C(n_59576), .D(n_59594), .Z(n_1793
		));
	notech_or4 i_1233(.A(n_2347), .B(n_2284), .C(n_2018), .D(n_59621), .Z(n_1792
		));
	notech_nand3 i_520(.A(n_2278), .B(n_2299), .C(n_3761), .Z(n_1791));
	notech_and4 i_78577136(.A(n_1778), .B(n_3280), .C(n_3109), .D(n_1785), .Z
		(n_1789));
	notech_and4 i_78177140(.A(n_1950), .B(n_1638), .C(n_738), .D(n_3994), .Z
		(n_1785));
	notech_and4 i_78077141(.A(n_811), .B(n_3098), .C(n_2579), .D(n_3079), .Z
		(n_1778));
	notech_and4 i_11577865(.A(n_2571), .B(n_4013), .C(n_2394), .D(n_2365), .Z
		(n_1770));
	notech_and4 i_67377222(.A(n_1741), .B(n_1738), .C(n_176196907), .D(n_34079
		), .Z(n_1762));
	notech_and4 i_67077223(.A(n_1745), .B(n_1744), .C(n_1759), .D(n_1702), .Z
		(n_176196907));
	notech_and4 i_66877225(.A(n_3993), .B(n_1757), .C(n_2305), .D(n_1751), .Z
		(n_1759));
	notech_and4 i_66077232(.A(n_1793), .B(n_2894), .C(n_2136), .D(n_3152), .Z
		(n_1757));
	notech_and4 i_65977233(.A(n_2609), .B(n_2928), .C(n_1792), .D(n_2629), .Z
		(n_1751));
	notech_ao4 i_65877234(.A(n_34143), .B(n_59585), .C(n_34142), .D(n_4072),
		 .Z(n_1745));
	notech_ao4 i_65677235(.A(n_34145), .B(n_1802), .C(n_2124), .D(n_59603), 
		.Z(n_1744));
	notech_and4 i_66277230(.A(n_34187), .B(n_69852396), .C(n_34030), .D(n_2365
		), .Z(n_1741));
	notech_and4 i_66177231(.A(n_4056), .B(n_4036), .C(n_872), .D(n_34070), .Z
		(n_1738));
	notech_and3 i_31377847(.A(n_4014), .B(n_208153600), .C(n_34049), .Z(n_1734
		));
	notech_and4 i_46577391(.A(n_2894), .B(n_4055), .C(n_1725), .D(n_1699), .Z
		(n_1730));
	notech_and4 i_46077395(.A(n_4030), .B(n_2569), .C(n_1950), .D(n_34043), 
		.Z(n_1725));
	notech_nand3 i_25477852(.A(n_2076), .B(n_4055), .C(n_2620), .Z(n_1722)
		);
	notech_ao3 i_46477392(.A(n_1719), .B(n_1714), .C(n_1640), .Z(n_1721));
	notech_and4 i_45977396(.A(n_4031), .B(n_1014), .C(n_3993), .D(n_34071), 
		.Z(n_1719));
	notech_and4 i_45877397(.A(n_4026), .B(n_2760), .C(n_2479), .D(n_2690), .Z
		(n_1714));
	notech_and4 i_31277849(.A(n_4007), .B(n_4047), .C(n_2340), .D(n_2609), .Z
		(n_1709));
	notech_and4 i_11677864(.A(n_4086), .B(n_2538), .C(n_34073), .D(n_1704), 
		.Z(n_1708));
	notech_and3 i_8177867(.A(n_4002), .B(n_4076), .C(n_4027), .Z(n_1704));
	notech_and4 i_73577817(.A(n_34063), .B(n_1958), .C(n_2377), .D(n_34042),
		 .Z(n_1702));
	notech_and2 i_62277829(.A(n_2365), .B(n_34040), .Z(n_1699));
	notech_and4 i_13977679(.A(n_1801), .B(n_3402), .C(n_1694), .D(n_4093), .Z
		(n_1695));
	notech_and4 i_13777681(.A(n_2664), .B(n_2637), .C(n_2357), .D(n_3124), .Z
		(n_1694));
	notech_or4 i_13877680(.A(n_1795), .B(n_4024), .C(n_1626), .D(n_1625), .Z
		(n_1689));
	notech_and4 i_12577693(.A(n_2611), .B(n_2949), .C(n_2166), .D(n_2463), .Z
		(n_1684));
	notech_and4 i_12677692(.A(n_3013), .B(n_2480), .C(n_2729), .D(n_2959), .Z
		(n_1681));
	notech_ao3 i_8777724(.A(n_2743), .B(n_2623), .C(n_1675), .Z(n_1676));
	notech_nand3 i_32677845(.A(n_2019), .B(n_1616), .C(n_1618), .Z(n_1675)
		);
	notech_and4 i_8577726(.A(n_1671), .B(n_1668), .C(n_1664), .D(n_1661), .Z
		(n_1673));
	notech_and4 i_8077729(.A(n_247296910), .B(n_2045), .C(n_2591), .D(n_4030
		), .Z(n_1671));
	notech_and4 i_7977730(.A(n_2588), .B(n_3360), .C(n_2627), .D(n_34031), .Z
		(n_1668));
	notech_and4 i_7877731(.A(n_2744), .B(n_2140), .C(n_2516), .D(n_1942), .Z
		(n_1664));
	notech_ao3 i_7777732(.A(n_34015), .B(n_1619), .C(n_34164), .Z(n_1661));
	notech_and4 i_5977748(.A(n_4048), .B(n_164996906), .C(n_2036), .D(n_1653
		), .Z(n_1654));
	notech_and4 i_5777750(.A(n_34187), .B(n_2831), .C(n_2450), .D(n_2426), .Z
		(n_1653));
	notech_and2 i_5077756(.A(n_2398), .B(n_1834), .Z(n_164996906));
	notech_and4 i_5877749(.A(n_1644), .B(n_2305), .C(n_1612), .D(n_3984), .Z
		(n_1647));
	notech_ao4 i_5377753(.A(n_2166), .B(n_2006), .C(n_4071), .D(n_1965), .Z(n_1644
		));
	notech_nand3 i_52377838(.A(n_4025), .B(n_2629), .C(n_34074), .Z(n_1640)
		);
	notech_and4 i_50277891(.A(n_1770), .B(n_1789), .C(n_1709), .D(n_3197), .Z
		(n_1639));
	notech_or2 i_77377146(.A(n_2151), .B(n_59511), .Z(n_1638));
	notech_or2 i_71177197(.A(n_3958), .B(n_2359), .Z(n_1637));
	notech_nand3 i_55377896(.A(n_1762), .B(n_1734), .C(n_1629), .Z(\udeco[33] 
		));
	notech_nand2 i_64477243(.A(modrm[4]), .B(n_221898892), .Z(n_1629));
	notech_and4 i_60377904(.A(n_1730), .B(n_1709), .C(n_1708), .D(n_1721), .Z
		(n_1628));
	notech_or4 i_77677933(.A(n_1689), .B(n_1621), .C(n_34183), .D(n_2102), .Z
		(\udeco[110] ));
	notech_and2 i_12977689(.A(adz), .B(n_34174), .Z(n_1626));
	notech_and2 i_12877690(.A(adz), .B(n_34069), .Z(n_1625));
	notech_and4 i_377803(.A(n_2484), .B(n_1684), .C(n_1681), .D(n_1995), .Z(n_1622
		));
	notech_and2 i_13077688(.A(opz[2]), .B(n_34208), .Z(n_1621));
	notech_and4 i_91577936(.A(n_1676), .B(n_1673), .C(n_34032), .D(n_2435), 
		.Z(n_1620));
	notech_or4 i_6877740(.A(n_2289), .B(n_59434), .C(n_59452), .D(n_34136), 
		.Z(n_1619));
	notech_or4 i_6577743(.A(n_2311), .B(n_59527), .C(n_59511), .D(n_34136), 
		.Z(n_1618));
	notech_nao3 i_6677742(.A(n_59527), .B(n_59538), .C(n_3277), .Z(n_1616)
		);
	notech_and4 i_94377937(.A(n_1654), .B(n_1647), .C(n_1613), .D(n_1606), .Z
		(n_1614));
	notech_nand2 i_4777759(.A(modrm[1]), .B(n_34209), .Z(n_1613));
	notech_or2 i_4577761(.A(n_4070), .B(n_59585), .Z(n_1612));
	notech_and4 i_077806(.A(n_4034), .B(n_1865), .C(n_1604), .D(n_2883), .Z(n_1608
		));
	notech_nand3 i_62507(.A(n_2398), .B(n_2380), .C(n_34036), .Z(\udeco[4] )
		);
	notech_and4 i_62740(.A(n_2366), .B(n_1960), .C(n_34073), .D(n_122998063)
		, .Z(udeco_73101168));
	notech_and2 i_1077796(.A(modrm[4]), .B(n_34093), .Z(n_118498020));
	notech_or4 i_62771(.A(n_4024), .B(n_214998833), .C(n_3971), .D(n_118498020
		), .Z(\udeco[84] ));
	notech_and2 i_1377793(.A(n_59479), .B(n_34093), .Z(n_118598021));
	notech_or4 i_62776(.A(n_3971), .B(n_4045), .C(n_118598021), .D(n_123498067
		), .Z(\udeco[85] ));
	notech_nao3 i_10377878(.A(n_1960), .B(n_3998), .C(n_4057), .Z(\udeco[88] 
		));
	notech_or2 i_62788(.A(\udeco[88] ), .B(\udeco[5] ), .Z(\udeco[89] ));
	notech_or4 i_6977877(.A(n_34132), .B(\udeco[5] ), .C(n_34108), .D(n_3971
		), .Z(\udeco[91] ));
	notech_nao3 i_62791(.A(n_34047), .B(n_34075), .C(n_34139), .Z(\udeco[92] 
		));
	notech_nao3 i_11377876(.A(n_3998), .B(n_34047), .C(n_34139), .Z(\udeco[90] 
		));
	notech_or2 i_62793(.A(n_4057), .B(\udeco[90] ), .Z(\udeco[93] ));
	notech_or2 i_62794(.A(n_4057), .B(\udeco[91] ), .Z(\udeco[95] ));
	notech_nao3 i_62795(.A(n_3998), .B(n_1960), .C(n_4010), .Z(\udeco[96] )
		);
	notech_or2 i_62797(.A(n_4010), .B(\udeco[88] ), .Z(\udeco[98] ));
	notech_or4 i_62799(.A(n_4024), .B(n_4057), .C(n_3971), .D(n_3985), .Z(\udeco[100] 
		));
	notech_and4 i_62800(.A(n_34148), .B(n_2623), .C(n_1960), .D(n_34075), .Z
		(udeco_101101167));
	notech_or4 i_62801(.A(n_4018), .B(n_3950), .C(\udeco[88] ), .D(n_4010), 
		.Z(\udeco[102] ));
	notech_nao3 i_28677938(.A(n_34210), .B(n_124598078), .C(n_124098073), .Z
		(\udeco[127] ));
	notech_nand3 i_277804(.A(n_2099), .B(n_3736), .C(n_1905), .Z(n_118698022
		));
	notech_nor2 i_9077721(.A(n_1984), .B(n_34193), .Z(n_118798023));
	notech_nand2 i_9177720(.A(n_59479), .B(n_3956), .Z(n_118898024));
	notech_and2 i_9277719(.A(modrm[2]), .B(n_118698022), .Z(n_118998025));
	notech_or4 i_88077935(.A(n_124098073), .B(n_126198091), .C(n_125498085),
		 .D(n_125198082), .Z(\udeco[118] ));
	notech_or4 i_69877934(.A(n_4024), .B(n_4057), .C(n_1675), .D(n_34085), .Z
		(\udeco[115] ));
	notech_or4 i_56177932(.A(n_128798112), .B(n_34088), .C(n_127398100), .D(n_207953599
		), .Z(\udeco[107] ));
	notech_nao3 i_16277659(.A(n_59538), .B(n_2397), .C(n_2403), .Z(n_119098026
		));
	notech_or4 i_16477658(.A(n_59416), .B(n_4090), .C(n_2315), .D(modrm[5]),
		 .Z(n_119198027));
	notech_nand2 i_16877655(.A(opz[2]), .B(n_34059), .Z(n_119298028));
	notech_nand3 i_20277931(.A(n_119198027), .B(n_119098026), .C(n_129798121
		), .Z(\udeco[106] ));
	notech_or2 i_17877647(.A(n_2278), .B(n_2052), .Z(n_119498029));
	notech_nand2 i_17977646(.A(opz[1]), .B(n_34059), .Z(n_119598030));
	notech_nand3 i_72577930(.A(n_119198027), .B(n_130998128), .C(n_119098026
		), .Z(\udeco[105] ));
	notech_and4 i_20577929(.A(n_1969), .B(n_2623), .C(n_1960), .D(n_34148), 
		.Z(udeco_103101166));
	notech_and2 i_19277633(.A(modrm[7]), .B(n_34093), .Z(n_119698031));
	notech_or4 i_72177928(.A(n_34139), .B(n_214998833), .C(n_3971), .D(n_119698031
		), .Z(\udeco[87] ));
	notech_and2 i_19577630(.A(modrm[6]), .B(n_34093), .Z(n_119798032));
	notech_or4 i_72110227(.A(n_34139), .B(n_214998833), .C(n_3971), .D(n_119798032
		), .Z(\udeco[86] ));
	notech_or4 i_62798(.A(n_4024), .B(n_4057), .C(n_4010), .D(n_3971), .Z(\udeco[99] 
		));
	notech_nand2 i_19977626(.A(modrm[3]), .B(n_34093), .Z(n_119898033));
	notech_or4 i_71877927(.A(n_214998833), .B(n_4009), .C(\udeco[99] ), .D(n_131598134
		), .Z(\udeco[83] ));
	notech_nand2 i_21177619(.A(modrm[2]), .B(n_34093), .Z(n_120198036));
	notech_nand3 i_71577926(.A(n_131898137), .B(n_131798136), .C(n_132298139
		), .Z(\udeco[82] ));
	notech_or4 i_21777613(.A(n_2386), .B(n_59493), .C(n_59603), .D(n_34080),
		 .Z(n_120298037));
	notech_or4 i_22077611(.A(n_59558), .B(n_2182), .C(n_59594), .D(n_59470),
		 .Z(n_120498039));
	notech_and2 i_22177610(.A(modrm[1]), .B(n_34093), .Z(n_120598040));
	notech_or4 i_71277925(.A(n_34186), .B(n_120598040), .C(n_34139), .D(n_133198145
		), .Z(\udeco[81] ));
	notech_or4 i_22277924(.A(n_4011), .B(n_4018), .C(\udeco[91] ), .D(n_34090
		), .Z(\udeco[80] ));
	notech_nao3 i_10477871(.A(n_122998063), .B(n_1960), .C(n_133798149), .Z(\udeco[74] 
		));
	notech_or4 i_21610230(.A(n_34035), .B(n_34034), .C(\udeco[74] ), .D(n_3968
		), .Z(\udeco[78] ));
	notech_nao3 i_20510233(.A(n_34077), .B(n_34210), .C(n_133898150), .Z(\udeco[77] 
		));
	notech_or4 i_22877923(.A(n_133898150), .B(n_1326), .C(n_3971), .D(n_3978
		), .Z(\udeco[75] ));
	notech_nand3 i_22210242(.A(n_131798136), .B(n_135398160), .C(n_122998063
		), .Z(\udeco[72] ));
	notech_or4 i_70977922(.A(n_124098073), .B(n_136298168), .C(n_34034), .D(n_3969
		), .Z(\udeco[70] ));
	notech_nao3 i_11477870(.A(n_34060), .B(n_34042), .C(n_136298168), .Z(\udeco[71] 
		));
	notech_or4 i_70577921(.A(n_4009), .B(n_3969), .C(n_136298168), .D(n_3968
		), .Z(\udeco[68] ));
	notech_or4 i_20977920(.A(n_34034), .B(\udeco[71] ), .C(\udeco[5] ), .D(n_214998833
		), .Z(\udeco[67] ));
	notech_or4 i_20210249(.A(n_4045), .B(n_136298168), .C(n_136398169), .D(n_34035
		), .Z(\udeco[69] ));
	notech_or2 i_70277919(.A(n_4057), .B(\udeco[69] ), .Z(\udeco[66] ));
	notech_or4 i_69810253(.A(n_135698162), .B(n_34113), .C(n_136098166), .D(n_137398178
		), .Z(\udeco[65] ));
	notech_or4 i_69810257(.A(n_135698162), .B(n_34113), .C(n_136098166), .D(n_137798182
		), .Z(\udeco[64] ));
	notech_or4 i_69477918(.A(n_4054), .B(n_139398195), .C(n_4015), .D(n_138998191
		), .Z(\udeco[63] ));
	notech_or4 i_68377917(.A(n_121198045), .B(n_139398195), .C(n_124098073),
		 .D(n_138998191), .Z(\udeco[62] ));
	notech_nao3 i_68977916(.A(n_140098202), .B(n_34092), .C(n_124098073), .Z
		(\udeco[61] ));
	notech_or4 i_59277915(.A(n_140598206), .B(n_140298204), .C(n_4015), .D(n_4054
		), .Z(\udeco[60] ));
	notech_nand3 i_68310262(.A(n_138498186), .B(n_141298213), .C(n_34091), .Z
		(\udeco[59] ));
	notech_nand3 i_67877914(.A(n_2579), .B(n_138498186), .C(n_142398222), .Z
		(\udeco[58] ));
	notech_or4 i_67277913(.A(n_135898164), .B(n_135798163), .C(n_140298204),
		 .D(n_142698224), .Z(\udeco[57] ));
	notech_ao4 i_105877809(.A(n_2210), .B(n_3959), .C(n_34144), .D(n_34007),
		 .Z(n_121198045));
	notech_or4 i_66777912(.A(n_142998227), .B(n_121198045), .C(n_143298230),
		 .D(n_140298204), .Z(\udeco[56] ));
	notech_or4 i_66210267(.A(n_144198238), .B(n_4011), .C(n_1640), .D(n_34176
		), .Z(\udeco[55] ));
	notech_nao3 i_65777911(.A(n_143898235), .B(n_144898245), .C(n_124098073)
		, .Z(\udeco[54] ));
	notech_or4 i_65277910(.A(n_34097), .B(n_146198257), .C(n_221898892), .D(n_34113
		), .Z(\udeco[53] ));
	notech_or4 i_64577909(.A(n_146498260), .B(n_34176), .C(n_34096), .D(n_122898062
		), .Z(\udeco[52] ));
	notech_or4 i_64177908(.A(n_135898164), .B(n_135798163), .C(n_34176), .D(n_148398273
		), .Z(\udeco[51] ));
	notech_ao3 i_39477457(.A(n_34201), .B(modrm[3]), .C(n_2113), .Z(n_121298046
		));
	notech_or4 i_63577907(.A(n_34113), .B(n_34097), .C(n_124098073), .D(n_149998287
		), .Z(\udeco[50] ));
	notech_or4 i_41177440(.A(n_2118), .B(n_59544), .C(n_59511), .D(n_59461),
		 .Z(n_121398047));
	notech_nao3 i_61977906(.A(n_150998296), .B(n_143898235), .C(n_34176), .Z
		(\udeco[48] ));
	notech_or4 i_62377905(.A(n_152498311), .B(n_151298299), .C(n_139198193),
		 .D(n_34081), .Z(\udeco[47] ));
	notech_or4 i_61910271(.A(n_1640), .B(n_34102), .C(n_152798313), .D(n_153698321
		), .Z(\udeco[46] ));
	notech_or4 i_61577903(.A(n_155198331), .B(n_151798304), .C(n_154998329),
		 .D(n_34081), .Z(\udeco[44] ));
	notech_or4 i_35377902(.A(n_221898892), .B(n_34078), .C(n_34107), .D(n_157298349
		), .Z(\udeco[43] ));
	notech_or2 i_49877358(.A(n_5254), .B(n_59443), .Z(n_121498048));
	notech_or4 i_60977901(.A(n_34107), .B(n_157498351), .C(n_159198365), .D(n_34082
		), .Z(\udeco[42] ));
	notech_or4 i_60310278(.A(n_34176), .B(n_151798304), .C(n_161098380), .D(n_135998165
		), .Z(\udeco[41] ));
	notech_ao4 i_477802(.A(n_4065), .B(n_2320), .C(n_59425), .D(n_2371), .Z(n_121898052
		));
	notech_nor2 i_54377320(.A(n_5254), .B(n_34200), .Z(n_121998053));
	notech_nor2 i_54477319(.A(n_2275), .B(n_121898052), .Z(n_122098054));
	notech_or4 i_59677900(.A(n_161698385), .B(n_162598391), .C(n_152798313),
		 .D(n_151298299), .Z(\udeco[40] ));
	notech_nand3 i_59210283(.A(n_163998402), .B(n_163698399), .C(n_163298396
		), .Z(\udeco[39] ));
	notech_or4 i_58777899(.A(n_164898411), .B(n_164598408), .C(n_155198331),
		 .D(n_34112), .Z(\udeco[38] ));
	notech_nao3 i_57577898(.A(n_1734), .B(n_166598425), .C(n_221898892), .Z(\udeco[36] 
		));
	notech_nao3 i_61077266(.A(n_59452), .B(n_59538), .C(n_2564), .Z(n_122198055
		));
	notech_and4 i_56877897(.A(n_1193), .B(n_168398442), .C(n_167598435), .D(n_1734
		), .Z(udeco_35101165));
	notech_nand3 i_53977895(.A(n_170798463), .B(n_169198450), .C(n_1960), .Z
		(\udeco[31] ));
	notech_or4 i_53177894(.A(n_221898892), .B(n_34125), .C(n_204853574), .D(n_172798479
		), .Z(\udeco[30] ));
	notech_and4 i_52277893(.A(n_169098449), .B(n_1770), .C(n_174398492), .D(n_3109
		), .Z(udeco_29101164));
	notech_and4 i_51277892(.A(n_175098498), .B(n_176298508), .C(n_3510), .D(n_169198450
		), .Z(udeco_28101163));
	notech_or4 i_78877133(.A(n_2347), .B(n_2338), .C(n_3961), .D(n_59621), .Z
		(n_122298056));
	notech_nao3 i_46177890(.A(n_179198527), .B(n_1699), .C(n_34121), .Z(\udeco[22] 
		));
	notech_and4 i_45177889(.A(n_179498530), .B(n_182098553), .C(n_1925), .D(n_222298895
		), .Z(udeco_21101162));
	notech_or4 i_42477888(.A(n_34125), .B(n_34176), .C(n_34124), .D(n_184398571
		), .Z(\udeco[19] ));
	notech_and4 i_37277887(.A(n_185998586), .B(n_185598583), .C(n_185398581)
		, .D(n_3403), .Z(udeco_15101161));
	notech_and4 i_36977886(.A(n_187298596), .B(n_186798593), .C(n_151898305)
		, .D(n_3403), .Z(udeco_14101160));
	notech_nor2 i_88677040(.A(n_3954), .B(n_3958), .Z(n_122398057));
	notech_and4 i_35310321(.A(n_188098604), .B(n_187798601), .C(n_189298616)
		, .D(n_34049), .Z(udeco_12101159));
	notech_nand2 i_29510326(.A(n_68), .B(n_34133), .Z(\udeco[6] ));
	notech_or2 i_91277014(.A(n_2398), .B(n_59511), .Z(n_122498058));
	notech_nand3 i_29077885(.A(n_122498058), .B(n_34057), .C(n_34133), .Z(\udeco[3] 
		));
	notech_nor2 i_91677011(.A(n_2398), .B(n_59470), .Z(n_122598059));
	notech_or4 i_29010330(.A(n_1967), .B(n_34134), .C(n_122598059), .D(n_189798621
		), .Z(\udeco[2] ));
	notech_nor2 i_92077007(.A(n_2398), .B(n_59585), .Z(n_122698060));
	notech_or4 i_28610335(.A(n_190098623), .B(n_4006), .C(n_122698060), .D(n_34135
		), .Z(\udeco[1] ));
	notech_nand2 i_35477844(.A(n_1958), .B(n_4066), .Z(n_122898062));
	notech_and3 i_68677824(.A(n_3992), .B(n_3876), .C(n_34083), .Z(n_122998063
		));
	notech_nao3 i_1577791(.A(n_1950), .B(n_2380), .C(n_214998833), .Z(n_123498067
		));
	notech_nao3 i_6377868(.A(n_34060), .B(n_34058), .C(n_1640), .Z(n_124098073
		));
	notech_and4 i_3477772(.A(n_4017), .B(n_1920), .C(n_2450), .D(n_34076), .Z
		(n_124398076));
	notech_and4 i_3677770(.A(n_4048), .B(n_2195), .C(n_124398076), .D(n_2435
		), .Z(n_124598078));
	notech_or4 i_10077711(.A(n_34101), .B(n_4003), .C(n_1180), .D(n_3985), .Z
		(n_125198082));
	notech_or4 i_10177710(.A(n_222598898), .B(n_34169), .C(n_34173), .D(n_4080
		), .Z(n_125498085));
	notech_and4 i_9977712(.A(n_2516), .B(n_3733), .C(n_2332), .D(n_118898024
		), .Z(n_125898089));
	notech_or4 i_10677707(.A(n_118798023), .B(n_118998025), .C(n_3974), .D(n_34084
		), .Z(n_126198091));
	notech_and4 i_11277701(.A(n_1543), .B(n_1923), .C(n_4061), .D(n_1545), .Z
		(n_126998096));
	notech_or4 i_15277667(.A(n_222998902), .B(n_34086), .C(n_1262), .D(n_34087
		), .Z(n_127398100));
	notech_and4 i_15377666(.A(n_4084), .B(n_3991), .C(n_2162), .D(n_4004), .Z
		(n_127698103));
	notech_nand2 i_14477674(.A(n_4061), .B(n_2792), .Z(n_128198108));
	notech_or4 i_15477665(.A(n_4024), .B(n_34061), .C(n_34048), .D(n_128198108
		), .Z(n_128398110));
	notech_or4 i_16077661(.A(n_34179), .B(n_4009), .C(n_128398110), .D(n_34121
		), .Z(n_128798112));
	notech_and4 i_17577650(.A(n_1678), .B(n_208398774), .C(n_2623), .D(n_34075
		), .Z(n_129698120));
	notech_and4 i_17677649(.A(n_129698120), .B(n_34060), .C(n_4087), .D(n_119298028
		), .Z(n_129798121));
	notech_and4 i_18577640(.A(n_4043), .B(n_4087), .C(n_1678), .D(n_208398774
		), .Z(n_130198123));
	notech_and3 i_18477641(.A(n_2049), .B(n_3998), .C(n_119598030), .Z(n_130798126
		));
	notech_and4 i_18777638(.A(n_119498029), .B(n_130798126), .C(n_130198123)
		, .D(n_2380), .Z(n_130998128));
	notech_nao3 i_20477624(.A(n_4093), .B(n_119898033), .C(n_34035), .Z(n_131598134
		));
	notech_and2 i_69177821(.A(n_2366), .B(n_34207), .Z(n_131798136));
	notech_ao4 i_21377617(.A(n_2383), .B(n_2167), .C(n_3963), .D(n_2182), .Z
		(n_131898137));
	notech_and4 i_21477616(.A(n_34077), .B(n_34073), .C(n_2357), .D(n_120198036
		), .Z(n_132298139));
	notech_ao4 i_22577607(.A(n_2383), .B(n_2182), .C(n_2167), .D(n_34136), .Z
		(n_133098144));
	notech_nand3 i_22777605(.A(n_120298037), .B(n_133098144), .C(n_34073), .Z
		(n_133198145));
	notech_ao4 i_23377601(.A(n_1953), .B(n_34198), .C(n_2577), .D(n_3935), .Z
		(n_133498147));
	notech_nao3 i_80377811(.A(n_2629), .B(n_1953), .C(n_4011), .Z(n_133798149
		));
	notech_nao3 i_16977858(.A(n_5254), .B(n_34083), .C(n_133798149), .Z(n_133898150
		));
	notech_and3 i_25077584(.A(n_3970), .B(n_120498039), .C(n_34143), .Z(n_134998156
		));
	notech_ao4 i_24977585(.A(n_34080), .B(n_2167), .C(n_59416), .D(n_2368), 
		.Z(n_135198158));
	notech_and4 i_25277582(.A(n_135198158), .B(n_2151), .C(n_34180), .D(n_134998156
		), .Z(n_135398160));
	notech_nand2 i_55177836(.A(n_2123), .B(n_4034), .Z(n_135698162));
	notech_or2 i_80577810(.A(n_135698162), .B(n_34113), .Z(n_135798163));
	notech_or2 i_25777579(.A(n_34068), .B(n_4024), .Z(n_135898164));
	notech_or4 i_15677861(.A(n_4024), .B(n_34068), .C(n_135698162), .D(n_34113
		), .Z(n_135998165));
	notech_nand3 i_64277827(.A(n_4056), .B(n_4044), .C(n_3964), .Z(n_136098166
		));
	notech_or4 i_235577807(.A(n_4091), .B(n_136098166), .C(n_135898164), .D(n_135798163
		), .Z(n_136298168));
	notech_or4 i_25977577(.A(n_4011), .B(n_1640), .C(n_4009), .D(n_3969), .Z
		(n_136398169));
	notech_nand3 i_65177825(.A(n_5254), .B(n_2377), .C(n_1958), .Z(n_136898174
		));
	notech_or2 i_73077819(.A(n_34068), .B(n_34108), .Z(n_136998175));
	notech_or4 i_27277565(.A(n_34132), .B(n_3978), .C(n_136998175), .D(n_136898174
		), .Z(n_137398178));
	notech_or4 i_27777560(.A(n_34132), .B(n_4091), .C(n_136998175), .D(n_133798149
		), .Z(n_137798182));
	notech_and4 i_8277866(.A(n_2094), .B(n_210398792), .C(n_2569), .D(n_1905
		), .Z(n_138498186));
	notech_and4 i_28577553(.A(n_3979), .B(n_34076), .C(n_34042), .D(n_1978),
		 .Z(n_138798189));
	notech_nand3 i_11777863(.A(n_138498186), .B(n_138798189), .C(n_1193), .Z
		(n_138998191));
	notech_and2 i_62077831(.A(n_34044), .B(n_34039), .Z(n_139098192));
	notech_or2 i_59777834(.A(n_4006), .B(n_4024), .Z(n_139198193));
	notech_or4 i_28877551(.A(n_4024), .B(n_4006), .C(n_4091), .D(n_34103), .Z
		(n_139398195));
	notech_and4 i_29777543(.A(n_2327), .B(n_2623), .C(n_34043), .D(n_2305), 
		.Z(n_139798199));
	notech_and4 i_30077540(.A(n_139798199), .B(n_131798136), .C(n_139098192)
		, .D(n_34091), .Z(n_140098202));
	notech_nand2 i_62177830(.A(n_2579), .B(n_138498186), .Z(n_140298204));
	notech_or4 i_30477536(.A(n_4006), .B(n_4091), .C(n_222498897), .D(n_34103
		), .Z(n_140598206));
	notech_and4 i_31177529(.A(n_1978), .B(n_34187), .C(n_2304), .D(n_1816), 
		.Z(n_141198212));
	notech_and4 i_31477528(.A(n_141198212), .B(n_1953), .C(n_2623), .D(n_34044
		), .Z(n_141298213));
	notech_and3 i_81477808(.A(n_34046), .B(n_34039), .C(n_2380), .Z(n_141598216
		));
	notech_and4 i_32177521(.A(n_139798199), .B(n_34187), .C(n_2357), .D(n_34094
		), .Z(n_142198220));
	notech_and4 i_32577518(.A(n_34091), .B(n_1193), .C(n_141598216), .D(n_142198220
		), .Z(n_142398222));
	notech_nao3 i_32977515(.A(n_34043), .B(n_139098192), .C(n_4091), .Z(n_142698224
		));
	notech_nao3 i_33577509(.A(n_1953), .B(n_1950), .C(n_4009), .Z(n_142998227
		));
	notech_or4 i_33677508(.A(n_4091), .B(n_2307), .C(n_34068), .D(n_2165), .Z
		(n_143298230));
	notech_and4 i_32277846(.A(n_4031), .B(n_69852396), .C(n_2304), .D(n_34057
		), .Z(n_143898235));
	notech_or4 i_34477500(.A(n_3986), .B(n_210198790), .C(n_34120), .D(n_34095
		), .Z(n_144198238));
	notech_and4 i_35077494(.A(n_34063), .B(n_34072), .C(n_2365), .D(n_1972),
		 .Z(n_144698243));
	notech_and4 i_35277492(.A(n_34149), .B(n_144698243), .C(n_34083), .D(n_34071
		), .Z(n_144898245));
	notech_nand2 i_35877488(.A(n_222798900), .B(n_4016), .Z(n_145198247));
	notech_and4 i_36477482(.A(n_2365), .B(n_2099), .C(n_2327), .D(n_34072), 
		.Z(n_145598251));
	notech_nao3 i_36777480(.A(n_145598251), .B(n_2380), .C(n_145198247), .Z(n_145698252
		));
	notech_or4 i_36677481(.A(n_4045), .B(n_210198790), .C(n_4091), .D(n_34069
		), .Z(n_145998255));
	notech_or4 i_37077478(.A(n_145998255), .B(n_34179), .C(n_4009), .D(n_145698252
		), .Z(n_146198257));
	notech_or4 i_37877472(.A(n_34181), .B(n_34165), .C(n_34167), .D(n_4024),
		 .Z(n_146498260));
	notech_and4 i_37977471(.A(n_3360), .B(n_2099), .C(n_69852396), .D(n_34042
		), .Z(n_146998263));
	notech_and4 i_38877463(.A(n_222798900), .B(n_1737), .C(n_5254), .D(n_4031
		), .Z(n_147998270));
	notech_and4 i_38977462(.A(n_3982), .B(n_147998270), .C(n_2614), .D(n_34057
		), .Z(n_148198271));
	notech_nand3 i_39177460(.A(n_148198271), .B(n_141598216), .C(n_1702), .Z
		(n_148398273));
	notech_or4 i_39577456(.A(n_4023), .B(n_34166), .C(n_34179), .D(n_3990), 
		.Z(n_148698276));
	notech_or4 i_40477447(.A(n_121298046), .B(n_148698276), .C(n_1326), .D(n_4045
		), .Z(n_148898278));
	notech_or4 i_40377448(.A(n_4091), .B(n_3968), .C(n_4088), .D(n_34099), .Z
		(n_149598284));
	notech_or4 i_40577446(.A(n_209698786), .B(n_4052), .C(n_145198247), .D(n_149598284
		), .Z(n_149798285));
	notech_or4 i_40877443(.A(n_148898278), .B(n_34120), .C(n_149798285), .D(n_135698162
		), .Z(n_149998287));
	notech_and4 i_41777434(.A(n_3979), .B(n_2366), .C(n_34187), .D(n_210098789
		), .Z(n_150398291));
	notech_ao3 i_41677435(.A(n_210498793), .B(n_121398047), .C(n_222398896),
		 .Z(n_150798294));
	notech_and4 i_41977432(.A(n_150398291), .B(n_150798294), .C(n_2380), .D(n_34073
		), .Z(n_150998296));
	notech_nand3 i_25377853(.A(n_843), .B(n_4047), .C(n_4067), .Z(n_151298299
		));
	notech_and4 i_42877424(.A(n_4051), .B(n_4007), .C(n_4025), .D(n_4085), .Z
		(n_151698303));
	notech_nand3 i_17477857(.A(n_3993), .B(n_4055), .C(n_151698303), .Z(n_151798304
		));
	notech_and2 i_73777816(.A(n_34065), .B(n_34050), .Z(n_151898305));
	notech_and4 i_43277420(.A(n_4019), .B(n_1014), .C(n_2116), .D(n_34071), 
		.Z(n_152198308));
	notech_nao3 i_43377419(.A(n_34060), .B(n_152198308), .C(n_4088), .Z(n_152298309
		));
	notech_or4 i_43677416(.A(n_4035), .B(n_151798304), .C(n_4033), .D(n_152298309
		), .Z(n_152498311));
	notech_nand2 i_73877815(.A(n_4085), .B(n_1704), .Z(n_152798313));
	notech_and4 i_44377409(.A(n_3982), .B(n_1623), .C(n_34060), .D(n_34072),
		 .Z(n_153398318));
	notech_and4 i_44477408(.A(n_3064), .B(n_3360), .C(n_153398318), .D(n_34039
		), .Z(n_153498319));
	notech_or2 i_44677406(.A(n_139198193), .B(n_34118), .Z(n_153698321));
	notech_and4 i_47377383(.A(n_2017), .B(n_34050), .C(n_34065), .D(n_3980),
		 .Z(n_154298324));
	notech_and4 i_47477382(.A(n_5254), .B(n_4019), .C(n_3064), .D(n_2304), .Z
		(n_154798327));
	notech_nao3 i_47677380(.A(n_154798327), .B(n_154298324), .C(n_151298299)
		, .Z(n_154998329));
	notech_or4 i_36577843(.A(n_4050), .B(n_4054), .C(n_4059), .D(n_4024), .Z
		(n_155198331));
	notech_or4 i_48777369(.A(n_4023), .B(n_4059), .C(n_34182), .D(n_223098903
		), .Z(n_155898337));
	notech_or4 i_49277364(.A(n_1987), .B(n_34153), .C(n_1722), .D(n_155898337
		), .Z(n_156098339));
	notech_nand3 i_48377373(.A(n_1798), .B(n_1796), .C(n_4025), .Z(n_156398341
		));
	notech_or4 i_48977367(.A(n_2307), .B(n_222398896), .C(n_34166), .D(n_34190
		), .Z(n_156798345));
	notech_or4 i_49177365(.A(n_34181), .B(n_4050), .C(n_156398341), .D(n_156798345
		), .Z(n_156898346));
	notech_or4 i_49577361(.A(n_156098339), .B(n_156898346), .C(n_1086), .D(n_34118
		), .Z(n_157298349));
	notech_or4 i_51077347(.A(n_4035), .B(n_4033), .C(n_34068), .D(n_34108), 
		.Z(n_157498351));
	notech_and4 i_50677351(.A(n_210398792), .B(n_69852396), .C(n_2365), .D(n_3993
		), .Z(n_158398357));
	notech_and4 i_50877349(.A(n_3994), .B(n_3996), .C(n_158398357), .D(n_121498048
		), .Z(n_158498358));
	notech_and4 i_50777350(.A(n_2623), .B(n_34076), .C(n_34077), .D(n_4030),
		 .Z(n_158898362));
	notech_and4 i_51377345(.A(n_158898362), .B(n_141598216), .C(n_2116), .D(n_34060
		), .Z(n_159098364));
	notech_nand3 i_51577343(.A(n_222298895), .B(n_158498358), .C(n_159098364
		), .Z(n_159198365));
	notech_ao4 i_52877332(.A(n_5254), .B(n_34201), .C(n_4065), .D(n_2018), .Z
		(n_159498367));
	notech_and4 i_52977331(.A(n_1728), .B(n_4032), .C(n_4056), .D(n_4082), .Z
		(n_159798370));
	notech_and4 i_53077330(.A(n_2760), .B(n_3064), .C(n_214598830), .D(n_34040
		), .Z(n_160198374));
	notech_and4 i_53277329(.A(n_2569), .B(n_34043), .C(n_222798900), .D(n_4086
		), .Z(n_160698377));
	notech_and4 i_53577326(.A(n_160698377), .B(n_160198374), .C(n_159798370)
		, .D(n_159498367), .Z(n_160898379));
	notech_nand2 i_53677325(.A(n_160898379), .B(n_1704), .Z(n_161098380));
	notech_or4 i_55677309(.A(n_156398341), .B(n_4006), .C(n_34184), .D(n_122098054
		), .Z(n_161698385));
	notech_and4 i_55277312(.A(n_1014), .B(n_1951), .C(n_4007), .D(n_1815), .Z
		(n_162298390));
	notech_or4 i_55577310(.A(n_4001), .B(n_2164), .C(n_121998053), .D(n_34109
		), .Z(n_162598391));
	notech_and4 i_57177297(.A(n_2036), .B(n_2569), .C(n_34042), .D(n_34207),
		 .Z(n_163298396));
	notech_and4 i_56977299(.A(n_1332), .B(n_3967), .C(n_212098806), .D(n_211798804
		), .Z(n_163698399));
	notech_and4 i_57077298(.A(n_2176), .B(n_3979), .C(n_901), .D(n_3965), .Z
		(n_163998402));
	notech_and4 i_58077289(.A(n_2176), .B(n_901), .C(n_894), .D(n_212498809)
		, .Z(n_164498407));
	notech_nand3 i_58277287(.A(n_2036), .B(n_164498407), .C(n_34073), .Z(n_164598408
		));
	notech_or4 i_58177288(.A(n_34173), .B(n_1987), .C(n_34181), .D(n_4060), 
		.Z(n_164898411));
	notech_and4 i_60177273(.A(n_2569), .B(n_2015), .C(n_214598830), .D(n_34044
		), .Z(n_165398415));
	notech_and4 i_59877275(.A(n_1329), .B(n_3977), .C(n_861), .D(n_1537), .Z
		(n_165898418));
	notech_and4 i_59177279(.A(n_2663), .B(n_2327), .C(n_214098825), .D(n_853
		), .Z(n_165998419));
	notech_and4 i_60277272(.A(n_3967), .B(n_3965), .C(n_165998419), .D(n_165898418
		), .Z(n_166298422));
	notech_and4 i_60677269(.A(n_166298422), .B(n_165398415), .C(n_34104), .D
		(n_3107), .Z(n_166598425));
	notech_and4 i_63077253(.A(n_69852396), .B(n_1816), .C(n_34077), .D(n_34072
		), .Z(n_166998429));
	notech_and4 i_62777256(.A(n_222698899), .B(n_4051), .C(n_4029), .D(n_872
		), .Z(n_167398433));
	notech_and4 i_63377250(.A(n_167398433), .B(n_166998429), .C(n_2305), .D(n_122198055
		), .Z(n_167598435));
	notech_and4 i_61477262(.A(n_3062), .B(n_2500), .C(n_3736), .D(n_1905), .Z
		(n_167798437));
	notech_and4 i_62977254(.A(n_3994), .B(n_1593), .C(n_1329), .D(n_34070), 
		.Z(n_168298441));
	notech_and4 i_63277251(.A(n_2076), .B(n_4036), .C(n_167798437), .D(n_168298441
		), .Z(n_168398442));
	notech_and4 i_68177215(.A(n_3970), .B(n_1806), .C(n_730), .D(n_3079), .Z
		(n_168898447));
	notech_and4 i_68477213(.A(n_733), .B(n_738), .C(n_168898447), .D(n_3197)
		, .Z(n_169098449));
	notech_and2 i_26977851(.A(n_3109), .B(n_169098449), .Z(n_169198450));
	notech_and4 i_70177204(.A(n_2327), .B(n_4032), .C(n_853), .D(n_214098825
		), .Z(n_169498453));
	notech_and4 i_69977206(.A(n_717), .B(n_2246), .C(n_4014), .D(n_4013), .Z
		(n_169798456));
	notech_and3 i_69277210(.A(n_1984), .B(n_1801), .C(n_1993), .Z(n_169898457
		));
	notech_and4 i_70377203(.A(n_4034), .B(n_169798456), .C(n_4085), .D(n_169898457
		), .Z(n_170398460));
	notech_and4 i_70777200(.A(n_222298895), .B(n_169498453), .C(n_208153600)
		, .D(n_170398460), .Z(n_170798463));
	notech_and4 i_72377189(.A(n_214398828), .B(n_3992), .C(n_202798726), .D(n_692
		), .Z(n_171698469));
	notech_nand3 i_72777186(.A(n_171698469), .B(n_2627), .C(n_34046), .Z(n_171798470
		));
	notech_and4 i_72477188(.A(n_709), .B(n_719), .C(n_703), .D(n_4008), .Z(n_172198473
		));
	notech_and4 i_72677187(.A(n_2760), .B(n_4032), .C(n_3143), .D(n_3980), .Z
		(n_172498476));
	notech_or4 i_73377182(.A(n_34116), .B(n_171798470), .C(n_155198331), .D(n_34115
		), .Z(n_172798479));
	notech_and4 i_74777171(.A(n_4041), .B(n_4036), .C(n_720), .D(n_673), .Z(n_173398483
		));
	notech_and4 i_74877170(.A(n_214398828), .B(n_4028), .C(n_1718), .D(n_222898901
		), .Z(n_173898487));
	notech_and2 i_74577173(.A(n_1332), .B(n_212098806), .Z(n_174098489));
	notech_and4 i_75177167(.A(n_222698899), .B(n_4029), .C(n_174098489), .D(n_173898487
		), .Z(n_174298491));
	notech_and4 i_75277166(.A(n_173398483), .B(n_174298491), .C(n_1950), .D(n_34047
		), .Z(n_174398492));
	notech_and4 i_76377155(.A(n_2099), .B(n_4016), .C(n_4026), .D(n_2538), .Z
		(n_174798496));
	notech_and4 i_76877151(.A(n_4055), .B(n_2894), .C(n_174798496), .D(n_1770
		), .Z(n_175098498));
	notech_and4 i_76177157(.A(n_1290), .B(n_4014), .C(n_720), .D(n_1999), .Z
		(n_175698502));
	notech_and4 i_76277156(.A(n_1718), .B(n_3967), .C(n_34070), .D(n_2760), 
		.Z(n_175998505));
	notech_and4 i_77077149(.A(n_175998505), .B(n_175698502), .C(n_1960), .D(n_34049
		), .Z(n_176298508));
	notech_and2 i_77577813(.A(n_1434), .B(n_122298056), .Z(n_176698511));
	notech_and4 i_79877124(.A(n_4053), .B(n_200298705), .C(n_4027), .D(n_1615
		), .Z(n_177598517));
	notech_and4 i_80177121(.A(n_493), .B(n_4084), .C(n_177598517), .D(n_497)
		, .Z(n_177698518));
	notech_and2 i_79377128(.A(n_4038), .B(n_191198633), .Z(n_178198520));
	notech_and4 i_80077122(.A(n_1537), .B(n_2760), .C(n_2928), .D(n_2571), .Z
		(n_178798524));
	notech_and4 i_80277120(.A(n_178198520), .B(n_178798524), .C(n_2080), .D(n_1996
		), .Z(n_178998525));
	notech_and4 i_80877116(.A(n_177698518), .B(n_176698511), .C(n_3280), .D(n_178998525
		), .Z(n_179198527));
	notech_and4 i_82877097(.A(n_2928), .B(n_853), .C(n_730), .D(n_4047), .Z(n_179498530
		));
	notech_and4 i_82377102(.A(n_2678), .B(n_2791), .C(n_533), .D(n_2884), .Z
		(n_180098535));
	notech_and4 i_81277112(.A(n_2631), .B(n_1780), .C(n_2137), .D(n_2757), .Z
		(n_180398538));
	notech_and4 i_82577100(.A(n_2157), .B(n_2212), .C(n_4049), .D(n_2029), .Z
		(n_180798542));
	notech_and4 i_83077095(.A(n_574), .B(n_466), .C(n_180398538), .D(n_180798542
		), .Z(n_180898543));
	notech_and4 i_83377092(.A(n_4004), .B(n_2538), .C(n_180098535), .D(n_180898543
		), .Z(n_180998544));
	notech_and4 i_82677099(.A(n_3987), .B(n_537), .C(n_202098721), .D(n_1777
		), .Z(n_181298547));
	notech_and4 i_82777098(.A(n_3973), .B(n_4037), .C(n_1504), .D(n_4005), .Z
		(n_181798550));
	notech_and4 i_83677089(.A(n_181798550), .B(n_181298547), .C(n_2435), .D(n_180998544
		), .Z(n_182098553));
	notech_and4 i_85677069(.A(n_2398), .B(n_4004), .C(n_4084), .D(n_1923), .Z
		(n_182498556));
	notech_and4 i_85177074(.A(n_4002), .B(n_4076), .C(n_2377), .D(n_4064), .Z
		(n_183098561));
	notech_and4 i_85277073(.A(n_1970), .B(n_1526), .C(n_530), .D(n_2058), .Z
		(n_183598565));
	notech_ao3 i_84377082(.A(n_2216), .B(n_455), .C(n_1987), .Z(n_183898567)
		);
	notech_and4 i_85877067(.A(n_183598565), .B(n_1603), .C(n_3975), .D(n_183898567
		), .Z(n_184198569));
	notech_and4 i_86177064(.A(n_4017), .B(n_183098561), .C(n_184198569), .D(n_2380
		), .Z(n_184298570));
	notech_nand3 i_86377062(.A(n_182498556), .B(n_176698511), .C(n_184298570
		), .Z(n_184398571));
	notech_ao4 i_84577080(.A(n_3957), .B(n_3954), .C(n_3963), .D(n_2517), .Z
		(n_184598573));
	notech_and4 i_85577070(.A(n_3993), .B(n_493), .C(n_3973), .D(n_4085), .Z
		(n_184998577));
	notech_and4 i_85977066(.A(n_1306), .B(n_184598573), .C(n_184998577), .D(n_1340
		), .Z(n_185098578));
	notech_and3 i_76677814(.A(n_2141), .B(n_4013), .C(n_2484), .Z(n_185398581
		));
	notech_and4 i_86977056(.A(n_3374), .B(n_3880), .C(n_4079), .D(n_3981), .Z
		(n_185598583));
	notech_and4 i_87077055(.A(n_4046), .B(n_4053), .C(n_2171), .D(n_4058), .Z
		(n_185998586));
	notech_and4 i_87877047(.A(n_4084), .B(n_2394), .C(n_520), .D(n_3982), .Z
		(n_186498591));
	notech_and4 i_88377043(.A(n_444), .B(n_4046), .C(n_186498591), .D(n_185398581
		), .Z(n_186798593));
	notech_and4 i_87977046(.A(n_2024), .B(n_2047), .C(n_1780), .D(n_201498717
		), .Z(n_187298596));
	notech_and4 i_89677030(.A(n_1346), .B(n_204), .C(n_1284), .D(n_215), .Z(n_187798601
		));
	notech_and4 i_89777029(.A(n_2171), .B(n_530), .C(n_218), .D(n_254), .Z(n_188098604
		));
	notech_and4 i_89877028(.A(n_3975), .B(n_4085), .C(n_34072), .D(n_1615), 
		.Z(n_188598609));
	notech_ao3 i_89577031(.A(n_1130), .B(n_34050), .C(n_122398057), .Z(n_188998613
		));
	notech_and3 i_89977027(.A(n_69852396), .B(n_4004), .C(n_188998613), .Z(n_189098614
		));
	notech_and4 i_90477022(.A(n_189098614), .B(n_185398581), .C(n_2434), .D(n_188598609
		), .Z(n_189298616));
	notech_nao3 i_90677020(.A(n_1919), .B(n_34071), .C(n_2164), .Z(n_189498618
		));
	notech_or4 i_90977017(.A(n_34051), .B(n_189498618), .C(n_34069), .D(n_34131
		), .Z(n_189698620));
	notech_or4 i_14877862(.A(n_4011), .B(n_1640), .C(n_4009), .D(n_189698620
		), .Z(n_189798621));
	notech_or4 i_15877860(.A(n_124098073), .B(n_34132), .C(\udeco[5] ), .D(n_189698620
		), .Z(n_190098623));
	notech_nand3 i_10397771(.A(n_3779), .B(n_1865), .C(n_194998666), .Z(n_190898630
		));
	notech_and4 i_10297772(.A(n_2352), .B(n_2654), .C(n_1856), .D(n_2344), .Z
		(n_190998631));
	notech_or4 i_118397774(.A(n_59558), .B(n_3935), .C(n_59576), .D(n_59585)
		, .Z(n_191198633));
	notech_nand2 i_114097776(.A(modrm[3]), .B(n_34137), .Z(n_191398635));
	notech_and2 i_113797777(.A(n_3763), .B(n_34055), .Z(n_191498636));
	notech_and2 i_113997778(.A(modrm[0]), .B(n_190898630), .Z(n_191598637)
		);
	notech_or4 i_92997779(.A(n_1321), .B(n_191498636), .C(n_191598637), .D(n_34147
		), .Z(\udeco[124] ));
	notech_and3 i_33697781(.A(n_2302), .B(n_34152), .C(n_34053), .Z(n_191798639
		));
	notech_or4 i_116497782(.A(n_2348), .B(n_59502), .C(n_59425), .D(n_191798639
		), .Z(n_191898640));
	notech_nao3 i_116397783(.A(n_34009), .B(n_34006), .C(n_2318), .Z(n_191998641
		));
	notech_and4 i_89297784(.A(n_199898701), .B(n_199498698), .C(n_2694), .D(n_1942
		), .Z(udeco_119101158));
	notech_nand3 i_14897785(.A(n_3736), .B(n_2099), .C(n_1905), .Z(n_192198642
		));
	notech_or4 i_141097787(.A(n_59558), .B(n_2316), .C(n_2389), .D(n_3761), 
		.Z(n_192698644));
	notech_nand2 i_141297788(.A(modrm[0]), .B(n_192198642), .Z(n_192798645)
		);
	notech_and2 i_140997789(.A(modrm[3]), .B(n_3773), .Z(n_192998646));
	notech_and2 i_141197790(.A(n_34056), .B(n_34119), .Z(n_193098647));
	notech_or4 i_85097791(.A(n_1321), .B(n_192998646), .C(n_34155), .D(n_193098647
		), .Z(\udeco[116] ));
	notech_or4 i_144397792(.A(n_59416), .B(n_2373), .C(n_59443), .D(n_2401),
		 .Z(n_193198648));
	notech_and4 i_84297793(.A(n_204598743), .B(n_201798719), .C(n_2684), .D(n_2890
		), .Z(udeco_114101157));
	notech_and4 i_82097794(.A(n_2704), .B(n_2684), .C(n_207798769), .D(n_2890
		), .Z(udeco_113101156));
	notech_or4 i_168297795(.A(n_59416), .B(n_2373), .C(n_3845), .D(n_59479),
		 .Z(n_193298649));
	notech_or4 i_168697796(.A(n_59558), .B(n_2313), .C(n_59493), .D(n_2348),
		 .Z(n_193398650));
	notech_and2 i_168597797(.A(opz[0]), .B(n_34059), .Z(n_193498651));
	notech_or4 i_66297798(.A(n_193498651), .B(n_209298783), .C(n_34164), .D(n_34161
		), .Z(\udeco[104] ));
	notech_and2 i_12697799(.A(n_3992), .B(n_3876), .Z(n_5254));
	notech_nao3 i_62897803(.A(n_211498802), .B(n_5254), .C(n_210198790), .Z(\udeco[49] 
		));
	notech_or4 i_172397804(.A(n_59416), .B(n_2037), .C(n_4072), .D(n_59479),
		 .Z(n_193898655));
	notech_and4 i_58297805(.A(n_193898655), .B(n_213898823), .C(n_1593), .D(n_894
		), .Z(udeco_37101155));
	notech_nao3 i_175097808(.A(n_34009), .B(n_34144), .C(n_2499), .Z(n_194198658
		));
	notech_or2 i_174797809(.A(n_2124), .B(n_59621), .Z(n_194298659));
	notech_or4 i_174997810(.A(n_59416), .B(n_2315), .C(n_59443), .D(n_3836),
		 .Z(n_194398660));
	notech_nao3 i_56110291(.A(n_216898847), .B(n_214398828), .C(n_1326), .Z(\udeco[34] 
		));
	notech_or2 i_182697811(.A(n_2151), .B(n_59470), .Z(n_194498661));
	notech_or2 i_182897812(.A(n_3697), .B(n_59621), .Z(n_194598662));
	notech_or2 i_182797813(.A(n_3728), .B(n_59443), .Z(n_194698663));
	notech_nao3 i_49497814(.A(n_717), .B(n_219698872), .C(n_1326), .Z(\udeco[26] 
		));
	notech_and4 i_47210313(.A(n_520), .B(n_537), .C(n_2567), .D(n_221598889)
		, .Z(udeco_23101154));
	notech_nao3 i_34697815(.A(n_1951), .B(n_2380), .C(n_4057), .Z(n_1326));
	notech_or4 i_17297817(.A(n_1326), .B(n_34169), .C(n_34052), .D(n_3978), 
		.Z(n_1321));
	notech_ao3 i_113197819(.A(n_3777), .B(n_3987), .C(n_3846), .Z(n_194998666
		));
	notech_ao4 i_114297823(.A(n_59527), .B(n_4070), .C(n_2348), .D(n_2338), 
		.Z(n_195698670));
	notech_ao4 i_114397824(.A(n_2166), .B(n_3760), .C(n_34136), .D(n_3935), 
		.Z(n_195798671));
	notech_and4 i_114697827(.A(n_195798671), .B(n_195698670), .C(n_3834), .D
		(n_247296910), .Z(n_196298674));
	notech_and4 i_114997830(.A(n_2450), .B(n_196298674), .C(n_1834), .D(n_191398635
		), .Z(n_196598677));
	notech_and3 i_116697834(.A(n_2676), .B(n_191998641), .C(n_191898640), .Z
		(n_197398681));
	notech_nand2 i_14397836(.A(n_2629), .B(n_34074), .Z(n_1249));
	notech_nand2 i_22197838(.A(n_34187), .B(n_34077), .Z(n_1180));
	notech_and4 i_26697841(.A(n_2216), .B(n_2709), .C(n_2151), .D(n_34143), 
		.Z(n_1130));
	notech_and4 i_133197842(.A(n_2231), .B(n_1833), .C(n_2188), .D(n_1907), 
		.Z(n_197798685));
	notech_and4 i_133397845(.A(n_2630), .B(n_3733), .C(n_3993), .D(n_197798685
		), .Z(n_198198688));
	notech_and4 i_133697848(.A(n_198198688), .B(n_2638), .C(n_1130), .D(n_2065
		), .Z(n_198598691));
	notech_and3 i_133897850(.A(n_4002), .B(n_2166), .C(n_2829), .Z(n_198898693
		));
	notech_and4 i_134097852(.A(n_2827), .B(n_198598691), .C(n_198898693), .D
		(n_2414), .Z(n_199098695));
	notech_and4 i_134697855(.A(n_2826), .B(n_199098695), .C(n_2707), .D(n_1920
		), .Z(n_199498698));
	notech_and4 i_134597858(.A(n_2522), .B(n_2831), .C(n_2510), .D(n_2605), 
		.Z(n_199898701));
	notech_and2 i_61097861(.A(n_4029), .B(n_3967), .Z(n_200298705));
	notech_ao4 i_141397862(.A(n_1984), .B(n_59527), .C(n_2383), .D(n_2865), 
		.Z(n_200398706));
	notech_and4 i_141697865(.A(n_200398706), .B(n_2857), .C(n_192698644), .D
		(n_34057), .Z(n_200698709));
	notech_and4 i_141897867(.A(n_2479), .B(n_200698709), .C(n_34075), .D(n_34148
		), .Z(n_200898711));
	notech_and4 i_142197870(.A(n_200298705), .B(n_200898711), .C(n_2884), .D
		(n_192798645), .Z(n_201198714));
	notech_and2 i_61297873(.A(n_1993), .B(n_4040), .Z(n_201498717));
	notech_and4 i_146697875(.A(n_1993), .B(n_4040), .C(n_2309), .D(n_2483), 
		.Z(n_201798719));
	notech_and4 i_25797877(.A(n_1886), .B(n_2686), .C(n_2572), .D(n_2899), .Z
		(n_202098721));
	notech_and4 i_71097882(.A(n_4007), .B(n_3672), .C(n_1537), .D(n_193198648
		), .Z(n_202798726));
	notech_and4 i_144897885(.A(n_2629), .B(n_3964), .C(n_2709), .D(n_34060),
		 .Z(n_203198729));
	notech_and4 i_145197888(.A(n_2765), .B(n_3867), .C(n_203198729), .D(n_2124
		), .Z(n_203498732));
	notech_and3 i_145397890(.A(n_1949), .B(n_1796), .C(n_3880), .Z(n_203698734
		));
	notech_and4 i_145697892(.A(n_3777), .B(n_203498732), .C(n_1526), .D(n_203698734
		), .Z(n_203898736));
	notech_and4 i_145997895(.A(n_203898736), .B(n_198898693), .C(n_2655), .D
		(n_202798726), .Z(n_204198739));
	notech_and4 i_146597898(.A(n_2903), .B(n_2605), .C(n_204198739), .D(n_1504
		), .Z(n_204498742));
	notech_and4 i_146797899(.A(n_2898), .B(n_202098721), .C(n_2893), .D(n_204498742
		), .Z(n_204598743));
	notech_and4 i_148697905(.A(n_3994), .B(n_2839), .C(n_202798726), .D(n_2852
		), .Z(n_205498749));
	notech_ao3 i_147297908(.A(n_2516), .B(n_34058), .C(n_4010), .Z(n_205798752
		));
	notech_and4 i_147597911(.A(n_2765), .B(n_3931), .C(n_3751), .D(n_205798752
		), .Z(n_206198755));
	notech_and4 i_147897914(.A(n_2625), .B(n_2176), .C(n_206198755), .D(n_2591
		), .Z(n_206498758));
	notech_and4 i_148297917(.A(n_2332), .B(n_206498758), .C(n_2534), .D(n_2539
		), .Z(n_206898761));
	notech_and4 i_148797919(.A(n_2572), .B(n_1969), .C(n_206898761), .D(n_2656
		), .Z(n_207098763));
	notech_and4 i_149097922(.A(n_2722), .B(n_2898), .C(n_207098763), .D(n_2850
		), .Z(n_207398766));
	notech_and4 i_149297923(.A(n_4040), .B(n_205498749), .C(n_207398766), .D
		(n_1993), .Z(n_207498767));
	notech_and4 i_149497925(.A(n_2834), .B(n_2893), .C(n_207498767), .D(n_2688
		), .Z(n_207798769));
	notech_and2 i_72097928(.A(n_3973), .B(n_4029), .Z(n_843));
	notech_and4 i_26497931(.A(n_2327), .B(n_193298649), .C(n_3665), .D(n_34207
		), .Z(n_208398774));
	notech_and4 i_168997934(.A(n_3998), .B(n_193398650), .C(n_3890), .D(n_34060
		), .Z(n_208698777));
	notech_and4 i_169297937(.A(n_208698777), .B(n_1290), .C(n_2162), .D(n_2380
		), .Z(n_208998780));
	notech_or4 i_169597940(.A(n_3820), .B(n_34061), .C(n_1249), .D(n_34162),
		 .Z(n_209298783));
	notech_nand3 i_4353(.A(n_223496909), .B(n_1792), .C(n_1999), .Z(n_209698786
		));
	notech_and4 i_4356(.A(n_34063), .B(n_4019), .C(n_34064), .D(n_1972), .Z(n_210098789
		));
	notech_or4 i_37397945(.A(n_34181), .B(n_34165), .C(n_34167), .D(n_1180),
		 .Z(n_210198790));
	notech_and2 i_4347(.A(n_4026), .B(n_3982), .Z(n_69852396));
	notech_and2 i_4298(.A(n_3838), .B(n_3987), .Z(n_210398792));
	notech_ao4 i_65097947(.A(n_2113), .B(n_2373), .C(n_2278), .D(n_2346), .Z
		(n_210498793));
	notech_ao4 i_170697948(.A(n_2275), .B(n_2118), .C(n_2564), .D(n_59461), 
		.Z(n_210598794));
	notech_and4 i_170997951(.A(n_210598794), .B(n_210498793), .C(n_4031), .D
		(n_1816), .Z(n_210898797));
	notech_and4 i_171397954(.A(n_2340), .B(n_210898797), .C(n_2099), .D(n_210398792
		), .Z(n_211198800));
	notech_and4 i_171597956(.A(n_4032), .B(n_4030), .C(n_211198800), .D(n_69852396
		), .Z(n_211498802));
	notech_and4 i_80797958(.A(n_4076), .B(n_193898655), .C(n_2615), .D(n_2091
		), .Z(n_211798804));
	notech_ao3 i_4572(.A(n_4014), .B(n_1329), .C(n_34012), .Z(n_212098806)
		);
	notech_and4 i_173897961(.A(n_872), .B(n_2500), .C(n_212098806), .D(n_200298705
		), .Z(n_212298808));
	notech_and2 i_74297962(.A(n_3994), .B(n_4085), .Z(n_692));
	notech_and3 i_4510(.A(n_2629), .B(n_4086), .C(n_34074), .Z(n_212498809)
		);
	notech_and4 i_172697966(.A(n_3973), .B(n_3736), .C(n_4031), .D(n_1114), 
		.Z(n_212898813));
	notech_and4 i_172997969(.A(n_212898813), .B(n_2743), .C(n_3061), .D(n_34065
		), .Z(n_213198816));
	notech_and4 i_173397972(.A(n_4034), .B(n_213198816), .C(n_2465), .D(n_861
		), .Z(n_213498819));
	notech_and4 i_173797974(.A(n_2036), .B(n_1014), .C(n_213498819), .D(n_34189
		), .Z(n_213698821));
	notech_and4 i_174097976(.A(n_3994), .B(n_213698821), .C(n_212298808), .D
		(n_4085), .Z(n_213898823));
	notech_and4 i_4614(.A(n_2192), .B(n_4017), .C(n_2500), .D(n_3981), .Z(n_214098825
		));
	notech_and4 i_4656(.A(n_2663), .B(n_2327), .C(n_214098825), .D(n_34148),
		 .Z(n_214398828));
	notech_ao3 i_4531(.A(n_4041), .B(n_1896), .C(n_222398896), .Z(n_214598830
		));
	notech_nand2 i_351097983(.A(n_34077), .B(n_34073), .Z(n_214998833));
	notech_ao4 i_175197984(.A(n_59470), .B(n_34143), .C(n_59443), .D(n_34185
		), .Z(n_215098834));
	notech_and4 i_175497987(.A(n_215098834), .B(n_3992), .C(n_194198658), .D
		(n_34180), .Z(n_215498837));
	notech_and4 i_175997990(.A(n_215498837), .B(n_194298659), .C(n_2017), .D
		(n_194398660), .Z(n_215898840));
	notech_and4 i_176097991(.A(n_811), .B(n_2340), .C(n_214598830), .D(n_215898840
		), .Z(n_215998841));
	notech_and4 i_176397993(.A(n_4055), .B(n_2538), .C(n_843), .D(n_215998841
		), .Z(n_216198843));
	notech_and4 i_176497994(.A(n_2099), .B(n_216198843), .C(n_3736), .D(n_2116
		), .Z(n_216298844));
	notech_and4 i_176797997(.A(n_960), .B(n_894), .C(n_2903), .D(n_216298844
		), .Z(n_216898847));
	notech_and3 i_184498000(.A(n_3102), .B(n_738), .C(n_2588), .Z(n_217298850
		));
	notech_and4 i_184898002(.A(n_34148), .B(n_217298850), .C(n_3098), .D(n_34044
		), .Z(n_217498852));
	notech_and4 i_183198006(.A(n_4026), .B(n_4041), .C(n_4013), .D(n_3980), 
		.Z(n_217998856));
	notech_and3 i_183498008(.A(n_217998856), .B(n_2305), .C(n_34070), .Z(n_218198858
		));
	notech_and4 i_183898010(.A(n_1290), .B(n_194498661), .C(n_218198858), .D
		(n_194598662), .Z(n_218498860));
	notech_and4 i_183998014(.A(n_3103), .B(n_853), .C(n_2099), .D(n_2533), .Z
		(n_218898864));
	notech_and4 i_184398016(.A(n_218898864), .B(n_2465), .C(n_218498860), .D
		(n_2015), .Z(n_219098866));
	notech_and4 i_184998019(.A(n_219098866), .B(n_222898901), .C(n_34071), .D
		(n_194698663), .Z(n_219398869));
	notech_and4 i_185298022(.A(n_703), .B(n_2246), .C(n_219398869), .D(n_217498852
		), .Z(n_219698872));
	notech_and4 i_195598026(.A(n_3049), .B(n_2723), .C(n_2928), .D(n_2024), 
		.Z(n_220098876));
	notech_and3 i_194798029(.A(n_4048), .B(n_4047), .C(n_4019), .Z(n_220398879
		));
	notech_and4 i_195098032(.A(n_2365), .B(n_3739), .C(n_4049), .D(n_220398879
		), .Z(n_220698882));
	notech_and4 i_195698035(.A(n_2212), .B(n_2522), .C(n_200298705), .D(n_220698882
		), .Z(n_220998885));
	notech_and4 i_195998037(.A(n_2157), .B(n_220998885), .C(n_3177), .D(n_220098876
		), .Z(n_221198887));
	notech_and4 i_196198039(.A(n_1993), .B(n_4040), .C(n_221198887), .D(n_530
		), .Z(n_221598889));
	notech_nand3 i_20077883(.A(n_2123), .B(n_4034), .C(n_4022), .Z(n_221898892
		));
	notech_and2 i_413977873(.A(n_34046), .B(n_4062), .Z(n_2219));
	notech_and3 i_4288(.A(n_3992), .B(n_3876), .C(n_2377), .Z(n_222198894)
		);
	notech_and3 i_61777832(.A(n_4067), .B(n_4022), .C(n_34064), .Z(n_222298895
		));
	notech_and4 i_177805(.A(n_2344), .B(n_3279), .C(n_3545), .D(n_1856), .Z(n_1607
		));
	notech_ao3 i_16198042(.A(n_34206), .B(n_3895), .C(n_2348), .Z(n_222398896
		));
	notech_or2 i_3625(.A(n_4089), .B(n_4024), .Z(n_222498897));
	notech_nand3 i_3834(.A(n_2073), .B(n_2202), .C(n_4082), .Z(n_222598898)
		);
	notech_ao4 i_4638(.A(n_2303), .B(n_34151), .C(n_34140), .D(n_2291), .Z(n_222698899
		));
	notech_nand2 i_4677760(.A(modrm[4]), .B(n_34226), .Z(n_1606));
	notech_ao4 i_41798043(.A(n_4072), .B(n_34138), .C(n_34142), .D(n_4090), 
		.Z(n_222798900));
	notech_ao4 i_55998044(.A(n_3954), .B(n_3957), .C(n_2339), .D(n_2299), .Z
		(n_222898901));
	notech_nand3 i_69598045(.A(n_2587), .B(n_197398681), .C(n_2722), .Z(n_222998902
		));
	notech_nand3 i_79798046(.A(n_4086), .B(n_4044), .C(n_34148), .Z(n_223098903
		));
	notech_nand2 i_4177765(.A(n_2390), .B(n_1791), .Z(n_1604));
	notech_inv i_35777(.A(n_1614), .Z(\udeco[125] ));
	notech_inv i_35778(.A(n_1620), .Z(\udeco[123] ));
	notech_inv i_35779(.A(n_1628), .Z(\udeco[45] ));
	notech_inv i_35780(.A(n_1802), .Z(n_34004));
	notech_inv i_35781(.A(n_1639), .Z(\udeco[27] ));
	notech_inv i_35782(.A(n_2027), .Z(n_34006));
	notech_inv i_35783(.A(n_2359), .Z(n_34007));
	notech_inv i_35784(.A(n_2469), .Z(n_34008));
	notech_inv i_35785(.A(n_2149), .Z(n_34009));
	notech_inv i_35786(.A(n_59461), .Z(n_34010));
	notech_inv i_35787(.A(n_2059), .Z(n_34011));
	notech_inv i_35788(.A(n_2005), .Z(n_34012));
	notech_inv i_35789(.A(n_2098), .Z(n_34013));
	notech_inv i_35790(.A(n_2202), .Z(n_34014));
	notech_inv i_35791(.A(n_2078), .Z(n_34015));
	notech_inv i_35792(.A(n_2013), .Z(n_34016));
	notech_inv i_35793(.A(n_2020), .Z(\udeco[112] ));
	notech_inv i_35794(.A(n_2055), .Z(\udeco[109] ));
	notech_inv i_35795(.A(n_2092), .Z(\udeco[32] ));
	notech_inv i_35796(.A(n_2127), .Z(\udeco[24] ));
	notech_inv i_35797(.A(n_2135), .Z(\udeco[20] ));
	notech_inv i_35798(.A(n_2146), .Z(\udeco[18] ));
	notech_inv i_35799(.A(n_2177), .Z(\udeco[17] ));
	notech_inv i_35800(.A(n_2208), .Z(\udeco[13] ));
	notech_inv i_35801(.A(n_221996908), .Z(\udeco[11] ));
	notech_inv i_35802(.A(n_2227), .Z(\udeco[10] ));
	notech_inv i_35803(.A(n_2241), .Z(\udeco[9] ));
	notech_inv i_35804(.A(n_2270), .Z(\udeco[0] ));
	notech_inv i_35805(.A(n_4003), .Z(n_34029));
	notech_inv i_35806(.A(n_4080), .Z(n_34030));
	notech_inv i_35807(.A(n_3974), .Z(n_34031));
	notech_inv i_35808(.A(n_207953599), .Z(n_34032));
	notech_inv i_35809(.A(n_4018), .Z(n_34033));
	notech_inv i_35810(.A(n_4093), .Z(n_34034));
	notech_inv i_35811(.A(n_4062), .Z(n_34035));
	notech_inv i_35812(.A(n_4057), .Z(n_34036));
	notech_inv i_35813(.A(n_4052), .Z(n_34037));
	notech_inv i_35814(.A(n_4091), .Z(n_34038));
	notech_inv i_35815(.A(n_4054), .Z(n_34039));
	notech_inv i_35816(.A(n_4050), .Z(n_34040));
	notech_inv i_35817(.A(n_4065), .Z(n_34041));
	notech_inv i_35818(.A(n_3969), .Z(n_34042));
	notech_inv i_35819(.A(n_4060), .Z(n_34043));
	notech_inv i_35820(.A(n_4015), .Z(n_34044));
	notech_inv i_35821(.A(n_4059), .Z(n_34045));
	notech_inv i_35822(.A(n_4045), .Z(n_34046));
	notech_inv i_35823(.A(n_3971), .Z(n_34047));
	notech_inv i_35824(.A(n_3981), .Z(n_34048));
	notech_inv i_35825(.A(n_204853574), .Z(n_34049));
	notech_inv i_35826(.A(n_4033), .Z(n_34050));
	notech_inv i_35827(.A(n_3984), .Z(n_34051));
	notech_inv i_35828(.A(n_4082), .Z(n_34052));
	notech_inv i_35829(.A(n_3908), .Z(n_34053));
	notech_inv i_35830(.A(n_3846), .Z(n_34054));
	notech_inv i_35831(.A(n_4071), .Z(n_34055));
	notech_inv i_35832(.A(n_3760), .Z(n_34056));
	notech_inv i_35833(.A(n_4006), .Z(n_34057));
	notech_inv i_35834(.A(n_4011), .Z(n_34058));
	notech_inv i_35835(.A(n_3955), .Z(n_34059));
	notech_inv i_35836(.A(n_4009), .Z(n_34060));
	notech_inv i_35837(.A(n_3972), .Z(n_34061));
	notech_inv i_35838(.A(n_3820), .Z(n_34062));
	notech_inv i_35839(.A(n_3990), .Z(n_34063));
	notech_inv i_35840(.A(n_4023), .Z(n_34064));
	notech_inv i_35841(.A(n_4035), .Z(n_34065));
	notech_inv i_35842(.A(n_3728), .Z(n_34066));
	notech_inv i_35843(.A(n_3697), .Z(n_34067));
	notech_inv i_35844(.A(n_3980), .Z(n_34068));
	notech_inv i_35845(.A(n_2305), .Z(n_34069));
	notech_inv i_35846(.A(n_4001), .Z(n_34070));
	notech_inv i_35847(.A(n_3986), .Z(n_34071));
	notech_inv i_35848(.A(n_4088), .Z(n_34072));
	notech_inv i_35849(.A(n_3978), .Z(n_34073));
	notech_inv i_35850(.A(n_3950), .Z(n_34074));
	notech_inv i_35851(.A(n_3985), .Z(n_34075));
	notech_inv i_35852(.A(n_4089), .Z(n_34076));
	notech_inv i_35853(.A(n_3968), .Z(n_34077));
	notech_inv i_35854(.A(n_4085), .Z(n_34078));
	notech_inv i_35855(.A(n_2102), .Z(n_34079));
	notech_inv i_35856(.A(n_2354), .Z(n_34080));
	notech_inv i_35857(.A(n_1708), .Z(n_34081));
	notech_inv i_35858(.A(n_1709), .Z(n_34082));
	notech_inv i_35859(.A(n_122898062), .Z(n_34083));
	notech_inv i_35860(.A(n_125898089), .Z(n_34084));
	notech_inv i_35861(.A(n_126998096), .Z(n_34085));
	notech_inv i_35862(.A(n_1712), .Z(n_34086));
	notech_inv i_35863(.A(n_1870), .Z(n_34087));
	notech_inv i_35864(.A(n_127698103), .Z(n_34088));
	notech_inv i_35865(.A(n_2397), .Z(n_34089));
	notech_inv i_35866(.A(n_133498147), .Z(n_34090));
	notech_inv i_35867(.A(n_136898174), .Z(n_34091));
	notech_inv i_35868(.A(n_138998191), .Z(n_34092));
	notech_inv i_35869(.A(n_1953), .Z(n_34093));
	notech_inv i_35870(.A(n_121198045), .Z(n_34094));
	notech_inv i_35871(.A(n_143898235), .Z(n_34095));
	notech_inv i_35872(.A(n_146998263), .Z(n_34096));
	notech_inv i_35873(.A(n_2614), .Z(n_34097));
	notech_inv i_35874(.A(n_2878), .Z(n_34098));
	notech_inv i_35875(.A(n_1978), .Z(n_34099));
	notech_inv i_35876(.A(n_2854), .Z(n_34100));
	notech_inv i_35877(.A(n_1623), .Z(n_34101));
	notech_inv i_35878(.A(n_153498319), .Z(n_34102));
	notech_inv i_35879(.A(n_2304), .Z(n_34103));
	notech_inv i_35880(.A(n_155198331), .Z(n_34104));
	notech_inv i_35881(.A(n_1981), .Z(n_34105));
	notech_inv i_35882(.A(n_1933), .Z(n_34106));
	notech_inv i_35883(.A(n_1704), .Z(n_34107));
	notech_inv i_35884(.A(n_1951), .Z(n_34108));
	notech_inv i_35885(.A(n_162298390), .Z(n_34109));
	notech_inv i_35886(.A(n_2759), .Z(n_34110));
	notech_inv i_35887(.A(n_2754), .Z(n_34111));
	notech_inv i_35888(.A(n_1702), .Z(n_34112));
	notech_inv i_35889(.A(n_3107), .Z(n_34113));
	notech_inv i_35890(.A(n_2713), .Z(n_34114));
	notech_inv i_35891(.A(n_172198473), .Z(n_34115));
	notech_inv i_35892(.A(n_172498476), .Z(n_34116));
	notech_inv i_35893(.A(n_2678), .Z(n_34117));
	notech_inv i_35894(.A(n_3510), .Z(n_34118));
	notech_inv i_35895(.A(n_1718), .Z(n_34119));
	notech_inv i_35896(.A(n_1699), .Z(n_34120));
	notech_inv i_35897(.A(n_1263), .Z(n_34121));
	notech_inv i_35898(.A(n_2620), .Z(n_34122));
	notech_inv i_35899(.A(n_2615), .Z(n_34123));
	notech_inv i_35900(.A(n_185098578), .Z(n_34124));
	notech_inv i_35901(.A(n_696), .Z(n_34125));
	notech_inv i_35902(.A(n_2543), .Z(n_34126));
	notech_inv i_35903(.A(n_2541), .Z(n_34127));
	notech_inv i_35904(.A(n_2536), .Z(n_34128));
	notech_inv i_35905(.A(n_1615), .Z(n_34129));
	notech_inv i_35906(.A(n_2296), .Z(n_34130));
	notech_inv i_35907(.A(n_1923), .Z(n_34131));
	notech_inv i_35908(.A(n_2022), .Z(n_34132));
	notech_inv i_35909(.A(n_190098623), .Z(n_34133));
	notech_inv i_35910(.A(n_2426), .Z(n_34134));
	notech_inv i_35911(.A(n_1969), .Z(n_34135));
	notech_inv i_35912(.A(n_2369), .Z(n_34136));
	notech_inv i_35913(.A(n_190998631), .Z(n_34137));
	notech_inv i_35914(.A(n_3959), .Z(n_34138));
	notech_inv i_35915(.A(n_1942), .Z(n_34139));
	notech_inv i_35916(.A(n_2390), .Z(n_34140));
	notech_inv i_35917(.A(n_2401), .Z(n_34141));
	notech_inv i_35918(.A(n_2210), .Z(n_34142));
	notech_inv i_35919(.A(n_1987), .Z(n_34143));
	notech_inv i_35920(.A(n_2355), .Z(n_34144));
	notech_inv i_35921(.A(n_2466), .Z(n_34145));
	notech_inv i_35922(.A(n_2463), .Z(n_34146));
	notech_inv i_35923(.A(n_196598677), .Z(n_34147));
	notech_inv i_35924(.A(n_1249), .Z(n_34148));
	notech_inv i_35925(.A(n_1180), .Z(n_34149));
	notech_inv i_35926(.A(n_2431), .Z(n_34150));
	notech_inv i_35927(.A(n_2418), .Z(n_34151));
	notech_inv i_35928(.A(n_2287), .Z(n_34152));
	notech_inv i_35929(.A(n_1905), .Z(n_34153));
	notech_inv i_35930(.A(n_2391), .Z(n_34154));
	notech_inv i_35931(.A(n_201198714), .Z(n_34155));
	notech_inv i_35932(.A(n_2852), .Z(n_34156));
	notech_inv i_35933(.A(n_2324), .Z(n_34157));
	notech_inv i_35934(.A(n_2321), .Z(n_34158));
	notech_inv i_35935(.A(n_2656), .Z(n_34159));
	notech_inv i_35936(.A(n_2850), .Z(n_34160));
	notech_inv i_35937(.A(n_208398774), .Z(n_34161));
	notech_inv i_35938(.A(n_208998780), .Z(n_34162));
	notech_inv i_35939(.A(n_2186), .Z(n_34163));
	notech_inv i_35940(.A(n_2792), .Z(n_34164));
	notech_inv i_35941(.A(n_1999), .Z(n_34165));
	notech_inv i_35942(.A(n_1972), .Z(n_34166));
	notech_inv i_35943(.A(n_210098789), .Z(n_34167));
	notech_inv i_35944(.A(n_2038), .Z(n_34168));
	notech_inv i_35945(.A(n_1816), .Z(n_34169));
	notech_inv i_35946(.A(n_2006), .Z(n_34170));
	notech_inv i_35947(.A(n_1986), .Z(n_34171));
	notech_inv i_35948(.A(n_1965), .Z(n_34172));
	notech_inv i_35949(.A(n_1624), .Z(n_34173));
	notech_inv i_35950(.A(n_2036), .Z(n_34174));
	notech_inv i_35951(.A(n_1943), .Z(n_34175));
	notech_inv i_35952(.A(n_1114), .Z(n_34176));
	notech_inv i_35953(.A(n_1841), .Z(n_34177));
	notech_inv i_35954(.A(n_1840), .Z(n_34178));
	notech_inv i_35955(.A(n_2116), .Z(n_34179));
	notech_inv i_35956(.A(n_214998833), .Z(n_34180));
	notech_inv i_35957(.A(n_2017), .Z(n_34181));
	notech_inv i_35958(.A(n_960), .Z(n_34182));
	notech_inv i_35959(.A(n_1695), .Z(n_34183));
	notech_inv i_35960(.A(n_2365), .Z(n_34184));
	notech_inv i_35961(.A(n_221898892), .Z(n_34185));
	notech_inv i_35962(.A(n_2357), .Z(n_34186));
	notech_inv i_35963(.A(n_222498897), .Z(n_34187));
	notech_inv i_35964(.A(n_2380), .Z(\udeco[5] ));
	notech_inv i_35965(.A(n_223098903), .Z(n_34189));
	notech_inv i_35966(.A(n_1950), .Z(n_34190));
	notech_inv i_35968(.A(n_59594), .Z(n_34192));
	notech_inv i_35969(.A(n_59580), .Z(n_34193));
	notech_inv i_35971(.A(n_59612), .Z(n_34195));
	notech_inv i_35972(.A(n_59634), .Z(n_34196));
	notech_inv i_35973(.A(op[7]), .Z(n_34197));
	notech_inv i_35974(.A(modrm[0]), .Z(n_34198));
	notech_inv i_35975(.A(modrm[1]), .Z(n_34199));
	notech_inv i_35976(.A(modrm[3]), .Z(n_34200));
	notech_inv i_35977(.A(modrm[4]), .Z(n_34201));
	notech_inv i_35978(.A(n_59479), .Z(n_34202));
	notech_inv i_35979(.A(modrm[6]), .Z(n_34203));
	notech_inv i_35980(.A(ipg_fault), .Z(n_34204));
	notech_inv i_35981(.A(twobyte), .Z(n_34205));
	notech_inv i_35982(.A(adz), .Z(n_34206));
	notech_inv i_35983(.A(n_4024), .Z(n_34207));
	notech_inv i_35984(.A(n_1622), .Z(n_34208));
	notech_inv i_35985(.A(n_1608), .Z(n_34209));
	notech_inv i_35986(.A(\udeco[91] ), .Z(n_34210));
	notech_inv i_35987(.A(udeco_73101168), .Z(\udeco[73] ));
	notech_inv i_35988(.A(udeco_101101167), .Z(\udeco[101] ));
	notech_inv i_35989(.A(udeco_103101166), .Z(\udeco[103] ));
	notech_inv i_35990(.A(udeco_35101165), .Z(\udeco[35] ));
	notech_inv i_35991(.A(udeco_29101164), .Z(\udeco[29] ));
	notech_inv i_35992(.A(udeco_28101163), .Z(\udeco[28] ));
	notech_inv i_35993(.A(udeco_21101162), .Z(\udeco[21] ));
	notech_inv i_35994(.A(udeco_15101161), .Z(\udeco[15] ));
	notech_inv i_35995(.A(udeco_14101160), .Z(\udeco[14] ));
	notech_inv i_35996(.A(udeco_12101159), .Z(\udeco[12] ));
	notech_inv i_35997(.A(udeco_119101158), .Z(\udeco[119] ));
	notech_inv i_35998(.A(udeco_114101157), .Z(\udeco[114] ));
	notech_inv i_35999(.A(udeco_113101156), .Z(\udeco[113] ));
	notech_inv i_36000(.A(udeco_37101155), .Z(\udeco[37] ));
	notech_inv i_36001(.A(udeco_23101154), .Z(\udeco[23] ));
	notech_inv i_36002(.A(n_1607), .Z(n_34226));
endmodule
module deco(clk, rstn, useq_ptr, in128, adz, pc_req, ivect, int_main, iack, ie, pg_fault
		, ipg_fault, cpl, cr0, valid_len, to_vliw, lenpc_out, immediate,
		 to_acu, operand_size, reps, over_seg, valid_op, term, start, ready_vliw
		);

	input clk;
	input rstn;
	output [3:0] useq_ptr;
	input [127:0] in128;
	input adz;
	input pc_req;
	input [7:0] ivect;
	input int_main;
	output iack;
	input ie;
	input pg_fault;
	input ipg_fault;
	input [1:0] cpl;
	input [31:0] cr0;
	input [5:0] valid_len;
	output [127:0] to_vliw;
	output [31:0] lenpc_out;
	output [63:0] immediate;
	output [210:0] to_acu;
	output [2:0] operand_size;
	output [2:0] reps;
	output [5:0] over_seg;
	output valid_op;
	input term;
	output start;
	input ready_vliw;

	wire [210:0] to_acu2;
	wire [2:0] opz2;
	wire [210:0] to_acu1;
	wire [127:0] inst_deco1;
	wire [127:0] inst_deco2;
	wire [2:0] reps2;
	wire [31:0] lenpc2;
	wire [3:0] i_ptr;
	wire [1:0] idx_deco;
	wire [5:0] int_excl;
	wire [7:0] ififo_rvect1;
	wire [4:0] fsm;
	wire [2:0] reps1;
	wire [2:0] opz1;
	wire [31:0] lenpc1;
	wire [210:0] to_acu0;
	wire [127:0] inst_deco;
	wire [2:0] opz0;
	wire [2:0] reps0;
	wire [31:0] lenpc;
	wire [7:0] ififo_rvect2;
	wire [7:0] ififo_rvect3;
	wire [7:0] ififo_rvect4;
	wire [127:0] udeco;
	wire [2:0] opz;
	wire [2:0] displc;
	wire [2:0] imm_sz;
	wire [4:0] pfx_sz;



	notech_inv i_15108(.A(n_63212), .Z(n_63275));
	notech_inv i_15106(.A(n_63212), .Z(n_63273));
	notech_inv i_15103(.A(n_63212), .Z(n_63270));
	notech_inv i_15101(.A(n_63212), .Z(n_63268));
	notech_inv i_15098(.A(n_63212), .Z(n_63265));
	notech_inv i_15096(.A(n_63212), .Z(n_63263));
	notech_inv i_15092(.A(n_63212), .Z(n_63259));
	notech_inv i_15090(.A(n_63212), .Z(n_63257));
	notech_inv i_15087(.A(n_63212), .Z(n_63254));
	notech_inv i_15085(.A(n_63212), .Z(n_63252));
	notech_inv i_15082(.A(n_63212), .Z(n_63249));
	notech_inv i_15080(.A(n_63212), .Z(n_63247));
	notech_inv i_15076(.A(n_63212), .Z(n_63243));
	notech_inv i_15074(.A(n_63212), .Z(n_63241));
	notech_inv i_15071(.A(n_63212), .Z(n_63238));
	notech_inv i_15069(.A(n_63212), .Z(n_63236));
	notech_inv i_15066(.A(n_63212), .Z(n_63233));
	notech_inv i_15064(.A(n_63212), .Z(n_63231));
	notech_inv i_15060(.A(n_63214), .Z(n_63227));
	notech_inv i_15058(.A(n_63214), .Z(n_63225));
	notech_inv i_15055(.A(n_63214), .Z(n_63222));
	notech_inv i_15053(.A(n_63214), .Z(n_63220));
	notech_inv i_15050(.A(n_63214), .Z(n_63217));
	notech_inv i_15048(.A(n_63214), .Z(n_63215));
	notech_inv i_15047(.A(n_63213), .Z(n_63214));
	notech_inv i_15046(.A(n_63212), .Z(n_63213));
	notech_inv i_15045(.A(clk), .Z(n_63212));
	notech_inv i_15043(.A(n_63147), .Z(n_63210));
	notech_inv i_15041(.A(n_63147), .Z(n_63208));
	notech_inv i_15038(.A(n_63147), .Z(n_63205));
	notech_inv i_15036(.A(n_63147), .Z(n_63203));
	notech_inv i_15033(.A(n_63147), .Z(n_63200));
	notech_inv i_15031(.A(n_63147), .Z(n_63198));
	notech_inv i_15027(.A(n_63147), .Z(n_63194));
	notech_inv i_15025(.A(n_63147), .Z(n_63192));
	notech_inv i_15022(.A(n_63147), .Z(n_63189));
	notech_inv i_15020(.A(n_63147), .Z(n_63187));
	notech_inv i_15017(.A(n_63147), .Z(n_63184));
	notech_inv i_15015(.A(n_63147), .Z(n_63182));
	notech_inv i_15011(.A(n_63147), .Z(n_63178));
	notech_inv i_15009(.A(n_63147), .Z(n_63176));
	notech_inv i_15006(.A(n_63147), .Z(n_63173));
	notech_inv i_15004(.A(n_63147), .Z(n_63171));
	notech_inv i_15001(.A(n_63147), .Z(n_63168));
	notech_inv i_14999(.A(n_63147), .Z(n_63166));
	notech_inv i_14995(.A(n_63149), .Z(n_63162));
	notech_inv i_14993(.A(n_63149), .Z(n_63160));
	notech_inv i_14990(.A(n_63149), .Z(n_63157));
	notech_inv i_14988(.A(n_63149), .Z(n_63155));
	notech_inv i_14985(.A(n_63149), .Z(n_63152));
	notech_inv i_14983(.A(n_63149), .Z(n_63150));
	notech_inv i_14982(.A(n_63171), .Z(n_63149));
	notech_inv i_14980(.A(clk), .Z(n_63147));
	notech_inv i_14978(.A(n_63082), .Z(n_63145));
	notech_inv i_14976(.A(n_63082), .Z(n_63143));
	notech_inv i_14973(.A(n_63082), .Z(n_63140));
	notech_inv i_14971(.A(n_63082), .Z(n_63138));
	notech_inv i_14968(.A(n_63082), .Z(n_63135));
	notech_inv i_14966(.A(n_63082), .Z(n_63133));
	notech_inv i_14962(.A(n_63082), .Z(n_63129));
	notech_inv i_14960(.A(n_63082), .Z(n_63127));
	notech_inv i_14957(.A(n_63082), .Z(n_63124));
	notech_inv i_14955(.A(n_63082), .Z(n_63122));
	notech_inv i_14952(.A(n_63082), .Z(n_63119));
	notech_inv i_14950(.A(n_63082), .Z(n_63117));
	notech_inv i_14946(.A(n_63082), .Z(n_63113));
	notech_inv i_14944(.A(n_63082), .Z(n_63111));
	notech_inv i_14941(.A(n_63082), .Z(n_63108));
	notech_inv i_14939(.A(n_63082), .Z(n_63106));
	notech_inv i_14936(.A(n_63082), .Z(n_63103));
	notech_inv i_14934(.A(n_63082), .Z(n_63101));
	notech_inv i_14930(.A(n_63084), .Z(n_63097));
	notech_inv i_14928(.A(n_63084), .Z(n_63095));
	notech_inv i_14925(.A(n_63084), .Z(n_63092));
	notech_inv i_14923(.A(n_63084), .Z(n_63090));
	notech_inv i_14920(.A(n_63084), .Z(n_63087));
	notech_inv i_14918(.A(n_63084), .Z(n_63085));
	notech_inv i_14917(.A(n_63106), .Z(n_63084));
	notech_inv i_14915(.A(clk), .Z(n_63082));
	notech_inv i_14531(.A(n_62614), .Z(n_62678));
	notech_inv i_14529(.A(n_62614), .Z(n_62676));
	notech_inv i_14528(.A(n_62614), .Z(n_62675));
	notech_inv i_14524(.A(n_62614), .Z(n_62671));
	notech_inv i_14523(.A(n_62614), .Z(n_62670));
	notech_inv i_14518(.A(n_62614), .Z(n_62665));
	notech_inv i_14514(.A(n_62614), .Z(n_62661));
	notech_inv i_14512(.A(n_62614), .Z(n_62659));
	notech_inv i_14509(.A(n_62614), .Z(n_62656));
	notech_inv i_14507(.A(n_62614), .Z(n_62654));
	notech_inv i_14504(.A(n_62614), .Z(n_62651));
	notech_inv i_14502(.A(n_62614), .Z(n_62649));
	notech_inv i_14498(.A(n_62614), .Z(n_62645));
	notech_inv i_14496(.A(n_62614), .Z(n_62643));
	notech_inv i_14493(.A(n_62614), .Z(n_62640));
	notech_inv i_14491(.A(n_62614), .Z(n_62638));
	notech_inv i_14488(.A(n_62614), .Z(n_62635));
	notech_inv i_14486(.A(n_62614), .Z(n_62633));
	notech_inv i_14482(.A(n_62616), .Z(n_62629));
	notech_inv i_14480(.A(n_62616), .Z(n_62627));
	notech_inv i_14477(.A(n_62616), .Z(n_62624));
	notech_inv i_14475(.A(n_62616), .Z(n_62622));
	notech_inv i_14472(.A(n_62616), .Z(n_62619));
	notech_inv i_14470(.A(n_62616), .Z(n_62617));
	notech_inv i_14469(.A(n_62615), .Z(n_62616));
	notech_inv i_14468(.A(n_62614), .Z(n_62615));
	notech_inv i_14467(.A(rstn), .Z(n_62614));
	notech_inv i_14465(.A(n_62549), .Z(n_62612));
	notech_inv i_14463(.A(n_62549), .Z(n_62610));
	notech_inv i_14460(.A(n_62549), .Z(n_62607));
	notech_inv i_14458(.A(n_62549), .Z(n_62605));
	notech_inv i_14455(.A(n_62549), .Z(n_62602));
	notech_inv i_14453(.A(n_62549), .Z(n_62600));
	notech_inv i_14449(.A(n_62549), .Z(n_62596));
	notech_inv i_14447(.A(n_62549), .Z(n_62594));
	notech_inv i_14444(.A(n_62549), .Z(n_62591));
	notech_inv i_14442(.A(n_62549), .Z(n_62589));
	notech_inv i_14439(.A(n_62549), .Z(n_62586));
	notech_inv i_14437(.A(n_62549), .Z(n_62584));
	notech_inv i_14433(.A(n_62549), .Z(n_62580));
	notech_inv i_14431(.A(n_62549), .Z(n_62578));
	notech_inv i_14428(.A(n_62549), .Z(n_62575));
	notech_inv i_14426(.A(n_62549), .Z(n_62573));
	notech_inv i_14423(.A(n_62549), .Z(n_62570));
	notech_inv i_14421(.A(n_62549), .Z(n_62568));
	notech_inv i_14417(.A(n_62551), .Z(n_62564));
	notech_inv i_14415(.A(n_62551), .Z(n_62562));
	notech_inv i_14412(.A(n_62551), .Z(n_62559));
	notech_inv i_14410(.A(n_62551), .Z(n_62557));
	notech_inv i_14407(.A(n_62551), .Z(n_62554));
	notech_inv i_14405(.A(n_62551), .Z(n_62552));
	notech_inv i_14404(.A(n_62573), .Z(n_62551));
	notech_inv i_14402(.A(rstn), .Z(n_62549));
	notech_inv i_14400(.A(n_62484), .Z(n_62547));
	notech_inv i_14398(.A(n_62484), .Z(n_62545));
	notech_inv i_14395(.A(n_62484), .Z(n_62542));
	notech_inv i_14393(.A(n_62484), .Z(n_62540));
	notech_inv i_14390(.A(n_62484), .Z(n_62537));
	notech_inv i_14388(.A(n_62484), .Z(n_62535));
	notech_inv i_14384(.A(n_62484), .Z(n_62531));
	notech_inv i_14382(.A(n_62484), .Z(n_62529));
	notech_inv i_14379(.A(n_62484), .Z(n_62526));
	notech_inv i_14377(.A(n_62484), .Z(n_62524));
	notech_inv i_14374(.A(n_62484), .Z(n_62521));
	notech_inv i_14372(.A(n_62484), .Z(n_62519));
	notech_inv i_14368(.A(n_62484), .Z(n_62515));
	notech_inv i_14366(.A(n_62484), .Z(n_62513));
	notech_inv i_14363(.A(n_62484), .Z(n_62510));
	notech_inv i_14361(.A(n_62484), .Z(n_62508));
	notech_inv i_14358(.A(n_62484), .Z(n_62505));
	notech_inv i_14356(.A(n_62484), .Z(n_62503));
	notech_inv i_14352(.A(n_62486), .Z(n_62499));
	notech_inv i_14350(.A(n_62486), .Z(n_62497));
	notech_inv i_14347(.A(n_62486), .Z(n_62494));
	notech_inv i_14345(.A(n_62486), .Z(n_62492));
	notech_inv i_14342(.A(n_62486), .Z(n_62489));
	notech_inv i_14340(.A(n_62486), .Z(n_62487));
	notech_inv i_14339(.A(n_62508), .Z(n_62486));
	notech_inv i_14337(.A(rstn), .Z(n_62484));
	notech_inv i_13932(.A(n_62013), .Z(n_62078));
	notech_inv i_13931(.A(n_62013), .Z(n_62077));
	notech_inv i_13926(.A(n_62013), .Z(n_62072));
	notech_inv i_13921(.A(n_62013), .Z(n_62067));
	notech_inv i_13920(.A(n_62013), .Z(n_62066));
	notech_inv i_13915(.A(n_62013), .Z(n_62061));
	notech_inv i_13910(.A(n_62013), .Z(n_62056));
	notech_inv i_13909(.A(n_62013), .Z(n_62055));
	notech_inv i_13904(.A(n_62013), .Z(n_62050));
	notech_inv i_13898(.A(n_62013), .Z(n_62044));
	notech_inv i_13897(.A(n_62013), .Z(n_62043));
	notech_inv i_13892(.A(n_62013), .Z(n_62038));
	notech_inv i_13887(.A(n_62013), .Z(n_62033));
	notech_inv i_13886(.A(n_62013), .Z(n_62032));
	notech_inv i_13881(.A(n_62013), .Z(n_62027));
	notech_inv i_13876(.A(n_62013), .Z(n_62022));
	notech_inv i_13875(.A(n_62013), .Z(n_62021));
	notech_inv i_13870(.A(n_62013), .Z(n_62016));
	notech_inv i_13867(.A(term), .Z(n_62013));
	notech_inv i_13864(.A(n_61979), .Z(n_62010));
	notech_inv i_13863(.A(n_61979), .Z(n_62009));
	notech_inv i_13858(.A(n_61979), .Z(n_62004));
	notech_inv i_13853(.A(n_61979), .Z(n_61999));
	notech_inv i_13852(.A(n_61979), .Z(n_61998));
	notech_inv i_13847(.A(n_61979), .Z(n_61993));
	notech_inv i_13842(.A(n_61979), .Z(n_61988));
	notech_inv i_13841(.A(n_61979), .Z(n_61987));
	notech_inv i_13836(.A(n_61979), .Z(n_61982));
	notech_inv i_13833(.A(term), .Z(n_61979));
	notech_inv i_12908(.A(n_60931), .Z(n_60949));
	notech_inv i_12906(.A(n_60931), .Z(n_60947));
	notech_inv i_12903(.A(n_60931), .Z(n_60944));
	notech_inv i_12901(.A(n_60931), .Z(n_60942));
	notech_inv i_12898(.A(n_60931), .Z(n_60939));
	notech_inv i_12896(.A(n_60931), .Z(n_60937));
	notech_inv i_12893(.A(n_60931), .Z(n_60934));
	notech_inv i_12891(.A(n_60931), .Z(n_60932));
	notech_inv i_12890(.A(n_2911), .Z(n_60931));
	notech_inv i_12881(.A(n_60920), .Z(n_60921));
	notech_inv i_12880(.A(n_2382), .Z(n_60920));
	notech_inv i_12877(.A(n_60851), .Z(n_60916));
	notech_inv i_12876(.A(n_60851), .Z(n_60915));
	notech_inv i_12871(.A(n_60851), .Z(n_60910));
	notech_inv i_12866(.A(n_60851), .Z(n_60905));
	notech_inv i_12865(.A(n_60851), .Z(n_60904));
	notech_inv i_12860(.A(n_60851), .Z(n_60899));
	notech_inv i_12855(.A(n_60851), .Z(n_60894));
	notech_inv i_12854(.A(n_60851), .Z(n_60893));
	notech_inv i_12849(.A(n_60851), .Z(n_60888));
	notech_inv i_12843(.A(n_60851), .Z(n_60882));
	notech_inv i_12842(.A(n_60851), .Z(n_60881));
	notech_inv i_12837(.A(n_60851), .Z(n_60876));
	notech_inv i_12832(.A(n_60851), .Z(n_60871));
	notech_inv i_12831(.A(n_60851), .Z(n_60870));
	notech_inv i_12826(.A(n_60851), .Z(n_60865));
	notech_inv i_12821(.A(n_60851), .Z(n_60860));
	notech_inv i_12820(.A(n_60851), .Z(n_60859));
	notech_inv i_12815(.A(n_60851), .Z(n_60854));
	notech_inv i_12812(.A(n_44738), .Z(n_60851));
	notech_inv i_12809(.A(n_60817), .Z(n_60848));
	notech_inv i_12808(.A(n_60817), .Z(n_60847));
	notech_inv i_12798(.A(n_60817), .Z(n_60837));
	notech_inv i_12797(.A(n_60817), .Z(n_60836));
	notech_inv i_12792(.A(n_60817), .Z(n_60831));
	notech_inv i_12786(.A(n_60817), .Z(n_60825));
	notech_inv i_12781(.A(n_60817), .Z(n_60820));
	notech_inv i_12778(.A(n_44738), .Z(n_60817));
	notech_inv i_12388(.A(n_60364), .Z(n_60418));
	notech_inv i_12387(.A(n_60364), .Z(n_60417));
	notech_inv i_12383(.A(n_60364), .Z(n_60413));
	notech_inv i_12379(.A(n_60364), .Z(n_60409));
	notech_inv i_12378(.A(n_60364), .Z(n_60408));
	notech_inv i_12374(.A(n_60364), .Z(n_60404));
	notech_inv i_12370(.A(n_60364), .Z(n_60400));
	notech_inv i_12369(.A(n_60364), .Z(n_60399));
	notech_inv i_12365(.A(n_60364), .Z(n_60395));
	notech_inv i_12360(.A(n_60364), .Z(n_60390));
	notech_inv i_12359(.A(n_60364), .Z(n_60389));
	notech_inv i_12355(.A(n_60364), .Z(n_60385));
	notech_inv i_12351(.A(n_60364), .Z(n_60381));
	notech_inv i_12350(.A(n_60364), .Z(n_60380));
	notech_inv i_12346(.A(n_60364), .Z(n_60376));
	notech_inv i_12342(.A(n_60364), .Z(n_60372));
	notech_inv i_12341(.A(n_60364), .Z(n_60371));
	notech_inv i_12337(.A(n_60364), .Z(n_60367));
	notech_inv i_12334(.A(n_5770), .Z(n_60364));
	notech_inv i_12332(.A(n_60336), .Z(n_60362));
	notech_inv i_12331(.A(n_60336), .Z(n_60361));
	notech_inv i_12318(.A(n_60347), .Z(n_60348));
	notech_inv i_12317(.A(n_60346), .Z(n_60347));
	notech_inv i_12316(.A(n_60336), .Z(n_60346));
	notech_inv i_12309(.A(n_60338), .Z(n_60339));
	notech_inv i_12308(.A(n_60337), .Z(n_60338));
	notech_inv i_12307(.A(n_60336), .Z(n_60337));
	notech_inv i_12306(.A(n_5770), .Z(n_60336));
	notech_inv i_12304(.A(n_60245), .Z(n_60333));
	notech_inv i_12302(.A(n_60245), .Z(n_60331));
	notech_inv i_12299(.A(n_60245), .Z(n_60328));
	notech_inv i_12297(.A(n_60245), .Z(n_60326));
	notech_inv i_12293(.A(n_60245), .Z(n_60322));
	notech_inv i_12291(.A(n_60245), .Z(n_60320));
	notech_inv i_12288(.A(n_60245), .Z(n_60317));
	notech_inv i_12286(.A(n_60245), .Z(n_60315));
	notech_inv i_12282(.A(n_60245), .Z(n_60311));
	notech_inv i_12280(.A(n_60245), .Z(n_60309));
	notech_inv i_12277(.A(n_60245), .Z(n_60306));
	notech_inv i_12275(.A(n_60245), .Z(n_60304));
	notech_inv i_12271(.A(n_60245), .Z(n_60300));
	notech_inv i_12269(.A(n_60245), .Z(n_60298));
	notech_inv i_12266(.A(n_60245), .Z(n_60295));
	notech_inv i_12264(.A(n_60245), .Z(n_60293));
	notech_inv i_12259(.A(n_60280), .Z(n_60288));
	notech_inv i_12257(.A(n_60280), .Z(n_60286));
	notech_inv i_12254(.A(n_60280), .Z(n_60283));
	notech_inv i_12252(.A(n_60280), .Z(n_60281));
	notech_inv i_12251(.A(n_60326), .Z(n_60280));
	notech_inv i_12248(.A(n_60280), .Z(n_60277));
	notech_inv i_12246(.A(n_60280), .Z(n_60275));
	notech_inv i_12243(.A(n_60280), .Z(n_60272));
	notech_inv i_12241(.A(n_60280), .Z(n_60270));
	notech_inv i_12237(.A(n_60280), .Z(n_60266));
	notech_inv i_12235(.A(n_60280), .Z(n_60264));
	notech_inv i_12232(.A(n_60280), .Z(n_60261));
	notech_inv i_12230(.A(n_60280), .Z(n_60259));
	notech_inv i_12226(.A(n_60245), .Z(n_60255));
	notech_inv i_12224(.A(n_60245), .Z(n_60253));
	notech_inv i_12221(.A(n_60245), .Z(n_60250));
	notech_inv i_12219(.A(n_60245), .Z(n_60248));
	notech_inv i_12216(.A(n_5769), .Z(n_60245));
	notech_inv i_12214(.A(n_60200), .Z(n_60243));
	notech_inv i_12212(.A(n_60200), .Z(n_60241));
	notech_inv i_12209(.A(n_60200), .Z(n_60238));
	notech_inv i_12207(.A(n_60200), .Z(n_60236));
	notech_inv i_12203(.A(n_60200), .Z(n_60232));
	notech_inv i_12201(.A(n_60200), .Z(n_60230));
	notech_inv i_12198(.A(n_60200), .Z(n_60227));
	notech_inv i_12196(.A(n_60200), .Z(n_60225));
	notech_inv i_12192(.A(n_60200), .Z(n_60221));
	notech_inv i_12190(.A(n_60200), .Z(n_60219));
	notech_inv i_12187(.A(n_60200), .Z(n_60216));
	notech_inv i_12185(.A(n_60200), .Z(n_60214));
	notech_inv i_12180(.A(n_60200), .Z(n_60209));
	notech_inv i_12179(.A(n_60200), .Z(n_60208));
	notech_inv i_12174(.A(n_60200), .Z(n_60203));
	notech_inv i_12171(.A(n_5769), .Z(n_60200));
	notech_inv i_12116(.A(n_60130), .Z(n_60148));
	notech_inv i_12114(.A(n_60130), .Z(n_60146));
	notech_inv i_12111(.A(n_60130), .Z(n_60143));
	notech_inv i_12109(.A(n_60130), .Z(n_60141));
	notech_inv i_12106(.A(n_60130), .Z(n_60138));
	notech_inv i_12104(.A(n_60130), .Z(n_60136));
	notech_inv i_12101(.A(n_60130), .Z(n_60133));
	notech_inv i_12099(.A(n_60130), .Z(n_60131));
	notech_inv i_12098(.A(n_3301), .Z(n_60130));
	notech_inv i_12096(.A(n_60109), .Z(n_60127));
	notech_inv i_12094(.A(n_60109), .Z(n_60125));
	notech_inv i_12091(.A(n_60109), .Z(n_60122));
	notech_inv i_12089(.A(n_60109), .Z(n_60120));
	notech_inv i_12086(.A(n_60109), .Z(n_60117));
	notech_inv i_12084(.A(n_60109), .Z(n_60115));
	notech_inv i_12081(.A(n_60109), .Z(n_60112));
	notech_inv i_12079(.A(n_60109), .Z(n_60110));
	notech_inv i_12078(.A(n_5768), .Z(n_60109));
	notech_inv i_11505(.A(n_59487), .Z(n_59489));
	notech_inv i_11504(.A(n_59487), .Z(n_59488));
	notech_inv i_11503(.A(in128[10]), .Z(n_59487));
	notech_inv i_11435(.A(n_1913), .Z(n_59410));
	notech_inv i_11430(.A(n_1913), .Z(n_59405));
	notech_inv i_11426(.A(n_59335), .Z(n_59400));
	notech_inv i_11425(.A(n_59335), .Z(n_59399));
	notech_inv i_11420(.A(n_59335), .Z(n_59394));
	notech_inv i_11415(.A(n_59335), .Z(n_59389));
	notech_inv i_11414(.A(n_59335), .Z(n_59388));
	notech_inv i_11409(.A(n_59335), .Z(n_59383));
	notech_inv i_11404(.A(n_59335), .Z(n_59378));
	notech_inv i_11403(.A(n_59335), .Z(n_59377));
	notech_inv i_11398(.A(n_59335), .Z(n_59372));
	notech_inv i_11392(.A(n_59335), .Z(n_59366));
	notech_inv i_11391(.A(n_59335), .Z(n_59365));
	notech_inv i_11386(.A(n_59335), .Z(n_59360));
	notech_inv i_11381(.A(n_59335), .Z(n_59355));
	notech_inv i_11380(.A(n_59335), .Z(n_59354));
	notech_inv i_11375(.A(n_59335), .Z(n_59349));
	notech_inv i_11370(.A(n_59335), .Z(n_59344));
	notech_inv i_11369(.A(n_59335), .Z(n_59343));
	notech_inv i_11364(.A(n_59335), .Z(n_59338));
	notech_inv i_11361(.A(\nbus_13544[0] ), .Z(n_59335));
	notech_inv i_11358(.A(n_59301), .Z(n_59332));
	notech_inv i_11357(.A(n_59301), .Z(n_59331));
	notech_inv i_11347(.A(n_59301), .Z(n_59321));
	notech_inv i_11346(.A(n_59301), .Z(n_59320));
	notech_inv i_11341(.A(n_59301), .Z(n_59315));
	notech_inv i_11336(.A(n_59301), .Z(n_59310));
	notech_inv i_11335(.A(n_59301), .Z(n_59309));
	notech_inv i_11330(.A(n_59301), .Z(n_59304));
	notech_inv i_11327(.A(\nbus_13544[0] ), .Z(n_59301));
	notech_inv i_11325(.A(n_59210), .Z(n_59298));
	notech_inv i_11323(.A(n_59210), .Z(n_59296));
	notech_inv i_11320(.A(n_59210), .Z(n_59293));
	notech_inv i_11318(.A(n_59210), .Z(n_59291));
	notech_inv i_11314(.A(n_59210), .Z(n_59287));
	notech_inv i_11312(.A(n_59210), .Z(n_59285));
	notech_inv i_11309(.A(n_59210), .Z(n_59282));
	notech_inv i_11307(.A(n_59210), .Z(n_59280));
	notech_inv i_11303(.A(n_59210), .Z(n_59276));
	notech_inv i_11301(.A(n_59210), .Z(n_59274));
	notech_inv i_11298(.A(n_59210), .Z(n_59271));
	notech_inv i_11296(.A(n_59210), .Z(n_59269));
	notech_inv i_11292(.A(n_59210), .Z(n_59265));
	notech_inv i_11290(.A(n_59210), .Z(n_59263));
	notech_inv i_11287(.A(n_59210), .Z(n_59260));
	notech_inv i_11285(.A(n_59210), .Z(n_59258));
	notech_inv i_11280(.A(n_59245), .Z(n_59253));
	notech_inv i_11278(.A(n_59245), .Z(n_59251));
	notech_inv i_11275(.A(n_59245), .Z(n_59248));
	notech_inv i_11273(.A(n_59245), .Z(n_59246));
	notech_inv i_11272(.A(n_59291), .Z(n_59245));
	notech_inv i_11269(.A(n_59245), .Z(n_59242));
	notech_inv i_11267(.A(n_59245), .Z(n_59240));
	notech_inv i_11264(.A(n_59245), .Z(n_59237));
	notech_inv i_11262(.A(n_59245), .Z(n_59235));
	notech_inv i_11258(.A(n_59245), .Z(n_59231));
	notech_inv i_11256(.A(n_59245), .Z(n_59229));
	notech_inv i_11253(.A(n_59245), .Z(n_59226));
	notech_inv i_11251(.A(n_59245), .Z(n_59224));
	notech_inv i_11247(.A(n_59210), .Z(n_59220));
	notech_inv i_11245(.A(n_59210), .Z(n_59218));
	notech_inv i_11242(.A(n_59210), .Z(n_59215));
	notech_inv i_11240(.A(n_59210), .Z(n_59213));
	notech_inv i_11237(.A(n_5406), .Z(n_59210));
	notech_inv i_11235(.A(n_59165), .Z(n_59208));
	notech_inv i_11233(.A(n_59165), .Z(n_59206));
	notech_inv i_11230(.A(n_59165), .Z(n_59203));
	notech_inv i_11228(.A(n_59165), .Z(n_59201));
	notech_inv i_11224(.A(n_59165), .Z(n_59197));
	notech_inv i_11222(.A(n_59165), .Z(n_59195));
	notech_inv i_11218(.A(n_59165), .Z(n_59191));
	notech_inv i_11212(.A(n_59165), .Z(n_59185));
	notech_inv i_11211(.A(n_59165), .Z(n_59184));
	notech_inv i_11207(.A(n_59165), .Z(n_59180));
	notech_inv i_11201(.A(n_59165), .Z(n_59174));
	notech_inv i_11200(.A(n_59165), .Z(n_59173));
	notech_inv i_11195(.A(n_59165), .Z(n_59168));
	notech_inv i_11192(.A(n_5406), .Z(n_59165));
	notech_inv i_11185(.A(n_59156), .Z(n_59157));
	notech_inv i_11184(.A(n_158456195), .Z(n_59156));
	notech_inv i_11182(.A(n_59137), .Z(n_59153));
	notech_inv i_11180(.A(n_59137), .Z(n_59151));
	notech_inv i_11179(.A(n_59137), .Z(n_59150));
	notech_inv i_11175(.A(n_59137), .Z(n_59146));
	notech_inv i_11173(.A(n_59137), .Z(n_59144));
	notech_inv i_11170(.A(n_59137), .Z(n_59141));
	notech_inv i_11168(.A(n_59137), .Z(n_59139));
	notech_inv i_11167(.A(n_59137), .Z(n_59138));
	notech_inv i_11166(.A(n_5276), .Z(n_59137));
	notech_inv i_11159(.A(n_59128), .Z(n_59129));
	notech_inv i_11158(.A(n_13699537), .Z(n_59128));
	notech_inv i_9876(.A(n_57723), .Z(n_57724));
	notech_inv i_9875(.A(n_2994), .Z(n_57723));
	notech_inv i_8994(.A(n_56812), .Z(n_56813));
	notech_inv i_8993(.A(n_1554100859), .Z(n_56812));
	notech_inv i_8984(.A(n_56801), .Z(n_56802));
	notech_inv i_8983(.A(\nbus_13546[0] ), .Z(n_56801));
	notech_inv i_8876(.A(n_56687), .Z(n_56688));
	notech_inv i_8875(.A(n_3302), .Z(n_56687));
	notech_inv i_8871(.A(n_56687), .Z(n_56683));
	notech_inv i_8867(.A(n_56687), .Z(n_56679));
	notech_inv i_8862(.A(n_56687), .Z(n_56674));
	notech_inv i_8858(.A(n_56687), .Z(n_56670));
	notech_inv i_8848(.A(n_56659), .Z(n_56660));
	notech_inv i_8847(.A(n_56640), .Z(n_56659));
	notech_inv i_8843(.A(n_56659), .Z(n_56655));
	notech_inv i_8839(.A(n_56659), .Z(n_56651));
	notech_inv i_8834(.A(n_56659), .Z(n_56646));
	notech_inv i_8830(.A(n_56659), .Z(n_56642));
	notech_inv i_8828(.A(n_56687), .Z(n_56640));
	notech_inv i_8820(.A(n_56631), .Z(n_56632));
	notech_inv i_8819(.A(n_56612), .Z(n_56631));
	notech_inv i_8815(.A(n_56631), .Z(n_56627));
	notech_inv i_8811(.A(n_56631), .Z(n_56623));
	notech_inv i_8806(.A(n_56631), .Z(n_56618));
	notech_inv i_8802(.A(n_56631), .Z(n_56614));
	notech_inv i_8800(.A(n_56687), .Z(n_56612));
	notech_inv i_8736(.A(n_56479), .Z(n_56544));
	notech_inv i_8735(.A(n_56479), .Z(n_56543));
	notech_inv i_8730(.A(n_56479), .Z(n_56538));
	notech_inv i_8725(.A(n_56479), .Z(n_56533));
	notech_inv i_8724(.A(n_56479), .Z(n_56532));
	notech_inv i_8719(.A(n_56479), .Z(n_56527));
	notech_inv i_8714(.A(n_56479), .Z(n_56522));
	notech_inv i_8713(.A(n_56479), .Z(n_56521));
	notech_inv i_8708(.A(n_56479), .Z(n_56516));
	notech_inv i_8702(.A(n_56479), .Z(n_56510));
	notech_inv i_8701(.A(n_56479), .Z(n_56509));
	notech_inv i_8696(.A(n_56479), .Z(n_56504));
	notech_inv i_8691(.A(n_56479), .Z(n_56499));
	notech_inv i_8690(.A(n_56479), .Z(n_56498));
	notech_inv i_8685(.A(n_56479), .Z(n_56493));
	notech_inv i_8680(.A(n_56479), .Z(n_56488));
	notech_inv i_8679(.A(n_56479), .Z(n_56487));
	notech_inv i_8674(.A(n_56479), .Z(n_56482));
	notech_inv i_8671(.A(\nbus_13540[0] ), .Z(n_56479));
	notech_inv i_8668(.A(n_56445), .Z(n_56476));
	notech_inv i_8667(.A(n_56445), .Z(n_56475));
	notech_inv i_8657(.A(n_56445), .Z(n_56465));
	notech_inv i_8656(.A(n_56445), .Z(n_56464));
	notech_inv i_8651(.A(n_56445), .Z(n_56459));
	notech_inv i_8646(.A(n_56445), .Z(n_56454));
	notech_inv i_8645(.A(n_56445), .Z(n_56453));
	notech_inv i_8640(.A(n_56445), .Z(n_56448));
	notech_inv i_8637(.A(\nbus_13540[0] ), .Z(n_56445));
	notech_inv i_7970(.A(n_55781), .Z(n_55782));
	notech_inv i_7969(.A(n_3303), .Z(n_55781));
	notech_inv i_7951(.A(n_55761), .Z(n_55762));
	notech_inv i_7950(.A(n_3246), .Z(n_55761));
	notech_inv i_7943(.A(n_55700), .Z(n_55701));
	notech_inv i_7942(.A(n_3236), .Z(n_55700));
	notech_ao4 i_226107(.A(n_60293), .B(n_44735), .C(n_59258), .D(n_43475), 
		.Z(n_3344));
	notech_ao4 i_126106(.A(n_60293), .B(n_44758), .C(n_59258), .D(n_43473), 
		.Z(n_3345));
	notech_ao4 i_4827835(.A(n_3246), .B(n_43838), .C(n_59258), .D(n_42839), 
		.Z(n_3346));
	notech_ao4 i_4727834(.A(n_3246), .B(n_43841), .C(n_59258), .D(n_42836), 
		.Z(n_3347));
	notech_ao4 i_4627833(.A(n_3246), .B(n_43845), .C(n_59258), .D(n_42834), 
		.Z(n_3348));
	notech_ao4 i_4527832(.A(n_3246), .B(n_43849), .C(n_59253), .D(n_42831), 
		.Z(n_3349));
	notech_ao4 i_4427831(.A(n_3246), .B(n_43851), .C(n_59253), .D(n_42829), 
		.Z(n_3350));
	notech_ao4 i_4327830(.A(n_3246), .B(n_43855), .C(n_59253), .D(n_42827), 
		.Z(n_3351));
	notech_ao4 i_4227829(.A(n_3246), .B(n_43857), .C(n_59258), .D(n_42824), 
		.Z(n_3352));
	notech_ao4 i_4127828(.A(n_3246), .B(n_43861), .C(n_59258), .D(n_42822), 
		.Z(n_3353));
	notech_ao4 i_4027827(.A(n_3236), .B(n_43879), .C(n_59258), .D(n_42819), 
		.Z(n_3354));
	notech_ao4 i_3827825(.A(n_3236), .B(n_43887), .C(n_59258), .D(n_42815), 
		.Z(n_3355));
	notech_ao4 i_3727824(.A(n_3236), .B(n_43893), .C(n_59260), .D(n_42812), 
		.Z(n_3356));
	notech_ao4 i_3627823(.A(n_3236), .B(n_43897), .C(n_59260), .D(n_42810), 
		.Z(n_3357));
	notech_ao4 i_3527822(.A(n_3236), .B(n_43899), .C(n_59260), .D(n_42807), 
		.Z(n_3358));
	notech_ao4 i_3427821(.A(n_3236), .B(n_43903), .C(n_59258), .D(n_42805), 
		.Z(n_3359));
	notech_ao4 i_3327820(.A(n_3236), .B(n_43905), .C(n_59258), .D(n_42803), 
		.Z(n_3360));
	notech_ao4 i_3227819(.A(n_60293), .B(n_2643), .C(n_59258), .D(n_42800), 
		.Z(n_3361));
	notech_ao4 i_3127818(.A(n_60293), .B(n_2635), .C(n_59258), .D(n_42798), 
		.Z(n_3362));
	notech_ao4 i_3027817(.A(n_60293), .B(n_2627), .C(n_59258), .D(n_42795), 
		.Z(n_3363));
	notech_ao4 i_2927816(.A(n_60288), .B(n_2619), .C(n_59253), .D(n_42793), 
		.Z(n_3364));
	notech_ao4 i_2827815(.A(n_60288), .B(n_2611), .C(n_59251), .D(n_42791), 
		.Z(n_3365));
	notech_ao4 i_2727814(.A(n_60288), .B(n_2603), .C(n_59251), .D(n_42788), 
		.Z(n_3366));
	notech_ao4 i_2527812(.A(n_60293), .B(n_2595), .C(n_59251), .D(n_42783), 
		.Z(n_3367));
	notech_ao4 i_2327810(.A(n_60288), .B(n_2577), .C(n_59251), .D(n_42779), 
		.Z(n_3368));
	notech_ao4 i_2027807(.A(n_60293), .B(n_2561), .C(n_59251), .D(n_42771), 
		.Z(n_3369));
	notech_ao4 i_1827805(.A(n_60293), .B(n_2545), .C(n_59251), .D(n_42767), 
		.Z(n_3370));
	notech_ao4 i_1727804(.A(n_60293), .B(n_2537), .C(n_59251), .D(n_42765), 
		.Z(n_3371));
	notech_ao4 i_1627803(.A(n_60295), .B(n_2527), .C(n_59251), .D(n_42763), 
		.Z(n_3372));
	notech_ao4 i_1327800(.A(n_60295), .B(n_2519), .C(n_59251), .D(n_42756), 
		.Z(n_3373));
	notech_ao4 i_1227799(.A(n_60293), .B(n_2511), .C(n_59251), .D(n_42753), 
		.Z(n_3374));
	notech_ao4 i_927796(.A(n_60293), .B(n_2495), .C(n_59253), .D(n_42747), .Z
		(n_3375));
	notech_ao4 i_527792(.A(n_60293), .B(n_2460), .C(n_59253), .D(n_42738), .Z
		(n_3376));
	notech_ao4 i_327790(.A(n_60293), .B(n_2444), .C(n_59253), .D(n_42733), .Z
		(n_3377));
	notech_ao4 i_223134(.A(n_60293), .B(n_44524), .C(n_59253), .D(n_43449), 
		.Z(n_3378));
	notech_ao4 i_123133(.A(n_60288), .B(n_44523), .C(n_59253), .D(n_43448), 
		.Z(n_3379));
	notech_nand3 i_12825766(.A(n_158456195), .B(n_60944), .C(n_1823), .Z(n_3380
		));
	notech_nao3 i_12725765(.A(n_60944), .B(n_1824), .C(n_1538), .Z(n_3381)
		);
	notech_nand3 i_12625764(.A(n_158456195), .B(n_60944), .C(n_1825), .Z(n_3382
		));
	notech_nao3 i_12525763(.A(n_60944), .B(n_1826), .C(n_1538), .Z(n_3383)
		);
	notech_nao3 i_12425762(.A(n_60944), .B(n_1827), .C(n_1538), .Z(n_3384)
		);
	notech_nand3 i_12325761(.A(n_60944), .B(n_13699537), .C(n_1828), .Z(n_3385
		));
	notech_nand2 i_12225760(.A(n_60944), .B(n_1829), .Z(n_3386));
	notech_nao3 i_12125759(.A(n_60944), .B(n_1830), .C(n_1538), .Z(n_3387)
		);
	notech_nand3 i_12025758(.A(n_158456195), .B(n_60944), .C(n_1831), .Z(n_3388
		));
	notech_nand3 i_11925757(.A(n_158456195), .B(n_60944), .C(n_1832), .Z(n_3389
		));
	notech_nand3 i_11825756(.A(n_158456195), .B(n_60944), .C(n_1833), .Z(n_3390
		));
	notech_nand3 i_11725755(.A(n_60944), .B(n_13699537), .C(n_1834), .Z(n_3391
		));
	notech_nand2 i_11625754(.A(n_60944), .B(n_1835), .Z(n_3392));
	notech_nand3 i_11525753(.A(n_1837), .B(n_1537), .C(n_1533), .Z(n_3393)
		);
	notech_nand3 i_11325751(.A(n_1912), .B(n_60944), .C(n_1838), .Z(n_3394)
		);
	notech_nand2 i_11225750(.A(n_60944), .B(n_1840), .Z(n_3395));
	notech_nand3 i_11125749(.A(n_158456195), .B(n_60944), .C(n_1841), .Z(n_3396
		));
	notech_nand2 i_11025748(.A(n_60942), .B(n_1842), .Z(n_3397));
	notech_nand2 i_10925747(.A(n_60942), .B(n_1843), .Z(n_3398));
	notech_nand3 i_10825746(.A(n_1537), .B(n_1533), .C(n_1844), .Z(n_3399)
		);
	notech_nand3 i_10725745(.A(n_60942), .B(n_1845), .C(n_1757), .Z(n_3400)
		);
	notech_nand2 i_10625744(.A(n_60942), .B(n_1847), .Z(n_3401));
	notech_nand3 i_10525743(.A(n_60942), .B(n_13699537), .C(n_1848), .Z(n_3402
		));
	notech_nand3 i_10425742(.A(n_60942), .B(n_13699537), .C(n_1849), .Z(n_3403
		));
	notech_nand3 i_10325741(.A(n_60942), .B(n_13699537), .C(n_1850), .Z(n_3404
		));
	notech_nand3 i_10225740(.A(n_60942), .B(n_13699537), .C(n_1851), .Z(n_3405
		));
	notech_nand2 i_10125739(.A(n_60942), .B(n_1852), .Z(n_3406));
	notech_nand2 i_10025738(.A(n_12254735), .B(n_1853), .Z(n_3407));
	notech_nand2 i_9925737(.A(n_1854), .B(n_12254735), .Z(n_3408));
	notech_nand2 i_9825736(.A(n_60942), .B(n_1855), .Z(n_3409));
	notech_nand2 i_9725735(.A(n_60942), .B(n_1856), .Z(n_3410));
	notech_nand2 i_9625734(.A(n_60942), .B(n_1857), .Z(n_3411));
	notech_nand2 i_9525733(.A(n_60942), .B(n_1858), .Z(n_3412));
	notech_nand2 i_9425732(.A(n_60942), .B(n_1859), .Z(n_3413));
	notech_nand2 i_9325731(.A(n_60942), .B(n_1860), .Z(n_3414));
	notech_nand2 i_9225730(.A(n_60947), .B(n_1861), .Z(n_3415));
	notech_nand2 i_9125729(.A(n_60949), .B(n_1862), .Z(n_3416));
	notech_nand2 i_9025728(.A(n_60949), .B(n_1863), .Z(n_3417));
	notech_nand2 i_8925727(.A(n_60949), .B(n_1864), .Z(n_3418));
	notech_nand3 i_8825726(.A(n_60949), .B(n_1865), .C(n_1710), .Z(n_3419)
		);
	notech_nand3 i_8725725(.A(n_60949), .B(n_1867), .C(n_1707), .Z(n_3420)
		);
	notech_nand3 i_8625724(.A(n_60949), .B(n_1869), .C(n_1704), .Z(n_3421)
		);
	notech_nand3 i_8525723(.A(n_60949), .B(n_1871), .C(n_1701), .Z(n_3422)
		);
	notech_nand3 i_8425722(.A(n_1533), .B(n_1873), .C(n_1698), .Z(n_3423));
	notech_nand3 i_8325721(.A(n_1533), .B(n_1875), .C(n_1695), .Z(n_3424));
	notech_nand3 i_8225720(.A(n_1533), .B(n_1877), .C(n_1692), .Z(n_3425));
	notech_nand3 i_8125719(.A(n_60949), .B(n_188198993), .C(n_1689), .Z(n_3426
		));
	notech_nand3 i_8025718(.A(n_60949), .B(n_13699537), .C(n_188398995), .Z(n_3427
		));
	notech_nand3 i_7925717(.A(n_60949), .B(n_13699537), .C(n_188498996), .Z(n_3428
		));
	notech_nand3 i_7825716(.A(n_60949), .B(n_13699537), .C(n_1885), .Z(n_3429
		));
	notech_nand3 i_7725715(.A(n_60949), .B(n_13699537), .C(n_1886), .Z(n_3430
		));
	notech_nand3 i_7625714(.A(n_60949), .B(n_13699537), .C(n_1887), .Z(n_3431
		));
	notech_nand2 i_7425712(.A(n_60949), .B(n_1888), .Z(n_3432));
	notech_nand2 i_7325711(.A(n_60949), .B(n_1889), .Z(n_3433));
	notech_nao3 i_7225710(.A(n_60949), .B(n_1890), .C(n_1538), .Z(n_3434));
	notech_nand3 i_7125709(.A(n_158456195), .B(n_60947), .C(n_1891), .Z(n_3435
		));
	notech_nand3 i_7025708(.A(n_158456195), .B(n_60947), .C(n_1893), .Z(n_3436
		));
	notech_nao3 i_6925707(.A(n_60947), .B(n_1894), .C(n_1538), .Z(n_3437));
	notech_nao3 i_6825706(.A(n_60947), .B(n_1895), .C(n_1538), .Z(n_3438));
	notech_nand3 i_6725705(.A(n_158456195), .B(n_60947), .C(n_1896), .Z(n_3439
		));
	notech_nand2 i_6625704(.A(n_60947), .B(n_1897), .Z(n_3440));
	notech_nand3 i_5925697(.A(n_158456195), .B(n_60947), .C(n_1911), .Z(n_3441
		));
	notech_nand3 i_5625694(.A(n_60947), .B(n_13699537), .C(n_1916), .Z(n_3442
		));
	notech_nand3 i_5125689(.A(n_158456195), .B(n_60947), .C(n_1917), .Z(n_3443
		));
	notech_nao3 i_4825686(.A(n_60947), .B(n_191898997), .C(n_1538), .Z(n_3444
		));
	notech_nand3 i_4725685(.A(n_59157), .B(n_60947), .C(n_191998998), .Z(n_3445
		));
	notech_nand3 i_4425682(.A(n_60947), .B(n_13699537), .C(n_192098999), .Z(n_3446
		));
	notech_nand3 i_3825676(.A(n_60947), .B(n_59129), .C(n_192199000), .Z(n_3447
		));
	notech_nand3 i_3325671(.A(n_60947), .B(n_59129), .C(n_192299001), .Z(n_3448
		));
	notech_nand3 i_3125669(.A(n_60947), .B(n_59129), .C(n_192399002), .Z(n_3449
		));
	notech_nand3 i_3025668(.A(n_60942), .B(n_59129), .C(n_192499003), .Z(n_3450
		));
	notech_nand2 i_2925667(.A(n_60934), .B(n_192599004), .Z(n_3451));
	notech_nand2 i_2825666(.A(n_60934), .B(n_192699005), .Z(n_3452));
	notech_nand3 i_2725665(.A(n_60934), .B(n_59129), .C(n_192799006), .Z(n_3453
		));
	notech_nand3 i_2625664(.A(n_60934), .B(n_59129), .C(n_192899007), .Z(n_3454
		));
	notech_nand2 i_2525663(.A(n_60934), .B(n_192999008), .Z(n_3455));
	notech_nand2 i_2125659(.A(n_60934), .B(n_193099009), .Z(n_3456));
	notech_nand2 i_1625654(.A(n_60934), .B(n_193199010), .Z(n_3457));
	notech_nand3 i_825646(.A(n_59157), .B(n_60934), .C(n_193299011), .Z(n_3458
		));
	notech_nand3 i_725645(.A(n_59157), .B(n_60934), .C(n_193399012), .Z(n_3459
		));
	notech_nand2 i_625644(.A(n_60934), .B(n_193499013), .Z(n_3460));
	notech_nand2 i_525643(.A(n_60934), .B(n_193599014), .Z(n_3461));
	notech_nand3 i_425642(.A(n_59157), .B(n_60934), .C(n_193699015), .Z(n_3462
		));
	notech_nand3 i_325641(.A(n_59157), .B(n_60934), .C(n_193799016), .Z(n_3463
		));
	notech_nand3 i_225640(.A(n_59157), .B(n_60934), .C(n_193899017), .Z(n_3464
		));
	notech_nand2 i_125639(.A(n_60934), .B(n_193999018), .Z(n_3465));
	notech_ao4 i_21126527(.A(n_60286), .B(n_44658), .C(n_59253), .D(n_44147)
		, .Z(n_3466));
	notech_ao4 i_8526401(.A(n_60286), .B(n_44736), .C(n_59253), .D(n_43965),
		 .Z(n_3467));
	notech_nao3 i_8(.A(n_60888), .B(n_44744), .C(n_60395), .Z(n_5768));
	notech_ao4 i_326108(.A(n_60286), .B(n_44748), .C(n_59253), .D(n_43477), 
		.Z(n_3343));
	notech_nand2 i_3(.A(n_2382), .B(n_60888), .Z(n_5406));
	notech_nand3 i_11(.A(n_60888), .B(n_44744), .C(n_59410), .Z(n_5276));
	notech_or4 i_56(.A(n_2975), .B(pc_req), .C(pg_fault), .D(n_42611), .Z(n_1912
		));
	notech_ao4 i_426109(.A(n_60286), .B(n_44747), .C(n_59253), .D(n_43478), 
		.Z(n_3342));
	notech_and3 i_70731(.A(n_1533), .B(n_230399382), .C(n_229699375), .Z(n_3468
		));
	notech_ao3 i_15679047(.A(n_60888), .B(in128[93]), .C(n_60395), .Z(n_3469
		));
	notech_nor2 i_20479046(.A(n_225599334), .B(n_60286), .Z(n_3470));
	notech_nor2 i_20879045(.A(n_225499333), .B(n_60286), .Z(n_3471));
	notech_nor2 i_20979044(.A(n_225399332), .B(n_60286), .Z(n_3472));
	notech_nor2 i_21679043(.A(n_225299331), .B(n_60286), .Z(n_3473));
	notech_nor2 i_22079042(.A(n_225199330), .B(n_60286), .Z(n_3474));
	notech_ao4 i_3227755(.A(n_2643), .B(n_60286), .C(n_59253), .D(n_42708), 
		.Z(n_3475));
	notech_ao4 i_2127744(.A(n_2569), .B(n_60288), .C(n_59265), .D(n_42697), 
		.Z(n_3476));
	notech_ao4 i_1727740(.A(n_2537), .B(n_60288), .C(n_59265), .D(n_42693), 
		.Z(n_3477));
	notech_ao4 i_12625508(.A(n_60288), .B(n_44520), .C(n_59265), .D(n_43073)
		, .Z(n_3478));
	notech_ao4 i_12425506(.A(n_60288), .B(n_44517), .C(n_59265), .D(n_43069)
		, .Z(n_3479));
	notech_ao4 i_12225504(.A(n_60288), .B(n_44515), .C(n_59265), .D(n_43065)
		, .Z(n_3480));
	notech_ao4 i_12025502(.A(n_60288), .B(n_44512), .C(n_59263), .D(n_43062)
		, .Z(n_3481));
	notech_ao4 i_11825500(.A(n_60286), .B(n_44510), .C(n_59263), .D(n_43058)
		, .Z(n_3482));
	notech_ao4 i_11725499(.A(n_60288), .B(n_44509), .C(n_59263), .D(n_43056)
		, .Z(n_3483));
	notech_ao4 i_11325495(.A(n_60288), .B(n_44504), .C(n_59265), .D(n_43049)
		, .Z(n_3484));
	notech_ao4 i_11225494(.A(n_60288), .B(n_44503), .C(n_59263), .D(n_43047)
		, .Z(n_3485));
	notech_ao4 i_11125493(.A(n_60295), .B(n_44502), .C(n_59265), .D(n_43045)
		, .Z(n_3486));
	notech_ao4 i_11025492(.A(n_60300), .B(n_44501), .C(n_59265), .D(n_43044)
		, .Z(n_3487));
	notech_ao4 i_10925491(.A(n_60300), .B(n_44500), .C(n_59265), .D(n_43041)
		, .Z(n_3488));
	notech_ao4 i_10725489(.A(n_60300), .B(n_44498), .C(n_59269), .D(n_43038)
		, .Z(n_3489));
	notech_ao4 i_10625488(.A(n_60300), .B(n_44497), .C(n_59269), .D(n_43037)
		, .Z(n_3490));
	notech_ao4 i_10525487(.A(n_60300), .B(n_44496), .C(n_59265), .D(n_43034)
		, .Z(n_3491));
	notech_ao4 i_10325485(.A(n_60298), .B(n_44493), .C(n_59265), .D(n_43029)
		, .Z(n_3492));
	notech_ao4 i_10125483(.A(n_60298), .B(n_44491), .C(n_59265), .D(n_43026)
		, .Z(n_3493));
	notech_ao4 i_10025482(.A(n_60298), .B(n_44490), .C(n_59265), .D(n_43025)
		, .Z(n_3494));
	notech_ao4 i_9925481(.A(n_60300), .B(n_44488), .C(n_59265), .D(n_43022),
		 .Z(n_3495));
	notech_ao4 i_9825480(.A(n_60298), .B(n_44487), .C(n_59263), .D(n_43021),
		 .Z(n_3496));
	notech_ao4 i_9725479(.A(n_60300), .B(n_44486), .C(n_59260), .D(n_43019),
		 .Z(n_3497));
	notech_ao4 i_8525467(.A(n_60300), .B(n_44472), .C(n_59260), .D(n_42997),
		 .Z(n_3498));
	notech_ao4 i_8425466(.A(n_60300), .B(n_44470), .C(n_59260), .D(n_42996),
		 .Z(n_3499));
	notech_ao4 i_8325465(.A(n_60304), .B(n_44469), .C(n_59260), .D(n_42993),
		 .Z(n_3500));
	notech_ao4 i_8225464(.A(n_60304), .B(n_44468), .C(n_59260), .D(n_42992),
		 .Z(n_3501));
	notech_ao4 i_8125463(.A(n_60300), .B(n_44467), .C(n_59260), .D(n_42990),
		 .Z(n_3502));
	notech_ao4 i_8025462(.A(n_60300), .B(n_44466), .C(n_59260), .D(n_42989),
		 .Z(n_3503));
	notech_ao4 i_7925461(.A(n_60300), .B(n_44464), .C(n_59260), .D(n_42986),
		 .Z(n_3504));
	notech_ao4 i_7825460(.A(n_60300), .B(n_44463), .C(n_59260), .D(n_42985),
		 .Z(n_3505));
	notech_ao4 i_7725459(.A(n_60300), .B(n_44462), .C(n_59260), .D(n_42983),
		 .Z(n_3506));
	notech_ao4 i_7625458(.A(n_60298), .B(n_44461), .C(n_59263), .D(n_42981),
		 .Z(n_3507));
	notech_ao4 i_7525457(.A(n_60295), .B(n_44460), .C(n_59263), .D(n_42979),
		 .Z(n_3508));
	notech_ao4 i_7425456(.A(n_60295), .B(n_44459), .C(n_59263), .D(n_42978),
		 .Z(n_3509));
	notech_ao4 i_7325455(.A(n_60295), .B(n_44458), .C(n_59263), .D(n_42975),
		 .Z(n_3510));
	notech_ao4 i_7225454(.A(n_60295), .B(n_44457), .C(n_59263), .D(n_42974),
		 .Z(n_3511));
	notech_ao4 i_7125453(.A(n_60295), .B(n_44456), .C(n_59263), .D(n_42972),
		 .Z(n_3512));
	notech_ao4 i_7025452(.A(n_60295), .B(n_44455), .C(n_59260), .D(n_42971),
		 .Z(n_3513));
	notech_ao4 i_6925451(.A(n_60295), .B(n_44454), .C(n_59263), .D(n_42968),
		 .Z(n_3514));
	notech_ao4 i_6825450(.A(n_60295), .B(n_44453), .C(n_59263), .D(n_42967),
		 .Z(n_3515));
	notech_ao4 i_6725449(.A(n_60295), .B(n_44452), .C(n_59263), .D(n_42965),
		 .Z(n_3516));
	notech_ao4 i_6625448(.A(n_60295), .B(n_44451), .C(n_59251), .D(n_42963),
		 .Z(n_3517));
	notech_ao4 i_6525447(.A(n_60298), .B(n_44450), .C(n_59240), .D(n_42961),
		 .Z(n_3518));
	notech_ao4 i_6425446(.A(n_60298), .B(n_44449), .C(n_59240), .D(n_42960),
		 .Z(n_3519));
	notech_ao4 i_6325445(.A(n_60298), .B(n_44448), .C(n_59240), .D(n_42957),
		 .Z(n_3520));
	notech_ao4 i_6225444(.A(n_60298), .B(n_44446), .C(n_59240), .D(n_42956),
		 .Z(n_3521));
	notech_ao4 i_6125443(.A(n_60298), .B(n_44445), .C(n_59240), .D(n_42954),
		 .Z(n_3522));
	notech_ao4 i_6025442(.A(n_60298), .B(n_44444), .C(n_59237), .D(n_42953),
		 .Z(n_3523));
	notech_ao4 i_5925441(.A(n_60295), .B(n_44443), .C(n_59237), .D(n_42950),
		 .Z(n_3524));
	notech_ao4 i_5825440(.A(n_60298), .B(n_44442), .C(n_59240), .D(n_42949),
		 .Z(n_3525));
	notech_ao4 i_5725439(.A(n_60298), .B(n_44440), .C(n_59240), .D(n_42947),
		 .Z(n_3526));
	notech_ao4 i_5625438(.A(n_60298), .B(n_44439), .C(n_59240), .D(n_42945),
		 .Z(n_3527));
	notech_ao4 i_5525437(.A(n_60275), .B(n_44438), .C(n_59242), .D(n_42943),
		 .Z(n_3528));
	notech_ao4 i_5425436(.A(n_60275), .B(n_44437), .C(n_59240), .D(n_42942),
		 .Z(n_3529));
	notech_ao4 i_5325435(.A(n_60275), .B(n_44436), .C(n_59242), .D(n_42939),
		 .Z(n_3530));
	notech_ao4 i_5225434(.A(n_60275), .B(n_44434), .C(n_59242), .D(n_42938),
		 .Z(n_3531));
	notech_ao4 i_5125433(.A(n_60275), .B(n_44433), .C(n_59242), .D(n_42936),
		 .Z(n_3532));
	notech_ao4 i_5025432(.A(n_60272), .B(n_44432), .C(n_59240), .D(n_42935),
		 .Z(n_3533));
	notech_ao4 i_4925431(.A(n_60272), .B(n_44431), .C(n_59240), .D(n_42932),
		 .Z(n_3534));
	notech_ao4 i_4825430(.A(n_60272), .B(n_44430), .C(n_59240), .D(n_42931),
		 .Z(n_3535));
	notech_ao4 i_4725429(.A(n_60275), .B(n_44429), .C(n_59240), .D(n_42929),
		 .Z(n_3536));
	notech_ao4 i_4125423(.A(n_60275), .B(n_44422), .C(n_59240), .D(n_42915),
		 .Z(n_3537));
	notech_ao4 i_4025422(.A(n_60275), .B(n_44421), .C(n_59237), .D(n_42913),
		 .Z(n_3538));
	notech_ao4 i_3925421(.A(n_60275), .B(n_44420), .C(n_59235), .D(n_42912),
		 .Z(n_3539));
	notech_ao4 i_3825420(.A(n_60277), .B(n_44419), .C(n_59235), .D(n_42909),
		 .Z(n_3540));
	notech_ao4 i_3725419(.A(n_60277), .B(n_44418), .C(n_59235), .D(n_42908),
		 .Z(n_3541));
	notech_ao4 i_3625418(.A(n_60277), .B(n_44416), .C(n_59237), .D(n_42906),
		 .Z(n_3542));
	notech_ao4 i_3525417(.A(n_60275), .B(n_44415), .C(n_59235), .D(n_42905),
		 .Z(n_3543));
	notech_ao4 i_3425416(.A(n_60275), .B(n_44414), .C(n_59235), .D(n_42902),
		 .Z(n_3544));
	notech_ao4 i_3325415(.A(n_60275), .B(n_44413), .C(n_59235), .D(n_42901),
		 .Z(n_3545));
	notech_ao4 i_3225414(.A(n_60275), .B(n_44412), .C(n_59235), .D(n_42899),
		 .Z(n_3546));
	notech_ao4 i_3125413(.A(n_60275), .B(n_44410), .C(n_59235), .D(n_42897),
		 .Z(n_3547));
	notech_ao4 i_3025412(.A(n_60272), .B(n_44409), .C(n_59235), .D(n_42895),
		 .Z(n_3548));
	notech_ao4 i_2925411(.A(n_60270), .B(n_44408), .C(n_59237), .D(n_42894),
		 .Z(n_3549));
	notech_ao4 i_2825410(.A(n_60270), .B(n_44407), .C(n_59237), .D(n_42891),
		 .Z(n_3550));
	notech_ao4 i_2725409(.A(n_60270), .B(n_44406), .C(n_59237), .D(n_42890),
		 .Z(n_3551));
	notech_ao4 i_2625408(.A(n_60270), .B(n_44404), .C(n_59237), .D(n_42888),
		 .Z(n_3552));
	notech_ao4 i_2525407(.A(n_60270), .B(n_44403), .C(n_59237), .D(n_42887),
		 .Z(n_3553));
	notech_ao4 i_2425406(.A(n_60270), .B(n_44402), .C(n_59237), .D(n_42884),
		 .Z(n_3554));
	notech_ao4 i_2325405(.A(n_60270), .B(n_44401), .C(n_59237), .D(n_42883),
		 .Z(n_3555));
	notech_ao4 i_2225404(.A(n_60270), .B(n_44400), .C(n_59237), .D(n_42881),
		 .Z(n_3556));
	notech_ao4 i_2125403(.A(n_60270), .B(n_44398), .C(n_59237), .D(n_42879),
		 .Z(n_3557));
	notech_ao4 i_2025402(.A(n_60270), .B(n_44397), .C(n_59237), .D(n_42877),
		 .Z(n_3558));
	notech_ao4 i_1925401(.A(n_60272), .B(n_44396), .C(n_59248), .D(n_42876),
		 .Z(n_3559));
	notech_ao4 i_1825400(.A(n_60272), .B(n_44395), .C(n_59248), .D(n_42873),
		 .Z(n_3560));
	notech_ao4 i_1725399(.A(n_60272), .B(n_44394), .C(n_59248), .D(n_42872),
		 .Z(n_3561));
	notech_ao4 i_1625398(.A(n_60272), .B(n_44392), .C(n_59248), .D(n_42870),
		 .Z(n_3562));
	notech_ao4 i_1525397(.A(n_60272), .B(n_44391), .C(n_59248), .D(n_42869),
		 .Z(n_3563));
	notech_ao4 i_1425396(.A(n_60272), .B(n_44390), .C(n_59246), .D(n_42866),
		 .Z(n_3564));
	notech_ao4 i_1325395(.A(n_60272), .B(n_44389), .C(n_59246), .D(n_42865),
		 .Z(n_3565));
	notech_ao4 i_1225394(.A(n_60272), .B(n_44388), .C(n_59246), .D(n_42863),
		 .Z(n_3566));
	notech_ao4 i_1125393(.A(n_60272), .B(n_44386), .C(n_59248), .D(n_42861),
		 .Z(n_3567));
	notech_ao4 i_1025392(.A(n_60272), .B(n_44385), .C(n_59248), .D(n_42859),
		 .Z(n_3568));
	notech_ao4 i_725389(.A(n_60277), .B(n_44382), .C(n_59248), .D(n_42853), 
		.Z(n_3569));
	notech_ao4 i_525387(.A(n_60283), .B(n_44379), .C(n_59248), .D(n_42848), 
		.Z(n_3570));
	notech_ao4 i_425386(.A(n_60283), .B(n_44378), .C(n_59251), .D(n_42847), 
		.Z(n_3571));
	notech_ao4 i_325385(.A(n_60283), .B(n_44377), .C(n_59251), .D(n_42845), 
		.Z(n_3572));
	notech_ao4 i_225384(.A(n_60283), .B(n_44376), .C(n_59251), .D(n_42843), 
		.Z(n_3573));
	notech_nand3 i_122688(.A(n_1912), .B(n_226099339), .C(n_225999338), .Z(n_3574
		));
	notech_ao4 i_223131(.A(n_60283), .B(n_43445), .C(n_59248), .D(n_43454), 
		.Z(n_3575));
	notech_ao4 i_123130(.A(n_44737), .B(n_43596), .C(n_59248), .D(n_43453), 
		.Z(n_3576));
	notech_ao4 i_20926314(.A(n_60281), .B(n_44655), .C(n_59248), .D(n_43823)
		, .Z(n_3577));
	notech_ao3 i_16278882(.A(n_60888), .B(in128[125]), .C(n_60395), .Z(n_3578
		));
	notech_ao4 i_20726312(.A(n_60281), .B(n_44653), .C(n_59248), .D(n_43819)
		, .Z(n_3579));
	notech_ao3 i_16478880(.A(n_60888), .B(in128[123]), .C(n_60395), .Z(n_3580
		));
	notech_ao4 i_20626311(.A(n_60281), .B(n_44652), .C(n_59248), .D(n_43818)
		, .Z(n_3581));
	notech_ao3 i_16578879(.A(n_60888), .B(in128[122]), .C(n_60395), .Z(n_3582
		));
	notech_ao4 i_20526310(.A(n_60283), .B(n_44650), .C(n_59246), .D(n_43817)
		, .Z(n_3583));
	notech_ao3 i_16678878(.A(n_60893), .B(in128[121]), .C(n_60395), .Z(n_3584
		));
	notech_ao4 i_20426309(.A(n_60283), .B(n_44649), .C(n_59242), .D(n_43815)
		, .Z(n_3585));
	notech_ao3 i_16778877(.A(n_60893), .B(in128[120]), .C(n_60395), .Z(n_3586
		));
	notech_ao4 i_20326308(.A(n_60283), .B(n_44648), .C(n_59242), .D(n_43813)
		, .Z(n_3587));
	notech_ao3 i_16878876(.A(n_60888), .B(in128[119]), .C(n_60395), .Z(n_3588
		));
	notech_ao4 i_20226307(.A(n_60283), .B(n_44647), .C(n_59242), .D(n_43812)
		, .Z(n_3589));
	notech_ao3 i_16978875(.A(n_60888), .B(in128[118]), .C(n_60395), .Z(n_3590
		));
	notech_ao4 i_20126306(.A(n_60286), .B(n_44646), .C(n_59242), .D(n_43811)
		, .Z(n_3591));
	notech_ao3 i_17078874(.A(n_60888), .B(in128[117]), .C(n_60395), .Z(n_3592
		));
	notech_ao4 i_20026305(.A(n_60286), .B(n_44644), .C(n_59242), .D(n_43809)
		, .Z(n_3593));
	notech_ao3 i_17178873(.A(n_60888), .B(in128[116]), .C(n_60395), .Z(n_3594
		));
	notech_ao4 i_19926304(.A(n_60286), .B(n_44643), .C(n_59242), .D(n_43808)
		, .Z(n_3595));
	notech_ao3 i_17278872(.A(n_60882), .B(in128[115]), .C(n_60390), .Z(n_3596
		));
	notech_ao4 i_19826303(.A(n_60283), .B(n_44642), .C(n_59242), .D(n_43807)
		, .Z(n_3597));
	notech_ao3 i_17378871(.A(n_60882), .B(in128[114]), .C(n_60390), .Z(n_3598
		));
	notech_ao4 i_19726302(.A(n_60283), .B(n_44641), .C(n_59242), .D(n_43806)
		, .Z(n_3599));
	notech_ao3 i_17478870(.A(n_60882), .B(in128[113]), .C(n_60390), .Z(n_3600
		));
	notech_ao4 i_19626301(.A(n_60283), .B(n_44640), .C(n_59242), .D(n_43805)
		, .Z(n_3601));
	notech_ao3 i_17578869(.A(n_60882), .B(in128[112]), .C(n_60390), .Z(n_3602
		));
	notech_ao4 i_19526300(.A(n_60283), .B(n_44638), .C(n_59242), .D(n_43803)
		, .Z(n_3603));
	notech_ao3 i_17678868(.A(n_60882), .B(in128[111]), .C(n_60390), .Z(n_3604
		));
	notech_ao4 i_19426299(.A(n_59246), .B(n_43802), .C(n_60283), .D(n_44637)
		, .Z(n_3605));
	notech_ao4 i_19026295(.A(n_59246), .B(n_43796), .C(n_60281), .D(n_44632)
		, .Z(n_3606));
	notech_ao4 i_18926294(.A(n_59246), .B(n_43795), .C(n_60277), .D(n_44631)
		, .Z(n_3607));
	notech_ao4 i_18826293(.A(n_59246), .B(n_43794), .C(n_60277), .D(n_44630)
		, .Z(n_3608));
	notech_ao4 i_18726292(.A(n_59246), .B(n_43793), .C(n_60277), .D(n_44629)
		, .Z(n_3609));
	notech_ao4 i_18626291(.A(n_59246), .B(n_43791), .C(n_60277), .D(n_44628)
		, .Z(n_3610));
	notech_ao4 i_18526290(.A(n_59246), .B(n_43790), .C(n_60277), .D(n_44626)
		, .Z(n_3611));
	notech_ao4 i_18426289(.A(n_59246), .B(n_43789), .C(n_60277), .D(n_44625)
		, .Z(n_3612));
	notech_ao4 i_17826283(.A(n_59246), .B(n_43781), .C(n_60277), .D(n_44618)
		, .Z(n_3613));
	notech_ao4 i_17626281(.A(n_59246), .B(n_43778), .C(n_60277), .D(n_44616)
		, .Z(n_3614));
	notech_ao4 i_17526280(.A(n_59269), .B(n_43777), .C(n_60277), .D(n_44614)
		, .Z(n_3615));
	notech_ao4 i_17426279(.A(n_59291), .B(n_43776), .C(n_60277), .D(n_44613)
		, .Z(n_3616));
	notech_ao4 i_17326278(.A(n_59291), .B(n_43775), .C(n_60281), .D(n_44612)
		, .Z(n_3617));
	notech_ao4 i_17226277(.A(n_59291), .B(n_43773), .C(n_60281), .D(n_44611)
		, .Z(n_3618));
	notech_ao4 i_17126276(.A(n_59291), .B(n_43772), .C(n_60281), .D(n_44610)
		, .Z(n_3619));
	notech_ao4 i_17026275(.A(n_59291), .B(n_43771), .C(n_60281), .D(n_44608)
		, .Z(n_3620));
	notech_ao4 i_16926274(.A(n_59287), .B(n_43770), .C(n_60281), .D(n_44607)
		, .Z(n_3621));
	notech_ao4 i_16826273(.A(n_59287), .B(n_43767), .C(n_60281), .D(n_44606)
		, .Z(n_3622));
	notech_ao4 i_16726272(.A(n_59287), .B(n_43765), .C(n_60281), .D(n_44605)
		, .Z(n_3623));
	notech_ao4 i_16626271(.A(n_59287), .B(n_43763), .C(n_60281), .D(n_44604)
		, .Z(n_3624));
	notech_ao4 i_16526270(.A(n_59287), .B(n_43760), .C(n_60281), .D(n_44602)
		, .Z(n_3625));
	notech_ao4 i_16426269(.A(n_59291), .B(n_43758), .C(n_60281), .D(n_44601)
		, .Z(n_3626));
	notech_ao4 i_16326268(.A(n_59291), .B(n_43755), .C(n_60326), .D(n_44600)
		, .Z(n_3627));
	notech_ao4 i_16226267(.A(n_59291), .B(n_43753), .C(n_60322), .D(n_44599)
		, .Z(n_3628));
	notech_ao4 i_16126266(.A(n_59293), .B(n_43751), .C(n_60326), .D(n_44598)
		, .Z(n_3629));
	notech_ao4 i_16026265(.A(n_59291), .B(n_43748), .C(n_60326), .D(n_44596)
		, .Z(n_3630));
	notech_ao4 i_15926264(.A(n_59291), .B(n_43746), .C(n_60326), .D(n_44595)
		, .Z(n_3631));
	notech_ao4 i_15826263(.A(n_59291), .B(n_43743), .C(n_60322), .D(n_44594)
		, .Z(n_3632));
	notech_ao4 i_15726262(.A(n_59291), .B(n_43741), .C(n_60322), .D(n_44593)
		, .Z(n_3633));
	notech_ao4 i_15626261(.A(n_59291), .B(n_43739), .C(n_60322), .D(n_44592)
		, .Z(n_3634));
	notech_ao4 i_15526260(.A(n_59291), .B(n_43736), .C(n_60322), .D(n_44590)
		, .Z(n_3635));
	notech_ao4 i_15426259(.A(n_59287), .B(n_43734), .C(n_60322), .D(n_44589)
		, .Z(n_3636));
	notech_ao4 i_15326258(.A(n_59285), .B(n_43731), .C(n_60326), .D(n_44588)
		, .Z(n_3637));
	notech_ao4 i_15226257(.A(n_59285), .B(n_43729), .C(n_60326), .D(n_44587)
		, .Z(n_3638));
	notech_ao4 i_15126256(.A(n_59285), .B(n_43727), .C(n_60326), .D(n_44586)
		, .Z(n_3639));
	notech_ao4 i_15026255(.A(n_59285), .B(n_43724), .C(n_60326), .D(n_44584)
		, .Z(n_3640));
	notech_ao4 i_14926254(.A(n_59285), .B(n_43722), .C(n_60326), .D(n_44583)
		, .Z(n_3641));
	notech_ao4 i_14826253(.A(n_59285), .B(n_43719), .C(n_60326), .D(n_44582)
		, .Z(n_3642));
	notech_ao4 i_14726252(.A(n_59285), .B(n_43717), .C(n_60326), .D(n_44581)
		, .Z(n_3643));
	notech_ao4 i_14626251(.A(n_59285), .B(n_43715), .C(n_60326), .D(n_44580)
		, .Z(n_3644));
	notech_ao4 i_14526250(.A(n_59285), .B(n_43712), .C(n_60326), .D(n_44578)
		, .Z(n_3645));
	notech_ao4 i_14426249(.A(n_59285), .B(n_43710), .C(n_60326), .D(n_44577)
		, .Z(n_3646));
	notech_ao4 i_14326248(.A(n_59287), .B(n_43707), .C(n_60322), .D(n_44576)
		, .Z(n_3647));
	notech_ao4 i_14226247(.A(n_59287), .B(n_43705), .C(n_60320), .D(n_44575)
		, .Z(n_3648));
	notech_ao4 i_14126246(.A(n_59287), .B(n_43703), .C(n_60320), .D(n_44574)
		, .Z(n_3649));
	notech_ao4 i_14026245(.A(n_59287), .B(n_43700), .C(n_60320), .D(n_44572)
		, .Z(n_3650));
	notech_ao4 i_13926244(.A(n_59287), .B(n_43698), .C(n_60320), .D(n_44571)
		, .Z(n_3651));
	notech_ao4 i_13826243(.A(n_59285), .B(n_43695), .C(n_60320), .D(n_44570)
		, .Z(n_3652));
	notech_ao4 i_13726242(.A(n_59285), .B(n_43693), .C(n_60320), .D(n_44569)
		, .Z(n_3653));
	notech_ao4 i_13626241(.A(n_59287), .B(n_43691), .C(n_60320), .D(n_44568)
		, .Z(n_3654));
	notech_ao4 i_13526240(.A(n_59287), .B(n_43688), .C(n_60320), .D(n_44566)
		, .Z(n_3655));
	notech_ao4 i_13426239(.A(n_59287), .B(n_43686), .C(n_60320), .D(n_44565)
		, .Z(n_3656));
	notech_ao4 i_13326238(.A(n_59298), .B(n_43683), .C(n_60320), .D(n_44564)
		, .Z(n_3657));
	notech_ao4 i_13226237(.A(n_59296), .B(n_43681), .C(n_60322), .D(n_44563)
		, .Z(n_3658));
	notech_ao4 i_13126236(.A(n_59298), .B(n_43679), .C(n_60322), .D(n_44562)
		, .Z(n_3659));
	notech_ao4 i_13026235(.A(n_59298), .B(n_43676), .C(n_60322), .D(n_44560)
		, .Z(n_3660));
	notech_ao4 i_12926234(.A(n_59298), .B(n_43674), .C(n_60322), .D(n_44559)
		, .Z(n_3661));
	notech_ao4 i_12826233(.A(n_59296), .B(n_43671), .C(n_60322), .D(n_44558)
		, .Z(n_3662));
	notech_ao4 i_12726232(.A(n_59296), .B(n_43669), .C(n_60320), .D(n_44557)
		, .Z(n_3663));
	notech_ao4 i_12626231(.A(n_59296), .B(n_43667), .C(n_60320), .D(n_44556)
		, .Z(n_3664));
	notech_ao4 i_12426229(.A(n_59296), .B(n_43662), .C(n_60320), .D(n_44553)
		, .Z(n_3665));
	notech_ao4 i_11426219(.A(n_59296), .B(n_43638), .C(n_60322), .D(n_44541)
		, .Z(n_3666));
	notech_ao4 i_10726212(.A(n_59298), .B(n_43623), .C(n_60322), .D(n_44533)
		, .Z(n_3667));
	notech_ao4 i_10526210(.A(n_59298), .B(n_43621), .C(n_60328), .D(n_44530)
		, .Z(n_3668));
	notech_ao4 i_10226207(.A(n_59298), .B(n_43617), .C(n_60333), .D(n_44527)
		, .Z(n_3669));
	notech_ao4 i_9926204(.A(n_60331), .B(n_44719), .C(n_59298), .D(n_43614),
		 .Z(n_3670));
	notech_ao3 i_7678966(.A(n_60882), .B(in128[15]), .C(n_60390), .Z(n_3671)
		);
	notech_ao4 i_9826203(.A(n_60333), .B(n_44721), .C(n_59298), .D(n_43613),
		 .Z(n_3672));
	notech_ao3 i_9778946(.A(n_60882), .B(in128[14]), .C(n_60390), .Z(n_3673)
		);
	notech_ao4 i_9726202(.A(n_60333), .B(n_44708), .C(n_59298), .D(n_43611),
		 .Z(n_3674));
	notech_ao3 i_6178980(.A(n_60882), .B(in128[13]), .C(n_60395), .Z(n_3675)
		);
	notech_ao4 i_9626201(.A(n_60333), .B(n_44709), .C(n_59298), .D(n_43610),
		 .Z(n_3676));
	notech_ao3 i_5578986(.A(n_60888), .B(in128[12]), .C(n_60390), .Z(n_3677)
		);
	notech_ao4 i_9526200(.A(n_60331), .B(n_44710), .C(n_59298), .D(n_43609),
		 .Z(n_3678));
	notech_ao3 i_7878964(.A(n_60882), .B(in128[11]), .C(n_60390), .Z(n_3679)
		);
	notech_ao4 i_9426199(.A(n_60331), .B(n_44720), .C(n_59298), .D(n_43608),
		 .Z(n_3680));
	notech_ao3 i_12078923(.A(n_60882), .B(n_59489), .C(n_60390), .Z(n_3681)
		);
	notech_ao4 i_9326198(.A(n_60331), .B(n_44723), .C(n_59298), .D(n_43607),
		 .Z(n_3682));
	notech_ao3 i_12178922(.A(n_60882), .B(in128[9]), .C(n_60395), .Z(n_3683)
		);
	notech_ao4 i_9226197(.A(n_60331), .B(n_44722), .C(n_59296), .D(n_43605),
		 .Z(n_3684));
	notech_ao3 i_7778965(.A(n_60893), .B(in128[8]), .C(n_60399), .Z(n_3685)
		);
	notech_ao4 i_9126196(.A(n_60331), .B(n_44674), .C(n_59293), .D(n_43604),
		 .Z(n_3686));
	notech_ao3 i_19478850(.A(n_60894), .B(in128[7]), .C(n_60400), .Z(n_3687)
		);
	notech_ao4 i_9026195(.A(n_60333), .B(n_44675), .C(n_59293), .D(n_43603),
		 .Z(n_3688));
	notech_ao3 i_19578849(.A(n_60894), .B(in128[6]), .C(n_60399), .Z(n_3689)
		);
	notech_ao4 i_8926194(.A(n_60333), .B(n_44676), .C(n_59293), .D(n_43602),
		 .Z(n_3690));
	notech_ao3 i_19678848(.A(n_60894), .B(in128[5]), .C(n_60399), .Z(n_3691)
		);
	notech_ao4 i_8826193(.A(n_60333), .B(n_44677), .C(n_59293), .D(n_43601),
		 .Z(n_3692));
	notech_ao3 i_19778847(.A(n_60893), .B(in128[4]), .C(n_60399), .Z(n_3693)
		);
	notech_ao4 i_8726192(.A(n_60333), .B(n_44678), .C(n_59293), .D(n_43599),
		 .Z(n_3694));
	notech_ao3 i_19878846(.A(n_60893), .B(in128[3]), .C(n_60400), .Z(n_3695)
		);
	notech_ao4 i_8626191(.A(n_60333), .B(n_44737), .C(n_59293), .D(n_43598),
		 .Z(n_3696));
	notech_ao3 i_9078952(.A(n_60894), .B(in128[2]), .C(n_60400), .Z(n_3697)
		);
	notech_ao4 i_8426189(.A(n_60333), .B(n_44659), .C(n_59293), .D(n_43595),
		 .Z(n_3698));
	notech_ao3 i_8178961(.A(n_60894), .B(in128[0]), .C(n_60400), .Z(n_3699)
		);
	notech_ao4 i_8326188(.A(n_60333), .B(n_44731), .C(n_59293), .D(n_43593),
		 .Z(n_3700));
	notech_ao3 i_15978885(.A(n_60894), .B(mod_dec), .C(n_60400), .Z(n_3701)
		);
	notech_ao4 i_8226187(.A(n_60333), .B(n_44730), .C(n_59293), .D(n_43592),
		 .Z(n_3702));
	notech_ao3 i_16078884(.A(n_60894), .B(sib_dec), .C(n_60400), .Z(n_3703)
		);
	notech_ao4 i_8126186(.A(n_60333), .B(n_44679), .C(n_59293), .D(n_43591),
		 .Z(n_3704));
	notech_ao3 i_14378900(.A(n_60894), .B(\to_acu2_0[80] ), .C(n_60400), .Z(n_3705
		));
	notech_ao4 i_8026185(.A(n_60333), .B(n_44705), .C(n_59296), .D(n_43590),
		 .Z(n_3706));
	notech_ao3 i_14178902(.A(n_60894), .B(\to_acu2_0[79] ), .C(n_60399), .Z(n_3707
		));
	notech_ao4 i_7926184(.A(n_60331), .B(n_44707), .C(n_59296), .D(n_43589),
		 .Z(n_3708));
	notech_ao3 i_14078903(.A(n_60894), .B(\to_acu2_0[78] ), .C(n_60399), .Z(n_3709
		));
	notech_ao4 i_7826183(.A(n_60328), .B(n_44660), .C(n_59296), .D(n_43587),
		 .Z(n_3710));
	notech_ao3 i_19978845(.A(n_60893), .B(\to_acu2_0[77] ), .C(n_60399), .Z(n_3711
		));
	notech_ao4 i_7726182(.A(n_60328), .B(n_44682), .C(n_59296), .D(n_43586),
		 .Z(n_3712));
	notech_ao3 i_13978904(.A(n_60893), .B(\to_acu2_0[76] ), .C(n_60395), .Z(n_3713
		));
	notech_ao4 i_7626181(.A(n_60328), .B(n_44673), .C(n_59296), .D(n_43585),
		 .Z(n_3714));
	notech_ao3 i_14578898(.A(n_60893), .B(\to_acu2_0[75] ), .C(n_60399), .Z(n_3715
		));
	notech_ao4 i_7526180(.A(n_60328), .B(n_44685), .C(n_59293), .D(n_43584),
		 .Z(n_3716));
	notech_ao3 i_10178942(.A(n_60893), .B(\to_acu2_0[74] ), .C(n_60399), .Z(n_3717
		));
	notech_ao4 i_7426179(.A(n_60328), .B(n_44684), .C(n_59293), .D(n_43583),
		 .Z(n_3718));
	notech_ao3 i_9878945(.A(n_60893), .B(\to_acu2_0[73] ), .C(n_60399), .Z(n_3719
		));
	notech_ao4 i_7326178(.A(n_60328), .B(n_44683), .C(n_59293), .D(n_43581),
		 .Z(n_3720));
	notech_ao3 i_13878905(.A(n_60893), .B(\to_acu2_0[72] ), .C(n_60399), .Z(n_3721
		));
	notech_ao4 i_7226177(.A(n_60328), .B(n_44671), .C(n_59296), .D(n_43580),
		 .Z(n_3722));
	notech_ao3 i_7278970(.A(n_60893), .B(\to_acu2_0[71] ), .C(n_60399), .Z(n_3723
		));
	notech_ao4 i_7126176(.A(n_60328), .B(n_44672), .C(n_59296), .D(n_43579),
		 .Z(n_3724));
	notech_ao3 i_14478899(.A(n_60893), .B(\to_acu2_0[70] ), .C(n_60399), .Z(n_3725
		));
	notech_ao4 i_7026175(.A(n_60328), .B(n_44725), .C(n_59285), .D(n_43578),
		 .Z(n_3726));
	notech_ao3 i_14978894(.A(n_60893), .B(\to_acu2_0[69] ), .C(n_60399), .Z(n_3727
		));
	notech_ao4 i_6926174(.A(n_60328), .B(n_44717), .C(n_59274), .D(n_43577),
		 .Z(n_3728));
	notech_ao3 i_13778906(.A(n_60893), .B(\to_acu2_0[68] ), .C(n_60390), .Z(n_3729
		));
	notech_ao4 i_6826173(.A(n_60331), .B(n_44661), .C(n_59274), .D(n_43575),
		 .Z(n_3730));
	notech_ao3 i_20078844(.A(n_60893), .B(\to_acu2_0[67] ), .C(n_60385), .Z(n_3731
		));
	notech_ao4 i_6726172(.A(n_60331), .B(n_44666), .C(n_59274), .D(n_43574),
		 .Z(n_3732));
	notech_ao3 i_20178843(.A(n_60893), .B(\to_acu2_0[66] ), .C(n_60385), .Z(n_3733
		));
	notech_ao4 i_6626171(.A(n_60331), .B(n_44662), .C(n_59274), .D(n_43573),
		 .Z(n_3734));
	notech_ao3 i_20278842(.A(n_60893), .B(\to_acu2_0[65] ), .C(n_60381), .Z(n_3735
		));
	notech_ao4 i_6526170(.A(n_60331), .B(n_44663), .C(n_59274), .D(n_43572),
		 .Z(n_3736));
	notech_ao3 i_20378841(.A(n_60882), .B(\to_acu2_0[64] ), .C(n_60381), .Z(n_3737
		));
	notech_ao4 i_6426169(.A(n_60331), .B(n_44667), .C(n_59271), .D(n_43571),
		 .Z(n_3738));
	notech_ao3 i_20578840(.A(n_60876), .B(\to_acu2_0[63] ), .C(n_60381), .Z(n_3739
		));
	notech_ao4 i_6326168(.A(n_60328), .B(n_44724), .C(n_59271), .D(n_43569),
		 .Z(n_3740));
	notech_ao3 i_15078893(.A(n_60876), .B(\to_acu2_0[62] ), .C(n_60385), .Z(n_3741
		));
	notech_ao4 i_6226167(.A(n_60328), .B(n_44706), .C(n_59271), .D(n_43568),
		 .Z(n_3742));
	notech_ao3 i_13678907(.A(n_60876), .B(\to_acu2_0[61] ), .C(n_60385), .Z(n_3743
		));
	notech_ao4 i_6126166(.A(n_60328), .B(n_44668), .C(n_59274), .D(n_43567),
		 .Z(n_3744));
	notech_ao3 i_20678839(.A(n_60871), .B(\to_acu2_0[60] ), .C(n_60385), .Z(n_3745
		));
	notech_ao4 i_6026165(.A(n_60331), .B(n_44692), .C(n_59271), .D(n_43566),
		 .Z(n_3746));
	notech_ao3 i_13578908(.A(n_60871), .B(\to_acu2_0[59] ), .C(n_60385), .Z(n_3747
		));
	notech_ao4 i_5926164(.A(n_60331), .B(n_44686), .C(n_59274), .D(n_43565),
		 .Z(n_3748));
	notech_ao3 i_6978973(.A(n_60876), .B(\to_acu2_0[58] ), .C(n_60385), .Z(n_3749
		));
	notech_ao4 i_5826163(.A(n_60309), .B(n_44687), .C(n_59274), .D(n_43563),
		 .Z(n_3750));
	notech_ao3 i_11778926(.A(n_60876), .B(\to_acu2_0[57] ), .C(n_60385), .Z(n_3751
		));
	notech_ao4 i_5726162(.A(n_60309), .B(n_44680), .C(n_59274), .D(n_43562),
		 .Z(n_3752));
	notech_ao3 i_14278901(.A(n_60876), .B(\to_acu2_0[56] ), .C(n_60381), .Z(n_3753
		));
	notech_ao4 i_5626161(.A(n_60309), .B(n_44691), .C(n_59276), .D(n_43561),
		 .Z(n_3754));
	notech_ao3 i_5778984(.A(n_60876), .B(\to_acu2_0[55] ), .C(n_60381), .Z(n_3755
		));
	notech_ao4 i_5426159(.A(n_60309), .B(n_44690), .C(n_59276), .D(n_43559),
		 .Z(n_3756));
	notech_ao3 i_8578957(.A(n_60876), .B(\to_acu2_0[53] ), .C(n_60381), .Z(n_3757
		));
	notech_ao4 i_5326158(.A(n_60309), .B(n_44688), .C(n_59274), .D(n_43557),
		 .Z(n_3758));
	notech_ao3 i_6878974(.A(n_60876), .B(\to_acu2_0[52] ), .C(n_60381), .Z(n_3759
		));
	notech_ao4 i_5226157(.A(n_60306), .B(n_44689), .C(n_59274), .D(n_43556),
		 .Z(n_3760));
	notech_ao3 i_8778955(.A(n_60876), .B(\to_acu2_0[51] ), .C(n_60381), .Z(n_3761
		));
	notech_ao4 i_5126156(.A(n_60306), .B(n_44681), .C(n_59274), .D(n_43555),
		 .Z(n_3762));
	notech_ao3 i_8478958(.A(n_60871), .B(\to_acu2_0[50] ), .C(n_60381), .Z(n_3763
		));
	notech_ao4 i_5026155(.A(n_60306), .B(n_44669), .C(n_59274), .D(n_43554),
		 .Z(n_3764));
	notech_ao3 i_20778838(.A(n_60871), .B(\to_acu2_0[49] ), .C(n_60381), .Z(n_3765
		));
	notech_ao4 i_4926154(.A(n_60306), .B(n_44693), .C(n_59274), .D(n_43553),
		 .Z(n_3766));
	notech_ao3 i_13478909(.A(n_60871), .B(\to_acu2_0[48] ), .C(n_60381), .Z(n_3767
		));
	notech_ao4 i_4826153(.A(n_60306), .B(n_44704), .C(n_59271), .D(n_43551),
		 .Z(n_3768));
	notech_ao3 i_8878954(.A(n_60871), .B(\to_acu2_0[47] ), .C(n_60381), .Z(n_3769
		));
	notech_ao4 i_4726152(.A(n_60309), .B(n_44703), .C(n_59269), .D(n_43550),
		 .Z(n_3770));
	notech_ao3 i_7078972(.A(n_60871), .B(\to_acu2_0[46] ), .C(n_60381), .Z(n_3771
		));
	notech_ao4 i_4526150(.A(n_60309), .B(n_44702), .C(n_59269), .D(n_43548),
		 .Z(n_3772));
	notech_ao3 i_5478987(.A(n_60871), .B(\to_acu2_0[44] ), .C(n_60381), .Z(n_3773
		));
	notech_ao4 i_4426149(.A(n_60309), .B(n_44700), .C(n_59269), .D(n_43547),
		 .Z(n_3774));
	notech_ao3 i_5278989(.A(n_60871), .B(\to_acu2_0[43] ), .C(n_60385), .Z(n_3775
		));
	notech_ao4 i_4326148(.A(n_60311), .B(n_44701), .C(n_59269), .D(n_43545),
		 .Z(n_3776));
	notech_ao3 i_15878886(.A(n_60871), .B(\to_acu2_0[42] ), .C(n_60389), .Z(n_3777
		));
	notech_ao4 i_4126146(.A(n_60309), .B(n_44698), .C(n_59269), .D(n_43543),
		 .Z(n_3778));
	notech_ao3 i_15778887(.A(n_60871), .B(\to_acu2_0[40] ), .C(n_60389), .Z(n_3779
		));
	notech_ao4 i_3926144(.A(n_60309), .B(n_44699), .C(n_59269), .D(n_43542),
		 .Z(n_3780));
	notech_ao3 i_15578888(.A(n_60871), .B(\to_acu2_0[38] ), .C(n_60389), .Z(n_3781
		));
	notech_ao4 i_3826143(.A(n_60309), .B(n_44696), .C(n_59269), .D(n_43541),
		 .Z(n_3782));
	notech_ao3 i_15478889(.A(n_60871), .B(\to_acu2_0[37] ), .C(n_60389), .Z(n_3783
		));
	notech_ao4 i_3726142(.A(n_60309), .B(n_44697), .C(n_59269), .D(n_43539),
		 .Z(n_3784));
	notech_ao3 i_15378890(.A(n_60871), .B(\to_acu2_0[36] ), .C(n_60389), .Z(n_3785
		));
	notech_ao4 i_3626141(.A(n_60309), .B(n_44694), .C(n_59269), .D(n_43538),
		 .Z(n_3786));
	notech_ao3 i_15278891(.A(n_60871), .B(\to_acu2_0[35] ), .C(n_60389), .Z(n_3787
		));
	notech_ao4 i_3526140(.A(n_60309), .B(n_44695), .C(n_59269), .D(n_43537),
		 .Z(n_3788));
	notech_ao3 i_15178892(.A(n_60876), .B(\to_acu2_0[34] ), .C(n_60390), .Z(n_3789
		));
	notech_ao4 i_3426139(.A(n_60306), .B(n_44670), .C(n_59271), .D(n_43536),
		 .Z(n_3790));
	notech_ao3 i_21078837(.A(n_60881), .B(\to_acu2_0[33] ), .C(n_60390), .Z(n_3791
		));
	notech_ao4 i_3326138(.A(n_60304), .B(n_44664), .C(n_59271), .D(n_43535),
		 .Z(n_3792));
	notech_ao3 i_21178836(.A(n_60881), .B(\to_acu2_0[32] ), .C(n_60390), .Z(n_3793
		));
	notech_ao4 i_3226137(.A(n_60304), .B(n_44665), .C(n_59271), .D(n_43532),
		 .Z(n_3794));
	notech_ao3 i_21278835(.A(n_60881), .B(\to_acu2_0[31] ), .C(n_60389), .Z(n_3795
		));
	notech_ao4 i_2627813(.A(n_225199330), .B(n_60304), .C(n_59271), .D(n_42786
		), .Z(n_3796));
	notech_ao4 i_2427811(.A(n_60304), .B(n_2585), .C(n_59271), .D(n_42781), 
		.Z(n_3797));
	notech_ao4 i_2227809(.A(n_225299331), .B(n_60304), .C(n_59271), .D(n_42776
		), .Z(n_3798));
	notech_ao4 i_2127808(.A(n_60304), .B(n_2569), .C(n_59269), .D(n_42774), 
		.Z(n_3799));
	notech_ao4 i_1927806(.A(n_60304), .B(n_2553), .C(n_59271), .D(n_42769), 
		.Z(n_3800));
	notech_ao4 i_1527802(.A(n_225399332), .B(n_60304), .C(n_59271), .D(n_42761
		), .Z(n_3801));
	notech_ao4 i_1427801(.A(n_225499333), .B(n_60304), .C(n_59271), .D(n_42759
		), .Z(n_3802));
	notech_ao4 i_1127798(.A(n_60304), .B(n_2503), .C(n_59282), .D(n_42751), 
		.Z(n_3803));
	notech_ao4 i_1027797(.A(n_225599334), .B(n_60306), .C(n_59282), .D(n_42749
		), .Z(n_3804));
	notech_ao4 i_827795(.A(n_60306), .B(n_2484), .C(n_59282), .D(n_42745), .Z
		(n_3805));
	notech_ao4 i_727794(.A(n_60306), .B(n_2476), .C(n_59282), .D(n_42743), .Z
		(n_3806));
	notech_ao4 i_627793(.A(n_60306), .B(n_2468), .C(n_59282), .D(n_42741), .Z
		(n_3807));
	notech_ao4 i_427791(.A(n_60306), .B(n_2452), .C(n_59280), .D(n_42736), .Z
		(n_3808));
	notech_ao4 i_227789(.A(n_60304), .B(n_2436), .C(n_59280), .D(n_42731), .Z
		(n_3809));
	notech_ao4 i_127788(.A(n_60304), .B(n_2428), .C(n_59280), .D(n_42729), .Z
		(n_3810));
	notech_ao4 i_13526451(.A(n_59280), .B(n_44050), .C(n_60306), .D(n_44566)
		, .Z(n_3811));
	notech_ao4 i_12426440(.A(n_59280), .B(n_44036), .C(n_60306), .D(n_44553)
		, .Z(n_3812));
	notech_ao4 i_12326439(.A(n_59282), .B(n_44035), .C(n_60306), .D(n_44552)
		, .Z(n_3813));
	notech_ao4 i_12226438(.A(n_59282), .B(n_44033), .C(n_60311), .D(n_44551)
		, .Z(n_3814));
	notech_ao4 i_12126437(.A(n_59282), .B(n_44030), .C(n_60317), .D(n_44550)
		, .Z(n_3815));
	notech_ao4 i_12026436(.A(n_59285), .B(n_44028), .C(n_60317), .D(n_44548)
		, .Z(n_3816));
	notech_ao4 i_11926435(.A(n_59282), .B(n_44025), .C(n_60317), .D(n_44547)
		, .Z(n_3817));
	notech_ao4 i_11826434(.A(n_59282), .B(n_44023), .C(n_60317), .D(n_44546)
		, .Z(n_3818));
	notech_ao4 i_11726433(.A(n_59282), .B(n_44021), .C(n_60317), .D(n_44545)
		, .Z(n_3819));
	notech_ao4 i_11626432(.A(n_59282), .B(n_44018), .C(n_60315), .D(n_44544)
		, .Z(n_3820));
	notech_ao4 i_11526431(.A(n_59282), .B(n_44016), .C(n_60315), .D(n_44542)
		, .Z(n_3821));
	notech_ao4 i_11426430(.A(n_59282), .B(n_44013), .C(n_60315), .D(n_44541)
		, .Z(n_3822));
	notech_ao4 i_11326429(.A(n_59280), .B(n_44012), .C(n_60315), .D(n_44540)
		, .Z(n_3823));
	notech_ao4 i_11226428(.A(n_59276), .B(n_44010), .C(n_60315), .D(n_44539)
		, .Z(n_3824));
	notech_ao4 i_11026426(.A(n_59276), .B(n_44005), .C(n_60317), .D(n_44536)
		, .Z(n_3825));
	notech_ao4 i_10826424(.A(n_59276), .B(n_44000), .C(n_60317), .D(n_44534)
		, .Z(n_3826));
	notech_ao4 i_10626422(.A(n_59276), .B(n_43997), .C(n_60317), .D(n_44532)
		, .Z(n_3827));
	notech_ao4 i_10526421(.A(n_59276), .B(n_43994), .C(n_60320), .D(n_44530)
		, .Z(n_3828));
	notech_ao4 i_10426420(.A(n_59276), .B(n_43993), .C(n_60317), .D(n_44529)
		, .Z(n_3829));
	notech_ao4 i_10326419(.A(n_59276), .B(n_43991), .C(n_60317), .D(n_44528)
		, .Z(n_3830));
	notech_ao4 i_10226418(.A(n_59276), .B(n_43988), .C(n_60317), .D(n_44527)
		, .Z(n_3831));
	notech_ao4 i_10126417(.A(n_59276), .B(n_43987), .C(n_60317), .D(n_44526)
		, .Z(n_3832));
	notech_ao4 i_9726413(.A(n_60317), .B(n_44708), .C(n_59276), .D(n_43980),
		 .Z(n_3833));
	notech_ao4 i_9626412(.A(n_60317), .B(n_44709), .C(n_59280), .D(n_43979),
		 .Z(n_3834));
	notech_ao4 i_9526411(.A(n_60315), .B(n_44710), .C(n_59280), .D(n_43977),
		 .Z(n_3835));
	notech_ao4 i_9426410(.A(n_60311), .B(n_44720), .C(n_59280), .D(n_43976),
		 .Z(n_3836));
	notech_ao4 i_9326409(.A(n_60311), .B(n_44723), .C(n_59280), .D(n_43975),
		 .Z(n_3837));
	notech_ao4 i_6726383(.A(n_60311), .B(n_44666), .C(n_59280), .D(n_43944),
		 .Z(n_3838));
	notech_ao4 i_6426380(.A(n_60311), .B(n_44667), .C(n_59276), .D(n_43940),
		 .Z(n_3839));
	notech_ao4 i_6226378(.A(n_60311), .B(n_44706), .C(n_59276), .D(n_43938),
		 .Z(n_3840));
	notech_ao4 i_6126377(.A(n_60311), .B(n_44668), .C(n_59280), .D(n_43937),
		 .Z(n_3841));
	notech_ao4 i_5826374(.A(n_60311), .B(n_44687), .C(n_59280), .D(n_43933),
		 .Z(n_3842));
	notech_ao4 i_5726373(.A(n_60311), .B(n_44680), .C(n_59280), .D(n_43932),
		 .Z(n_3843));
	notech_ao4 i_5626372(.A(n_60311), .B(n_44691), .C(n_59197), .D(n_43931),
		 .Z(n_3844));
	notech_ao4 i_5326369(.A(n_60311), .B(n_44688), .C(n_59197), .D(n_43927),
		 .Z(n_3845));
	notech_ao4 i_5226368(.A(n_60315), .B(n_44689), .C(n_59191), .D(n_43926),
		 .Z(n_3846));
	notech_ao4 i_5126367(.A(n_60315), .B(n_44681), .C(n_59191), .D(n_43925),
		 .Z(n_3847));
	notech_ao4 i_5026366(.A(n_60315), .B(n_44669), .C(n_59191), .D(n_43923),
		 .Z(n_3848));
	notech_ao4 i_4226358(.A(n_59197), .B(n_43913), .C(n_60315), .D(n_44749),
		 .Z(n_3849));
	notech_ao4 i_4126357(.A(n_60315), .B(n_44698), .C(n_59185), .D(n_43909),
		 .Z(n_3850));
	notech_ao4 i_3526351(.A(n_60311), .B(n_44695), .C(n_59197), .D(n_43901),
		 .Z(n_3851));
	notech_ao4 i_3426350(.A(n_60311), .B(n_44670), .C(n_59197), .D(n_43898),
		 .Z(n_3852));
	notech_ao4 i_2926345(.A(n_59197), .B(n_43886), .C(n_60315), .D(n_44757),
		 .Z(n_3853));
	notech_ao4 i_2826344(.A(n_59191), .B(n_43884), .C(n_60315), .D(n_44746),
		 .Z(n_3854));
	notech_ao4 i_2726343(.A(n_59191), .B(n_43881), .C(n_60315), .D(n_44743),
		 .Z(n_3855));
	notech_ao4 i_2626342(.A(n_59191), .B(n_43878), .C(n_60270), .D(n_44755),
		 .Z(n_3856));
	notech_ao4 i_2526341(.A(n_59191), .B(n_43875), .C(n_60225), .D(n_44756),
		 .Z(n_3857));
	notech_ao4 i_2426340(.A(n_59191), .B(n_43873), .C(n_60225), .D(n_44741),
		 .Z(n_3858));
	notech_ao4 i_2326339(.A(n_59191), .B(n_43871), .C(n_60225), .D(n_44740),
		 .Z(n_3859));
	notech_ao4 i_2226338(.A(n_59191), .B(n_43868), .C(n_60225), .D(n_44742),
		 .Z(n_3860));
	notech_ao4 i_2026336(.A(n_59191), .B(n_43863), .C(n_60225), .D(n_44753),
		 .Z(n_3861));
	notech_ao4 i_526110(.A(n_60225), .B(n_44751), .C(n_59191), .D(n_43481), 
		.Z(n_3341));
	notech_nand2 i_6257(.A(n_43431), .B(idx_deco[1]), .Z(n_1669));
	notech_and2 i_66549(.A(n_43434), .B(idx_deco[0]), .Z(n_5405));
	notech_ao4 i_65958(.A(n_2398), .B(n_3028), .C(n_42549), .D(n_3025), .Z(n_1915
		));
	notech_ao3 i_127188(.A(n_60881), .B(\nbus_12406[0] ), .C(n_60389), .Z(n_1914
		));
	notech_ao4 i_1(.A(n_2975), .B(n_2401), .C(n_2976), .D(n_2970), .Z(n_1913
		));
	notech_ao3 i_132(.A(n_60881), .B(\to_acu2_0[6] ), .C(n_60385), .Z(n_1910
		));
	notech_ao3 i_191(.A(n_60881), .B(repz), .C(n_60385), .Z(n_1909));
	notech_ao3 i_290(.A(n_60882), .B(\to_acu2_0[3] ), .C(n_60385), .Z(n_1908
		));
	notech_ao4 i_626111(.A(n_60221), .B(n_44734), .C(n_59191), .D(n_43482), 
		.Z(n_3340));
	notech_ao3 i_293(.A(n_60882), .B(opz[0]), .C(n_60385), .Z(n_1907));
	notech_ao3 i_300(.A(n_60882), .B(\to_acu2_0[4] ), .C(n_60385), .Z(n_1906
		));
	notech_ao4 i_726112(.A(n_60225), .B(n_44733), .C(n_59185), .D(n_43484), 
		.Z(n_3339));
	notech_ao3 i_321(.A(in128[1]), .B(in128[2]), .C(n_60225), .Z(n_1905));
	notech_ao3 i_324(.A(n_60882), .B(\to_acu2_0[0] ), .C(n_60389), .Z(n_1904
		));
	notech_ao4 i_826113(.A(n_60225), .B(n_44759), .C(n_59185), .D(n_43485), 
		.Z(n_3338));
	notech_ao3 i_335(.A(n_60882), .B(\to_acu2_0[2] ), .C(n_60389), .Z(n_1903
		));
	notech_ao3 i_38180639(.A(n_60882), .B(\to_acu2_0[7] ), .C(n_60389), .Z(n_3337
		));
	notech_ao3 i_336(.A(n_60881), .B(opz[1]), .C(n_60389), .Z(n_1902));
	notech_ao3 i_342(.A(n_60881), .B(\to_acu2_0[1] ), .C(n_60389), .Z(n_1901
		));
	notech_ao3 i_373(.A(n_60881), .B(\to_acu2_0[5] ), .C(n_60389), .Z(n_1900
		));
	notech_ao3 i_397(.A(n_60881), .B(\to_acu2_0[54] ), .C(n_60413), .Z(n_1899
		));
	notech_and2 i_104(.A(twobyte), .B(n_44729), .Z(n_1898));
	notech_ao4 i_926114(.A(n_60227), .B(n_44726), .C(n_59185), .D(n_43488), 
		.Z(n_3336));
	notech_ao3 i_26180640(.A(n_60876), .B(\to_acu2_0[8] ), .C(n_60413), .Z(n_3335
		));
	notech_ao4 i_1026115(.A(n_60227), .B(n_44728), .C(n_59185), .D(n_43489),
		 .Z(n_3334));
	notech_ao3 i_190(.A(n_60881), .B(in128[127]), .C(n_60413), .Z(n_48352)
		);
	notech_ao3 i_105(.A(n_60881), .B(in128[1]), .C(n_60413), .Z(n_47596));
	notech_ao3 i_34380641(.A(n_60881), .B(\to_acu2_0[9] ), .C(n_60413), .Z(n_3333
		));
	notech_ao3 i_225256(.A(n_60881), .B(udeco[1]), .C(n_60413), .Z(n_41886)
		);
	notech_ao3 i_325257(.A(n_60881), .B(udeco[2]), .C(n_60417), .Z(n_41892)
		);
	notech_ao3 i_425258(.A(n_60881), .B(udeco[3]), .C(n_60417), .Z(n_41898)
		);
	notech_ao3 i_525259(.A(n_60881), .B(udeco[4]), .C(n_60417), .Z(n_41904)
		);
	notech_ao3 i_725261(.A(n_60881), .B(udeco[6]), .C(n_60417), .Z(n_41916)
		);
	notech_ao3 i_1025264(.A(n_60894), .B(udeco[9]), .C(n_60417), .Z(n_41934)
		);
	notech_ao3 i_1125265(.A(n_60915), .B(udeco[10]), .C(n_60413), .Z(n_41940
		));
	notech_ao3 i_1225266(.A(n_60915), .B(udeco[11]), .C(n_60413), .Z(n_41946
		));
	notech_ao3 i_1325267(.A(n_60915), .B(udeco[12]), .C(n_60409), .Z(n_41952
		));
	notech_ao3 i_1425268(.A(n_60910), .B(udeco[13]), .C(n_60409), .Z(n_41958
		));
	notech_ao3 i_1525269(.A(n_60910), .B(udeco[14]), .C(n_60409), .Z(n_41964
		));
	notech_ao3 i_1625270(.A(n_60915), .B(udeco[15]), .C(n_60413), .Z(n_41970
		));
	notech_ao3 i_1725271(.A(n_60915), .B(udeco[16]), .C(n_60413), .Z(n_41976
		));
	notech_ao3 i_1825272(.A(n_60915), .B(udeco[17]), .C(n_60413), .Z(n_41982
		));
	notech_ao3 i_1925273(.A(n_60915), .B(udeco[18]), .C(n_60413), .Z(n_41988
		));
	notech_ao3 i_2025274(.A(n_60915), .B(udeco[19]), .C(n_60413), .Z(n_41994
		));
	notech_ao3 i_2125275(.A(n_60915), .B(udeco[20]), .C(n_60413), .Z(n_42000
		));
	notech_ao3 i_2225276(.A(n_60915), .B(udeco[21]), .C(n_60417), .Z(n_42006
		));
	notech_ao3 i_2325277(.A(n_60910), .B(udeco[22]), .C(n_60418), .Z(n_42012
		));
	notech_ao3 i_2425278(.A(n_60910), .B(udeco[23]), .C(n_60418), .Z(n_42018
		));
	notech_ao3 i_2525279(.A(n_60910), .B(udeco[24]), .C(n_60418), .Z(n_42024
		));
	notech_ao3 i_2625280(.A(n_60910), .B(udeco[25]), .C(n_60418), .Z(n_42030
		));
	notech_ao3 i_2725281(.A(n_60905), .B(udeco[26]), .C(n_60418), .Z(n_42036
		));
	notech_ao3 i_2825282(.A(n_60905), .B(udeco[27]), .C(n_60418), .Z(n_42042
		));
	notech_ao3 i_2925283(.A(n_60905), .B(udeco[28]), .C(n_60418), .Z(n_42048
		));
	notech_ao3 i_3025284(.A(n_60910), .B(udeco[29]), .C(n_60418), .Z(n_42054
		));
	notech_ao3 i_3125285(.A(n_60910), .B(udeco[30]), .C(n_60418), .Z(n_42060
		));
	notech_ao3 i_3225286(.A(n_60910), .B(udeco[31]), .C(n_60418), .Z(n_42066
		));
	notech_ao3 i_3325287(.A(n_60910), .B(udeco[32]), .C(n_60418), .Z(n_42072
		));
	notech_ao3 i_3425288(.A(n_60910), .B(udeco[33]), .C(n_60417), .Z(n_42078
		));
	notech_ao3 i_3525289(.A(n_60910), .B(udeco[34]), .C(n_60417), .Z(n_42084
		));
	notech_ao3 i_3625290(.A(n_60915), .B(udeco[35]), .C(n_60417), .Z(n_42090
		));
	notech_ao3 i_3725291(.A(n_60916), .B(udeco[36]), .C(n_60417), .Z(n_42096
		));
	notech_ao3 i_3825292(.A(n_60916), .B(udeco[37]), .C(n_60417), .Z(n_42102
		));
	notech_ao3 i_3925293(.A(n_60916), .B(udeco[38]), .C(n_60417), .Z(n_42108
		));
	notech_ao3 i_4025294(.A(n_60916), .B(udeco[39]), .C(n_60418), .Z(n_42114
		));
	notech_ao3 i_4125295(.A(n_60916), .B(udeco[40]), .C(n_60418), .Z(n_42120
		));
	notech_ao3 i_4725301(.A(n_60916), .B(udeco[46]), .C(n_60418), .Z(n_42156
		));
	notech_ao3 i_4825302(.A(n_60916), .B(udeco[47]), .C(n_60417), .Z(n_42162
		));
	notech_ao3 i_4925303(.A(n_60916), .B(udeco[48]), .C(n_60417), .Z(n_42168
		));
	notech_ao3 i_5025304(.A(n_60916), .B(udeco[49]), .C(n_60409), .Z(n_42174
		));
	notech_ao3 i_5125305(.A(n_60916), .B(udeco[50]), .C(n_60404), .Z(n_42180
		));
	notech_ao3 i_5225306(.A(n_60916), .B(udeco[51]), .C(n_60404), .Z(n_42186
		));
	notech_ao3 i_5325307(.A(n_60916), .B(udeco[52]), .C(n_60404), .Z(n_42192
		));
	notech_ao3 i_5425308(.A(n_60916), .B(udeco[53]), .C(n_60404), .Z(n_42198
		));
	notech_ao3 i_5525309(.A(n_60915), .B(udeco[54]), .C(n_60404), .Z(n_42204
		));
	notech_ao3 i_5625310(.A(n_60915), .B(udeco[55]), .C(n_60404), .Z(n_42210
		));
	notech_ao3 i_5725311(.A(n_60915), .B(udeco[56]), .C(n_60404), .Z(n_42216
		));
	notech_ao3 i_5825312(.A(n_60915), .B(udeco[57]), .C(n_60408), .Z(n_42222
		));
	notech_ao3 i_5925313(.A(n_60915), .B(udeco[58]), .C(n_60404), .Z(n_42228
		));
	notech_ao3 i_6025314(.A(n_60915), .B(udeco[59]), .C(n_60404), .Z(n_42234
		));
	notech_ao3 i_6125315(.A(n_60916), .B(udeco[60]), .C(n_60404), .Z(n_42240
		));
	notech_ao3 i_6225316(.A(n_60916), .B(udeco[61]), .C(n_60400), .Z(n_42246
		));
	notech_ao3 i_6325317(.A(n_60916), .B(udeco[62]), .C(n_60400), .Z(n_42252
		));
	notech_ao3 i_6425318(.A(n_60915), .B(udeco[63]), .C(n_60400), .Z(n_42258
		));
	notech_ao3 i_6525319(.A(n_60916), .B(udeco[64]), .C(n_60400), .Z(n_42264
		));
	notech_ao3 i_6625320(.A(n_60916), .B(udeco[65]), .C(n_60400), .Z(n_42270
		));
	notech_ao3 i_6725321(.A(n_60905), .B(udeco[66]), .C(n_60400), .Z(n_42276
		));
	notech_ao3 i_6825322(.A(n_60899), .B(udeco[67]), .C(n_60404), .Z(n_42282
		));
	notech_ao3 i_6925323(.A(n_60899), .B(udeco[68]), .C(n_60404), .Z(n_42288
		));
	notech_ao3 i_7025324(.A(n_60899), .B(udeco[69]), .C(n_60404), .Z(n_42294
		));
	notech_ao3 i_7125325(.A(n_60899), .B(udeco[70]), .C(n_60400), .Z(n_42300
		));
	notech_ao3 i_7225326(.A(n_60899), .B(udeco[71]), .C(n_60404), .Z(n_42306
		));
	notech_ao3 i_7325327(.A(n_60899), .B(udeco[72]), .C(n_60408), .Z(n_42312
		));
	notech_ao3 i_7425328(.A(n_60904), .B(udeco[73]), .C(n_60409), .Z(n_42318
		));
	notech_ao3 i_7525329(.A(n_60904), .B(udeco[74]), .C(n_60409), .Z(n_42324
		));
	notech_ao3 i_7625330(.A(n_60904), .B(udeco[75]), .C(n_60409), .Z(n_42330
		));
	notech_ao3 i_7725331(.A(n_60904), .B(udeco[76]), .C(n_60408), .Z(n_42336
		));
	notech_ao3 i_7825332(.A(n_60904), .B(udeco[77]), .C(n_60409), .Z(n_42342
		));
	notech_ao3 i_7925333(.A(n_60904), .B(udeco[78]), .C(n_60409), .Z(n_42348
		));
	notech_ao3 i_8025334(.A(n_60899), .B(udeco[79]), .C(n_60409), .Z(n_42354
		));
	notech_ao3 i_8125335(.A(n_60894), .B(udeco[80]), .C(n_60409), .Z(n_42360
		));
	notech_ao3 i_8225336(.A(n_60894), .B(udeco[81]), .C(n_60409), .Z(n_42366
		));
	notech_ao3 i_8325337(.A(n_60894), .B(udeco[82]), .C(n_60409), .Z(n_42372
		));
	notech_ao3 i_8425338(.A(n_60894), .B(udeco[83]), .C(n_60409), .Z(n_42378
		));
	notech_ao3 i_8525339(.A(n_60894), .B(udeco[84]), .C(n_60408), .Z(n_42384
		));
	notech_ao3 i_9725351(.A(n_60894), .B(udeco[96]), .C(n_60408), .Z(n_42456
		));
	notech_ao3 i_9825352(.A(n_60899), .B(udeco[97]), .C(n_60408), .Z(n_42462
		));
	notech_ao3 i_9925353(.A(n_60899), .B(udeco[98]), .C(n_60408), .Z(n_42468
		));
	notech_ao3 i_10025354(.A(n_60899), .B(udeco[99]), .C(n_60408), .Z(n_42474
		));
	notech_ao3 i_10125355(.A(n_60894), .B(udeco[100]), .C(n_60408), .Z(n_42480
		));
	notech_ao3 i_10325357(.A(n_60899), .B(udeco[102]), .C(n_60408), .Z(n_42492
		));
	notech_ao3 i_10525359(.A(n_60899), .B(udeco[104]), .C(n_60408), .Z(n_42504
		));
	notech_ao3 i_10625360(.A(n_60904), .B(udeco[105]), .C(n_60408), .Z(n_42510
		));
	notech_ao3 i_10725361(.A(n_60905), .B(udeco[106]), .C(n_60408), .Z(n_42516
		));
	notech_ao3 i_10925363(.A(n_60905), .B(udeco[108]), .C(n_60408), .Z(n_42528
		));
	notech_ao3 i_11025364(.A(n_60905), .B(udeco[109]), .C(n_60346), .Z(n_42534
		));
	notech_ao3 i_11125365(.A(n_60905), .B(udeco[110]), .C(n_60346), .Z(n_42540
		));
	notech_ao3 i_11225366(.A(n_60905), .B(udeco[111]), .C(n_60346), .Z(n_42546
		));
	notech_ao3 i_11325367(.A(n_60905), .B(udeco[112]), .C(n_60346), .Z(n_42552
		));
	notech_ao3 i_11725371(.A(n_60905), .B(udeco[116]), .C(n_60346), .Z(n_42576
		));
	notech_ao3 i_11825372(.A(n_60905), .B(udeco[117]), .C(n_60346), .Z(n_42582
		));
	notech_ao3 i_12025374(.A(n_60905), .B(udeco[119]), .C(n_60346), .Z(n_42594
		));
	notech_ao3 i_12225376(.A(n_60905), .B(udeco[121]), .C(n_60346), .Z(n_42606
		));
	notech_ao3 i_12425378(.A(n_60905), .B(udeco[123]), .C(n_60346), .Z(n_42618
		));
	notech_ao3 i_12625380(.A(n_60905), .B(udeco[125]), .C(n_60346), .Z(n_42630
		));
	notech_nor2 i_195(.A(n_2428), .B(n_60227), .Z(n_44375));
	notech_nor2 i_196(.A(n_2436), .B(n_60227), .Z(n_44381));
	notech_nor2 i_197(.A(n_2444), .B(n_60227), .Z(n_44387));
	notech_nor2 i_198(.A(n_2452), .B(n_60225), .Z(n_44393));
	notech_nor2 i_199(.A(n_2460), .B(n_60225), .Z(n_44399));
	notech_nor2 i_200(.A(n_2468), .B(n_60225), .Z(n_44405));
	notech_nor2 i_201(.A(n_2476), .B(n_60225), .Z(n_44411));
	notech_nor2 i_202(.A(n_2484), .B(n_60225), .Z(n_44417));
	notech_nor2 i_203(.A(n_2495), .B(n_60221), .Z(n_44423));
	notech_nor2 i_205(.A(n_2503), .B(n_60219), .Z(n_44435));
	notech_nor2 i_206(.A(n_2511), .B(n_60219), .Z(n_44441));
	notech_nor2 i_207(.A(n_2519), .B(n_60219), .Z(n_44447));
	notech_nor2 i_210(.A(n_2527), .B(n_60221), .Z(n_44465));
	notech_nor2 i_211(.A(n_2537), .B(n_60221), .Z(n_44471));
	notech_nor2 i_212(.A(n_2545), .B(n_60219), .Z(n_44477));
	notech_nor2 i_213(.A(n_2553), .B(n_60219), .Z(n_44483));
	notech_nor2 i_214(.A(n_2561), .B(n_60219), .Z(n_44489));
	notech_nor2 i_215(.A(n_2569), .B(n_60219), .Z(n_44495));
	notech_nor2 i_217(.A(n_2577), .B(n_60219), .Z(n_44507));
	notech_nor2 i_218(.A(n_2585), .B(n_60221), .Z(n_44513));
	notech_nor2 i_219(.A(n_2595), .B(n_60221), .Z(n_44519));
	notech_nor2 i_221(.A(n_2603), .B(n_60221), .Z(n_44531));
	notech_nor2 i_222(.A(n_2611), .B(n_60221), .Z(n_44537));
	notech_nor2 i_223(.A(n_2619), .B(n_60221), .Z(n_44543));
	notech_nor2 i_224(.A(n_2627), .B(n_60221), .Z(n_44549));
	notech_nor2 i_225(.A(n_2635), .B(n_60221), .Z(n_44555));
	notech_nor2 i_226(.A(n_2643), .B(n_60221), .Z(n_44561));
	notech_nor2 i_227(.A(n_3236), .B(n_43905), .Z(n_44567));
	notech_nor2 i_228(.A(n_3236), .B(n_43903), .Z(n_44573));
	notech_nor2 i_229(.A(n_3236), .B(n_43899), .Z(n_44579));
	notech_nor2 i_230(.A(n_3236), .B(n_43897), .Z(n_44585));
	notech_nor2 i_231(.A(n_3236), .B(n_43893), .Z(n_44591));
	notech_nor2 i_232(.A(n_55701), .B(n_43887), .Z(n_44597));
	notech_nor2 i_234(.A(n_55701), .B(n_43879), .Z(n_44609));
	notech_nor2 i_235(.A(n_3246), .B(n_43861), .Z(n_44615));
	notech_nor2 i_236(.A(n_3246), .B(n_43857), .Z(n_44621));
	notech_nor2 i_237(.A(n_3246), .B(n_43855), .Z(n_44627));
	notech_nor2 i_238(.A(n_3246), .B(n_43851), .Z(n_44633));
	notech_nor2 i_239(.A(n_55762), .B(n_43849), .Z(n_44639));
	notech_nor2 i_240(.A(n_55762), .B(n_43845), .Z(n_44645));
	notech_nor2 i_241(.A(n_55762), .B(n_43841), .Z(n_44651));
	notech_nor2 i_242(.A(n_55762), .B(n_43838), .Z(n_44657));
	notech_nor2 i_418(.A(n_5745), .B(n_1898), .Z(n_1892));
	notech_nor2 i_67(.A(twobyte), .B(fpu), .Z(n_5745));
	notech_and2 i_95611435(.A(\to_acu2_0[0] ), .B(\to_acu2_0[1] ), .Z(n_5712
		));
	notech_nand2 i_65686(.A(n_2967), .B(n_2964), .Z(n_1879));
	notech_and2 i_65692(.A(n_44683), .B(n_44682), .Z(n_1878));
	notech_nor2 i_233(.A(n_55701), .B(n_43832), .Z(n_44603));
	notech_ao3 i_3439(.A(n_60905), .B(udeco[127]), .C(n_60346), .Z(n_42642)
		);
	notech_ao3 i_3438(.A(n_60904), .B(udeco[126]), .C(n_60348), .Z(n_42636)
		);
	notech_ao3 i_3436(.A(n_60904), .B(udeco[124]), .C(n_60348), .Z(n_42624)
		);
	notech_ao3 i_3434(.A(n_60904), .B(udeco[122]), .C(n_60348), .Z(n_42612)
		);
	notech_ao3 i_3432(.A(n_60904), .B(udeco[120]), .C(n_60348), .Z(n_42600)
		);
	notech_ao3 i_3430(.A(n_60904), .B(udeco[118]), .C(n_60348), .Z(n_42588)
		);
	notech_ao3 i_3427(.A(n_60904), .B(udeco[115]), .C(n_60348), .Z(n_42570)
		);
	notech_ao3 i_3426(.A(n_60904), .B(udeco[114]), .C(n_60346), .Z(n_42564)
		);
	notech_ao3 i_3425(.A(n_60904), .B(udeco[113]), .C(n_60346), .Z(n_42558)
		);
	notech_ao3 i_3419(.A(n_60905), .B(udeco[107]), .C(n_60346), .Z(n_42522)
		);
	notech_ao3 i_112(.A(n_60904), .B(udeco[103]), .C(n_60348), .Z(n_42498)
		);
	notech_ao3 i_3413(.A(n_60904), .B(udeco[101]), .C(n_60348), .Z(n_42486)
		);
	notech_ao3 i_3407(.A(n_60904), .B(udeco[95]), .C(n_60346), .Z(n_42450)
		);
	notech_ao3 i_3406(.A(n_60837), .B(udeco[94]), .C(n_60362), .Z(n_42444)
		);
	notech_ao3 i_3405(.A(n_60837), .B(udeco[93]), .C(n_60361), .Z(n_42438)
		);
	notech_ao3 i_3404(.A(n_60837), .B(udeco[92]), .C(n_60362), .Z(n_42432)
		);
	notech_ao3 i_3403(.A(n_60837), .B(udeco[91]), .C(n_60362), .Z(n_42426)
		);
	notech_ao3 i_3402(.A(n_60837), .B(udeco[90]), .C(n_60362), .Z(n_42420)
		);
	notech_ao3 i_3401(.A(n_60837), .B(udeco[89]), .C(n_60361), .Z(n_42414)
		);
	notech_ao3 i_3400(.A(n_60837), .B(udeco[88]), .C(n_60361), .Z(n_42408)
		);
	notech_ao3 i_3399(.A(n_60837), .B(udeco[87]), .C(n_60361), .Z(n_42402)
		);
	notech_ao3 i_3398(.A(n_60837), .B(udeco[86]), .C(n_60361), .Z(n_42396)
		);
	notech_ao3 i_3397(.A(n_60837), .B(udeco[85]), .C(n_60361), .Z(n_42390)
		);
	notech_ao4 i_1226117(.A(n_60221), .B(n_44727), .C(n_59185), .D(n_43494),
		 .Z(n_3332));
	notech_ao3 i_25980643(.A(n_60837), .B(\to_acu2_0[11] ), .C(n_60361), .Z(n_3331
		));
	notech_ao3 i_130(.A(udeco[103]), .B(rep), .C(n_60221), .Z(n_49797));
	notech_nor2 i_131(.A(n_60227), .B(n_43466), .Z(n_45639));
	notech_ao4 i_1326118(.A(n_60232), .B(n_44716), .C(n_59185), .D(n_43495),
		 .Z(n_3330));
	notech_nor2 i_3730155(.A(int_excl[2]), .B(n_1734), .Z(n_1755));
	notech_or4 i_3830156(.A(int_excl[1]), .B(int_excl[0]), .C(int_excl[2]), 
		.D(int_excl[3]), .Z(n_1754));
	notech_nor2 i_1398051(.A(n_2994), .B(pc_req), .Z(n_41609));
	notech_nao3 i_27(.A(db67), .B(n_60837), .C(n_2994), .Z(n_5721));
	notech_ao3 i_28080644(.A(n_60836), .B(\to_acu2_0[12] ), .C(n_60361), .Z(n_3329
		));
	notech_nand2 i_31(.A(n_2339), .B(n_44684), .Z(n_1744));
	notech_or2 i_60(.A(int_excl[1]), .B(int_excl[0]), .Z(n_1734));
	notech_and2 i_63(.A(n_3007), .B(n_44747), .Z(n_1733));
	notech_or2 i_73(.A(int_excl[4]), .B(n_1754), .Z(n_1730));
	notech_nand2 i_94(.A(n_2342), .B(n_2341), .Z(n_1724));
	notech_ao4 i_1426119(.A(n_60232), .B(n_44713), .C(n_59184), .D(n_43497),
		 .Z(n_3328));
	notech_nand3 i_128(.A(n_60361), .B(n_2975), .C(n_60836), .Z(n_1714));
	notech_or4 i_6244(.A(fsm[2]), .B(n_2969), .C(fsm[0]), .D(n_43437), .Z(n_5770
		));
	notech_ao3 i_39580645(.A(n_60836), .B(\to_acu2_0[13] ), .C(n_60346), .Z(n_3327
		));
	notech_ao4 i_1526120(.A(n_60232), .B(n_44712), .C(n_59184), .D(n_43499),
		 .Z(n_3326));
	notech_ao3 i_25880646(.A(n_60836), .B(\to_acu2_0[14] ), .C(n_60346), .Z(n_3325
		));
	notech_ao4 i_1626121(.A(n_60232), .B(n_44711), .C(n_59184), .D(n_43501),
		 .Z(n_3324));
	notech_ao3 i_25780647(.A(n_60836), .B(\to_acu2_0[15] ), .C(n_60346), .Z(n_3323
		));
	notech_ao4 i_1726122(.A(n_60232), .B(n_44718), .C(n_59185), .D(n_43502),
		 .Z(n_3322));
	notech_ao3 i_33480648(.A(n_60836), .B(\to_acu2_0[16] ), .C(n_60361), .Z(n_3321
		));
	notech_ao4 i_1826123(.A(n_60232), .B(n_44715), .C(n_59185), .D(n_43505),
		 .Z(n_3320));
	notech_ao3 i_25680649(.A(n_60836), .B(\to_acu2_0[17] ), .C(n_60362), .Z(n_3319
		));
	notech_ao4 i_1926124(.A(n_60230), .B(n_44714), .C(n_59185), .D(n_43506),
		 .Z(n_3318));
	notech_ao3 i_25580650(.A(n_60836), .B(\to_acu2_0[18] ), .C(n_60362), .Z(n_3317
		));
	notech_ao4 i_5526160(.A(n_60232), .B(n_44732), .C(n_59185), .D(n_43560),
		 .Z(n_3316));
	notech_ao4 i_8526190(.A(n_60232), .B(n_44736), .C(n_59185), .D(n_43597),
		 .Z(n_3315));
	notech_ao4 i_17926284(.A(n_60232), .B(n_44619), .C(n_59185), .D(n_43782)
		, .Z(n_3314));
	notech_ao3 i_15880651(.A(n_60836), .B(in128[95]), .C(n_60361), .Z(n_3313
		));
	notech_ao4 i_18026285(.A(n_60236), .B(n_44620), .C(n_59185), .D(n_43783)
		, .Z(n_3312));
	notech_ao3 i_15980652(.A(n_60836), .B(in128[96]), .C(n_60361), .Z(n_3311
		));
	notech_ao4 i_18126286(.A(n_60236), .B(n_44622), .C(n_59185), .D(n_43784)
		, .Z(n_3310));
	notech_ao3 i_16080653(.A(n_60836), .B(in128[97]), .C(n_60361), .Z(n_3309
		));
	notech_ao4 i_18226287(.A(n_60236), .B(n_44623), .C(n_59185), .D(n_43785)
		, .Z(n_3308));
	notech_ao3 i_16180654(.A(n_60836), .B(in128[98]), .C(n_60348), .Z(n_3307
		));
	notech_ao4 i_18326288(.A(n_60236), .B(n_44624), .C(n_59185), .D(n_43788)
		, .Z(n_3306));
	notech_or2 i_080662(.A(n_60339), .B(pc_req), .Z(n_5769));
	notech_ao3 i_16280655(.A(n_60836), .B(in128[99]), .C(n_60339), .Z(n_3305
		));
	notech_ao4 i_21126316(.A(n_60236), .B(n_44658), .C(n_59185), .D(n_43825)
		, .Z(n_3304));
	notech_nao3 i_6241(.A(n_2380), .B(n_44729), .C(twobyte), .Z(n_1676));
	notech_nand3 i_10380656(.A(n_5745), .B(n_2379), .C(n_2380), .Z(n_17054783
		));
	notech_and2 i_12780657(.A(n_1600), .B(n_1813), .Z(n_3303));
	notech_and3 i_4780658(.A(n_60934), .B(n_5767), .C(n_2402), .Z(n_5765));
	notech_and3 i_7580660(.A(n_60932), .B(n_194199020), .C(n_1600), .Z(n_3302
		));
	notech_and3 i_72449(.A(n_1600), .B(n_1813), .C(n_1533), .Z(n_3301));
	notech_and2 i_74312(.A(n_5765), .B(n_1601), .Z(n_3300));
	notech_and4 i_75510(.A(n_1813), .B(n_1812), .C(n_1817), .D(n_1800), .Z(n_3299
		));
	notech_and2 i_70766(.A(n_5765), .B(n_1604), .Z(n_3298));
	notech_and2 i_72060(.A(n_60932), .B(n_2387), .Z(n_3297));
	notech_ao3 i_70704(.A(n_5765), .B(n_2381), .C(n_1605), .Z(n_3296));
	notech_ao3 i_70920(.A(n_5765), .B(n_44369), .C(n_1803), .Z(n_3295));
	notech_ao3 i_71390(.A(n_5765), .B(n_2386), .C(n_1605), .Z(n_3294));
	notech_nor2 i_73501(.A(n_1606), .B(n_1607), .Z(n_3293));
	notech_and2 i_70750(.A(n_5765), .B(n_43787), .Z(n_3292));
	notech_nand3 i_1225(.A(n_2336), .B(n_2998), .C(n_3020), .Z(n_3289));
	notech_ao4 i_1219(.A(ipg_fault), .B(n_43465), .C(pc_req), .D(n_3017), .Z
		(n_3288));
	notech_ao4 i_1183(.A(n_2866), .B(n_44729), .C(n_2865), .D(n_43465), .Z(n_3284
		));
	notech_or4 i_1176(.A(\fpu_indrm[3] ), .B(\fpu_indrm[2] ), .C(\fpu_indrm[4] 
		), .D(n_2412), .Z(n_3283));
	notech_nao3 i_1169(.A(n_3280), .B(n_43797), .C(n_2845), .Z(n_3281));
	notech_ao4 i_99(.A(n_43827), .B(n_3279), .C(n_3256), .D(n_3278), .Z(n_3280
		));
	notech_nand3 i_1163(.A(n_2859), .B(n_5712), .C(n_44751), .Z(n_3279));
	notech_nao3 i_1161(.A(n_2859), .B(\to_acu2_0[4] ), .C(n_3015), .Z(n_3278
		));
	notech_ao4 i_1155(.A(n_43827), .B(n_3271), .C(n_2850), .D(n_43814), .Z(n_3272
		));
	notech_nand3 i_1154(.A(n_2859), .B(n_5712), .C(\to_acu2_0[4] ), .Z(n_3271
		));
	notech_ao3 i_37(.A(n_2859), .B(n_42548), .C(n_43827), .Z(n_3270));
	notech_and4 i_70(.A(db67), .B(n_3014), .C(n_41609), .D(n_44729), .Z(n_3266
		));
	notech_or4 i_118(.A(n_3256), .B(\to_acu2_0[4] ), .C(\to_acu2_0[3] ), .D(n_3015
		), .Z(n_3263));
	notech_ao4 i_945(.A(n_2706), .B(in128[46]), .C(n_2705), .D(in128[54]), .Z
		(n_3260));
	notech_or4 i_933(.A(\fpu_indrm[3] ), .B(\fpu_indrm[2] ), .C(n_2412), .D(n_42645
		), .Z(n_3258));
	notech_or2 i_48(.A(db67), .B(n_43465), .Z(n_3256));
	notech_ao4 i_893(.A(n_2692), .B(in128[55]), .C(n_2705), .D(in128[63]), .Z
		(n_3254));
	notech_ao4 i_888(.A(n_2689), .B(in128[54]), .C(n_2705), .D(in128[62]), .Z
		(n_3253));
	notech_ao4 i_883(.A(n_2686), .B(in128[53]), .C(n_2705), .D(in128[61]), .Z
		(n_3252));
	notech_ao4 i_878(.A(n_2683), .B(in128[52]), .C(n_2705), .D(in128[60]), .Z
		(n_3251));
	notech_ao4 i_873(.A(n_2680), .B(in128[51]), .C(n_2705), .D(in128[59]), .Z
		(n_3250));
	notech_ao4 i_868(.A(n_2677), .B(in128[50]), .C(n_2705), .D(in128[58]), .Z
		(n_3249));
	notech_ao4 i_863(.A(n_2674), .B(in128[49]), .C(n_2705), .D(in128[57]), .Z
		(n_3248));
	notech_ao4 i_858(.A(n_2671), .B(in128[48]), .C(n_2705), .D(in128[56]), .Z
		(n_3247));
	notech_nao3 i_7(.A(n_60837), .B(n_2670), .C(n_60339), .Z(n_3246));
	notech_and4 i_87(.A(n_3118), .B(n_3197), .C(n_3061), .D(n_3076), .Z(n_3245
		));
	notech_ao4 i_851(.A(n_2667), .B(in128[47]), .C(n_2705), .D(in128[55]), .Z
		(n_3243));
	notech_ao4 i_846(.A(n_2664), .B(in128[45]), .C(n_2705), .D(in128[53]), .Z
		(n_3242));
	notech_ao4 i_841(.A(n_2661), .B(in128[44]), .C(n_2705), .D(in128[52]), .Z
		(n_3241));
	notech_ao4 i_836(.A(n_2658), .B(in128[43]), .C(n_2705), .D(in128[51]), .Z
		(n_3240));
	notech_ao4 i_831(.A(n_2655), .B(in128[42]), .C(n_2705), .D(in128[50]), .Z
		(n_3239));
	notech_ao4 i_826(.A(n_2652), .B(in128[41]), .C(n_2705), .D(in128[49]), .Z
		(n_3238));
	notech_ao4 i_821(.A(n_2649), .B(in128[40]), .C(n_2705), .D(in128[48]), .Z
		(n_3237));
	notech_nao3 i_2(.A(n_60847), .B(n_2648), .C(n_60339), .Z(n_3236));
	notech_and4 i_89(.A(n_3061), .B(n_3118), .C(n_3076), .D(n_43910), .Z(n_3235
		));
	notech_ao4 i_812(.A(n_3164), .B(n_44590), .C(n_3163), .D(n_44610), .Z(n_3232
		));
	notech_and2 i_807(.A(n_2642), .B(n_3229), .Z(n_3230));
	notech_ao4 i_806(.A(n_3157), .B(n_44600), .C(n_3156), .D(n_44581), .Z(n_3229
		));
	notech_ao4 i_799(.A(n_3164), .B(n_44589), .C(n_3163), .D(n_44608), .Z(n_3227
		));
	notech_and2 i_794(.A(n_2634), .B(n_3224), .Z(n_3225));
	notech_ao4 i_793(.A(n_3157), .B(n_44599), .C(n_3156), .D(n_44580), .Z(n_3224
		));
	notech_ao4 i_786(.A(n_3164), .B(n_44588), .C(n_3163), .D(n_44607), .Z(n_3222
		));
	notech_and2 i_781(.A(n_2626), .B(n_3219), .Z(n_3220));
	notech_ao4 i_780(.A(n_3157), .B(n_44598), .C(n_3156), .D(n_44578), .Z(n_3219
		));
	notech_ao4 i_773(.A(n_3164), .B(n_44587), .C(n_3163), .D(n_44606), .Z(n_3217
		));
	notech_and2 i_768(.A(n_2618), .B(n_3214), .Z(n_3215));
	notech_ao4 i_767(.A(n_3157), .B(n_44596), .C(n_3156), .D(n_44577), .Z(n_3214
		));
	notech_ao4 i_760(.A(n_3164), .B(n_44586), .C(n_3163), .D(n_44605), .Z(n_3212
		));
	notech_and2 i_755(.A(n_2610), .B(n_3209), .Z(n_3210));
	notech_ao4 i_754(.A(n_3157), .B(n_44595), .C(n_3156), .D(n_44576), .Z(n_3209
		));
	notech_ao4 i_747(.A(n_3164), .B(n_44584), .C(n_3163), .D(n_44604), .Z(n_3207
		));
	notech_and2 i_742(.A(n_2602), .B(n_3204), .Z(n_3205));
	notech_ao4 i_741(.A(n_3157), .B(n_44594), .C(n_3156), .D(n_44575), .Z(n_3204
		));
	notech_ao4 i_734(.A(n_3164), .B(n_44582), .C(n_3163), .D(n_44601), .Z(n_3202
		));
	notech_and2 i_729(.A(n_2594), .B(n_3199), .Z(n_3200));
	notech_ao4 i_728(.A(n_3157), .B(n_44592), .C(n_3156), .D(n_44572), .Z(n_3199
		));
	notech_or2 i_88(.A(n_3158), .B(n_2590), .Z(n_3198));
	notech_mux2 i_81(.S(imm_sz[1]), .A(n_44371), .B(imm_sz[2]), .Z(n_3197)
		);
	notech_ao4 i_718(.A(n_3164), .B(n_44581), .C(n_3163), .D(n_44600), .Z(n_3195
		));
	notech_and2 i_713(.A(n_2584), .B(n_3192), .Z(n_3193));
	notech_ao4 i_712(.A(n_3158), .B(n_44552), .C(n_3157), .D(n_44590), .Z(n_3192
		));
	notech_ao4 i_705(.A(n_3164), .B(n_44580), .C(n_3163), .D(n_44599), .Z(n_3190
		));
	notech_and2 i_700(.A(n_2576), .B(n_3187), .Z(n_3188));
	notech_ao4 i_699(.A(n_3158), .B(n_44551), .C(n_3157), .D(n_44589), .Z(n_3187
		));
	notech_ao4 i_692(.A(n_3164), .B(n_44577), .C(n_3163), .D(n_44596), .Z(n_3185
		));
	notech_and2 i_687(.A(n_2568), .B(n_3182), .Z(n_3183));
	notech_ao4 i_686(.A(n_3158), .B(n_44548), .C(n_3157), .D(n_44587), .Z(n_3182
		));
	notech_ao4 i_679(.A(n_3164), .B(n_44576), .C(n_3163), .D(n_44595), .Z(n_3180
		));
	notech_and2 i_674(.A(n_2560), .B(n_3177), .Z(n_3178));
	notech_ao4 i_673(.A(n_3158), .B(n_44547), .C(n_3157), .D(n_44586), .Z(n_3177
		));
	notech_ao4 i_666(.A(n_3164), .B(n_44575), .C(n_3163), .D(n_44594), .Z(n_3175
		));
	notech_and2 i_661(.A(n_2552), .B(n_3172), .Z(n_3173));
	notech_ao4 i_660(.A(n_3158), .B(n_44546), .C(n_3157), .D(n_44584), .Z(n_3172
		));
	notech_ao4 i_653(.A(n_3164), .B(n_44574), .C(n_3163), .D(n_44593), .Z(n_3170
		));
	notech_and2 i_648(.A(n_2544), .B(n_3167), .Z(n_3168));
	notech_ao4 i_647(.A(n_3158), .B(n_44545), .C(n_3157), .D(n_44583), .Z(n_3167
		));
	notech_ao4 i_640(.A(n_3164), .B(n_44572), .C(n_3163), .D(n_44592), .Z(n_3165
		));
	notech_or4 i_52(.A(imm_sz[0]), .B(imm_sz[1]), .C(n_3060), .D(n_44158), .Z
		(n_3164));
	notech_nand2 i_51(.A(n_3117), .B(n_44159), .Z(n_3163));
	notech_nao3 i_50(.A(n_3060), .B(n_2531), .C(n_44158), .Z(n_3162));
	notech_and2 i_635(.A(n_2536), .B(n_3159), .Z(n_3160));
	notech_ao4 i_634(.A(n_3158), .B(n_44544), .C(n_3157), .D(n_44582), .Z(n_3159
		));
	notech_or4 i_91(.A(n_3068), .B(n_2532), .C(n_2418), .D(n_2417), .Z(n_3158
		));
	notech_or4 i_55(.A(imm_sz[0]), .B(imm_sz[1]), .C(n_3060), .D(n_3068), .Z
		(n_3157));
	notech_nao3 i_53(.A(n_3057), .B(n_3117), .C(n_3064), .Z(n_3156));
	notech_or4 i_59(.A(imm_sz[0]), .B(imm_sz[1]), .C(n_3057), .D(n_3064), .Z
		(n_3155));
	notech_ao4 i_625(.A(n_44542), .B(n_3132), .C(n_3130), .D(n_44581), .Z(n_3153
		));
	notech_and2 i_620(.A(n_3150), .B(n_2526), .Z(n_3151));
	notech_ao4 i_619(.A(n_3125), .B(n_44571), .C(n_3124), .D(n_44590), .Z(n_3150
		));
	notech_ao4 i_612(.A(n_3132), .B(n_44539), .C(n_3130), .D(n_44577), .Z(n_3148
		));
	notech_and2 i_607(.A(n_3145), .B(n_2518), .Z(n_3146));
	notech_ao4 i_606(.A(n_3125), .B(n_44568), .C(n_3124), .D(n_44587), .Z(n_3145
		));
	notech_ao4 i_599(.A(n_3132), .B(n_44538), .C(n_3130), .D(n_44576), .Z(n_3143
		));
	notech_and2 i_594(.A(n_3140), .B(n_2510), .Z(n_3141));
	notech_ao4 i_593(.A(n_3125), .B(n_44566), .C(n_3124), .D(n_44586), .Z(n_3140
		));
	notech_ao4 i_586(.A(n_3132), .B(n_44536), .C(n_3130), .D(n_44575), .Z(n_3138
		));
	notech_and2 i_581(.A(n_3135), .B(n_2502), .Z(n_3136));
	notech_ao4 i_580(.A(n_3125), .B(n_44565), .C(n_3124), .D(n_44584), .Z(n_3135
		));
	notech_ao4 i_573(.A(n_3132), .B(n_44534), .C(n_3130), .D(n_44572), .Z(n_3133
		));
	notech_nao3 i_82(.A(n_3060), .B(n_2488), .C(n_3068), .Z(n_3132));
	notech_ao3 i_46(.A(n_2490), .B(n_3061), .C(n_3117), .Z(n_3131));
	notech_or2 i_84(.A(n_3118), .B(n_3069), .Z(n_3130));
	notech_or4 i_83(.A(n_2420), .B(n_2419), .C(n_3064), .D(n_3118), .Z(n_3129
		));
	notech_and2 i_568(.A(n_3126), .B(n_2494), .Z(n_3127));
	notech_ao4 i_567(.A(n_3125), .B(n_44563), .C(n_3124), .D(n_44582), .Z(n_3126
		));
	notech_or2 i_90(.A(n_3118), .B(n_3078), .Z(n_3125));
	notech_or2 i_85(.A(n_3118), .B(n_3072), .Z(n_3124));
	notech_nao3 i_92(.A(n_3060), .B(n_2489), .C(n_44158), .Z(n_3123));
	notech_nand3 i_830111(.A(imm_sz[1]), .B(n_44371), .C(imm_sz[2]), .Z(n_3121
		));
	notech_or2 i_86(.A(n_3118), .B(n_3065), .Z(n_3119));
	notech_and2 i_4(.A(n_2490), .B(n_44105), .Z(n_3118));
	notech_nor2 i_630108(.A(imm_sz[1]), .B(imm_sz[0]), .Z(n_3117));
	notech_ao4 i_554(.A(n_44157), .B(n_44719), .C(n_3078), .D(n_44562), .Z(n_3115
		));
	notech_and2 i_549(.A(n_3112), .B(n_2483), .Z(n_3113));
	notech_ao4 i_548(.A(n_3072), .B(n_44581), .C(n_3069), .D(n_44571), .Z(n_3112
		));
	notech_ao4 i_541(.A(n_44157), .B(n_44721), .C(n_44560), .D(n_3078), .Z(n_3110
		));
	notech_and2 i_536(.A(n_3107), .B(n_2475), .Z(n_3108));
	notech_ao4 i_535(.A(n_3072), .B(n_44580), .C(n_44570), .D(n_3069), .Z(n_3107
		));
	notech_ao4 i_528(.A(n_44157), .B(n_44708), .C(n_3078), .D(n_44559), .Z(n_3105
		));
	notech_and2 i_523(.A(n_3102), .B(n_2467), .Z(n_3103));
	notech_ao4 i_522(.A(n_3072), .B(n_44578), .C(n_3069), .D(n_44569), .Z(n_3102
		));
	notech_ao4 i_515(.A(n_44157), .B(n_44709), .C(n_3078), .D(n_44558), .Z(n_3100
		));
	notech_and2 i_510(.A(n_3097), .B(n_2459), .Z(n_3098));
	notech_ao4 i_509(.A(n_3072), .B(n_44577), .C(n_3069), .D(n_44568), .Z(n_3097
		));
	notech_ao3 i_26080642(.A(n_60847), .B(\to_acu2_0[10] ), .C(n_60339), .Z(n_11899519
		));
	notech_nao3 i_30280355(.A(cpl[0]), .B(cpl[1]), .C(n_59157), .Z(n_13699537
		));
	notech_nao3 i_39180269(.A(n_2379), .B(\to_acu2_0[71] ), .C(n_1676), .Z(n_16599551
		));
	notech_nao3 i_39380267(.A(idx_deco[0]), .B(n_43434), .C(n_5767), .Z(n_16799552
		));
	notech_nao3 i_126079401(.A(n_2379), .B(\to_acu2_0[75] ), .C(n_1676), .Z(n_1097100405
		));
	notech_nao3 i_126179400(.A(n_2379), .B(\to_acu2_0[70] ), .C(n_1676), .Z(n_1098100406
		));
	notech_and3 i_279298191(.A(n_2382), .B(to_acu1[39]), .C(n_60847), .Z(n_1099100407
		));
	notech_nand3 i_28180376(.A(n_2995), .B(inst_deco1[113]), .C(n_59410), .Z
		(n_1178100486));
	notech_and2 i_293298192(.A(lenpc1[6]), .B(n_59410), .Z(n_1181100489));
	notech_and2 i_293398193(.A(lenpc1[7]), .B(n_59410), .Z(n_1182100490));
	notech_and2 i_293498194(.A(lenpc1[8]), .B(n_59410), .Z(n_1183100491));
	notech_and2 i_293598195(.A(lenpc1[9]), .B(n_59410), .Z(n_1184100492));
	notech_and2 i_293698196(.A(lenpc1[10]), .B(n_59410), .Z(n_1185100493));
	notech_and2 i_293798197(.A(lenpc1[11]), .B(n_59410), .Z(n_1186100494));
	notech_and2 i_293898198(.A(lenpc1[12]), .B(n_59410), .Z(n_1187100495));
	notech_and2 i_293998199(.A(lenpc1[13]), .B(n_59410), .Z(n_1188100496));
	notech_and2 i_294098200(.A(lenpc1[14]), .B(n_59410), .Z(n_1189100497));
	notech_and2 i_294198201(.A(lenpc1[15]), .B(n_59410), .Z(n_1190100498));
	notech_and2 i_294298202(.A(lenpc1[16]), .B(n_59410), .Z(n_1191100499));
	notech_and2 i_294398203(.A(lenpc1[17]), .B(n_59410), .Z(n_1192100500));
	notech_and2 i_294498204(.A(lenpc1[18]), .B(n_59410), .Z(n_1193100501));
	notech_and2 i_294698205(.A(lenpc1[20]), .B(n_59410), .Z(n_1194100502));
	notech_and3 i_298398206(.A(n_2382), .B(lenpc2[31]), .C(n_60831), .Z(n_1195100503
		));
	notech_and3 i_299798207(.A(n_2382), .B(to_acu2[39]), .C(n_60831), .Z(n_1196100504
		));
	notech_ao4 i_138679275(.A(n_60122), .B(n_44505), .C(n_1912), .D(n_42555)
		, .Z(n_1198100506));
	notech_ao4 i_133679325(.A(n_59150), .B(n_43259), .C(n_60122), .D(n_44460
		), .Z(n_1200100508));
	notech_ao4 i_132679335(.A(n_59150), .B(n_43235), .C(n_60122), .D(n_44450
		), .Z(n_1201100509));
	notech_ao4 i_132579336(.A(n_59150), .B(n_43232), .C(n_60122), .D(n_44449
		), .Z(n_1202100510));
	notech_ao4 i_132479337(.A(n_59150), .B(n_43230), .C(n_60122), .D(n_44448
		), .Z(n_1204100511));
	notech_ao4 i_132379338(.A(n_59150), .B(n_43227), .C(n_60122), .D(n_44446
		), .Z(n_1205100512));
	notech_ao4 i_132279339(.A(n_59150), .B(n_43225), .C(n_60122), .D(n_44445
		), .Z(n_1206100513));
	notech_ao4 i_132179340(.A(n_59150), .B(n_43223), .C(n_60122), .D(n_44444
		), .Z(n_1207100514));
	notech_ao4 i_131979342(.A(n_59151), .B(n_43218), .C(n_60122), .D(n_44442
		), .Z(n_1208100515));
	notech_ao4 i_131879343(.A(n_59151), .B(n_43215), .C(n_60122), .D(n_44440
		), .Z(n_1209100516));
	notech_ao4 i_131679345(.A(n_59151), .B(n_43211), .C(n_60122), .D(n_44438
		), .Z(n_1210100517));
	notech_ao4 i_131579346(.A(n_59150), .B(n_43208), .C(n_60122), .D(n_44437
		), .Z(n_1211100518));
	notech_ao4 i_131479347(.A(n_59150), .B(n_43206), .C(n_60122), .D(n_44436
		), .Z(n_1212100519));
	notech_ao4 i_131379348(.A(n_59150), .B(n_43203), .C(n_60122), .D(n_44434
		), .Z(n_1213100520));
	notech_ao4 i_131179350(.A(n_59150), .B(n_43199), .C(n_60122), .D(n_44432
		), .Z(n_1214100521));
	notech_ao4 i_131079351(.A(n_59150), .B(n_43196), .C(n_60122), .D(n_44431
		), .Z(n_1215100522));
	notech_ao4 i_130779354(.A(n_59146), .B(n_43189), .C(n_60120), .D(n_44428
		), .Z(n_1216100523));
	notech_ao4 i_130679355(.A(n_59146), .B(n_43187), .C(n_60120), .D(n_44427
		), .Z(n_1217100524));
	notech_ao4 i_130479357(.A(n_59146), .B(n_43181), .C(n_60120), .D(n_44425
		), .Z(n_1218100525));
	notech_ao4 i_130379358(.A(n_59146), .B(n_43177), .C(n_60120), .D(n_44424
		), .Z(n_1219100526));
	notech_ao4 i_130279359(.A(n_59146), .B(n_43175), .C(n_60120), .D(n_44422
		), .Z(n_1220100527));
	notech_ao4 i_130179360(.A(n_59146), .B(n_43172), .C(n_60120), .D(n_44421
		), .Z(n_1221100528));
	notech_ao4 i_130079361(.A(n_59146), .B(n_43170), .C(n_60120), .D(n_44420
		), .Z(n_1222100529));
	notech_ao4 i_129879363(.A(n_59150), .B(n_43165), .C(n_60120), .D(n_44418
		), .Z(n_1223100530));
	notech_ao4 i_129779364(.A(n_59150), .B(n_43163), .C(n_60120), .D(n_44416
		), .Z(n_1224100531));
	notech_ao4 i_129679365(.A(n_59150), .B(n_43160), .C(n_60120), .D(n_44415
		), .Z(n_1225100532));
	notech_ao4 i_129579366(.A(n_59150), .B(n_43158), .C(n_60120), .D(n_44414
		), .Z(n_1226100533));
	notech_ao4 i_129379368(.A(n_59146), .B(n_43153), .C(n_60120), .D(n_44412
		), .Z(n_1227100534));
	notech_ao4 i_128579376(.A(n_59146), .B(n_43134), .C(n_60120), .D(n_44402
		), .Z(n_1228100535));
	notech_ao4 i_128479377(.A(n_59146), .B(n_43131), .C(n_60120), .D(n_44401
		), .Z(n_1229100536));
	notech_ao4 i_128279379(.A(n_59153), .B(n_43125), .C(n_60120), .D(n_44397
		), .Z(n_1230100537));
	notech_ao4 i_128179380(.A(n_59153), .B(n_43123), .C(n_60120), .D(n_44396
		), .Z(n_1231100538));
	notech_ao4 i_128079381(.A(n_59153), .B(n_43119), .C(n_60127), .D(n_44394
		), .Z(n_1232100539));
	notech_ao4 i_127879383(.A(n_59153), .B(n_43115), .C(n_60127), .D(n_44391
		), .Z(n_1233100540));
	notech_ao4 i_127779384(.A(n_59153), .B(n_43112), .C(n_60127), .D(n_44390
		), .Z(n_1234100541));
	notech_ao4 i_127679385(.A(n_59153), .B(n_43110), .C(n_60127), .D(n_44389
		), .Z(n_1235100542));
	notech_ao4 i_127579386(.A(n_59153), .B(n_43107), .C(n_60127), .D(n_44388
		), .Z(n_1236100543));
	notech_ao4 i_127479387(.A(n_59153), .B(n_43105), .C(n_60127), .D(n_44386
		), .Z(n_1237100544));
	notech_ao4 i_127379388(.A(n_59153), .B(n_43103), .C(n_60127), .D(n_44385
		), .Z(n_1238100545));
	notech_ao4 i_127279389(.A(n_59153), .B(n_43100), .C(n_60127), .D(n_44384
		), .Z(n_1239100546));
	notech_or4 i_66520(.A(trig_it), .B(intff), .C(n_43379), .D(n_44768), .Z(n_1240100547
		));
	notech_nand3 i_22778822(.A(n_1553100858), .B(n_1552100857), .C(n_1478100784
		), .Z(n_1241100548));
	notech_ao4 i_3279009(.A(n_2413), .B(n_42721), .C(n_5745), .D(n_1898), .Z
		(n_1477100783));
	notech_nand2 i_77578274(.A(n_2847), .B(fpu), .Z(n_1478100784));
	notech_nao3 i_79178258(.A(idx_deco[1]), .B(n_43431), .C(n_5767), .Z(n_1481100787
		));
	notech_and2 i_294798208(.A(lenpc1[21]), .B(n_59410), .Z(n_1482100788));
	notech_and2 i_294898209(.A(lenpc1[22]), .B(n_59410), .Z(n_1483100789));
	notech_and2 i_294998210(.A(lenpc1[23]), .B(n_59410), .Z(n_1484100790));
	notech_and2 i_295098211(.A(lenpc1[24]), .B(n_59410), .Z(n_1485100791));
	notech_and2 i_295198212(.A(lenpc1[25]), .B(n_59405), .Z(n_1486100792));
	notech_and2 i_295298213(.A(lenpc1[26]), .B(n_59405), .Z(n_1487100793));
	notech_and2 i_295398214(.A(lenpc1[27]), .B(n_59405), .Z(n_1488100794));
	notech_and2 i_295498215(.A(lenpc1[28]), .B(n_59405), .Z(n_1489100795));
	notech_and2 i_295598216(.A(lenpc1[29]), .B(n_59405), .Z(n_1490100796));
	notech_and2 i_295698217(.A(lenpc1[30]), .B(n_59405), .Z(n_1491100797));
	notech_and2 i_295798218(.A(lenpc1[31]), .B(n_59405), .Z(n_1492100798));
	notech_and3 i_295898219(.A(lenpc2[6]), .B(n_2382), .C(n_60847), .Z(n_1493100799
		));
	notech_and3 i_296098220(.A(n_2382), .B(lenpc2[8]), .C(n_60847), .Z(n_1494100800
		));
	notech_and3 i_296198221(.A(n_2382), .B(lenpc2[9]), .C(n_60847), .Z(n_1495100801
		));
	notech_and3 i_296398222(.A(n_2382), .B(lenpc2[11]), .C(n_60847), .Z(n_1496100802
		));
	notech_and3 i_296498223(.A(n_2382), .B(lenpc2[12]), .C(n_60847), .Z(n_1497100803
		));
	notech_and3 i_296598224(.A(n_2382), .B(lenpc2[13]), .C(n_60847), .Z(n_1498100804
		));
	notech_and3 i_296698225(.A(n_2382), .B(lenpc2[14]), .C(n_60847), .Z(n_1499100805
		));
	notech_and3 i_296798226(.A(n_2382), .B(lenpc2[15]), .C(n_60831), .Z(n_1500100806
		));
	notech_and3 i_296898227(.A(n_2382), .B(lenpc2[16]), .C(n_60831), .Z(n_1501100807
		));
	notech_and3 i_296998228(.A(n_2382), .B(lenpc2[17]), .C(n_60831), .Z(n_1502100808
		));
	notech_and3 i_297098229(.A(n_2382), .B(lenpc2[18]), .C(n_60831), .Z(n_1503100809
		));
	notech_and3 i_297198230(.A(n_2382), .B(lenpc2[19]), .C(n_60837), .Z(n_1504100810
		));
	notech_and3 i_297298231(.A(n_60921), .B(lenpc2[20]), .C(n_60837), .Z(n_1505100811
		));
	notech_and3 i_297398232(.A(n_60921), .B(lenpc2[21]), .C(n_60837), .Z(n_1506100812
		));
	notech_and3 i_297498233(.A(n_60921), .B(lenpc2[22]), .C(n_60831), .Z(n_1507100813
		));
	notech_and3 i_297598234(.A(n_60921), .B(lenpc2[23]), .C(n_60831), .Z(n_1508100814
		));
	notech_and3 i_297698235(.A(n_60921), .B(lenpc2[24]), .C(n_60831), .Z(n_1509100815
		));
	notech_and3 i_297798236(.A(n_60921), .B(lenpc2[25]), .C(n_60831), .Z(n_1510100816
		));
	notech_and3 i_297898237(.A(n_60921), .B(lenpc2[26]), .C(n_60831), .Z(n_1511100817
		));
	notech_and3 i_297998238(.A(n_60921), .B(lenpc2[27]), .C(n_60831), .Z(n_1512100818
		));
	notech_and3 i_298098239(.A(n_60921), .B(lenpc2[28]), .C(n_60836), .Z(n_1513100819
		));
	notech_and3 i_298198240(.A(n_60921), .B(lenpc2[29]), .C(n_60820), .Z(n_1514100820
		));
	notech_and3 i_298298241(.A(n_60921), .B(lenpc2[30]), .C(n_60820), .Z(n_1515100821
		));
	notech_ao3 i_298598242(.A(n_60820), .B(\nbus_12406[1] ), .C(n_60339), .Z
		(n_1516100822));
	notech_ao3 i_298698243(.A(n_60820), .B(\nbus_12406[2] ), .C(n_60337), .Z
		(n_1518100823));
	notech_ao3 i_298798244(.A(n_60820), .B(\nbus_12406[3] ), .C(n_60337), .Z
		(n_1519100824));
	notech_ao3 i_298898245(.A(n_60820), .B(\nbus_12406[4] ), .C(n_60337), .Z
		(n_1520100825));
	notech_ao3 i_12978914(.A(n_60825), .B(\to_acu2_0[20] ), .C(n_60339), .Z(n_1521100826
		));
	notech_ao3 i_21478833(.A(n_60825), .B(\to_acu2_0[29] ), .C(n_60337), .Z(n_1522100827
		));
	notech_ao3 i_21378834(.A(n_60825), .B(\to_acu2_0[30] ), .C(n_60339), .Z(n_1523100828
		));
	notech_ao3 i_5878983(.A(n_60820), .B(\to_acu2_0[45] ), .C(n_60339), .Z(n_1524100829
		));
	notech_ao3 i_12578918(.A(n_60825), .B(in128[16]), .C(n_60339), .Z(n_1525100830
		));
	notech_ao3 i_5078991(.A(n_60825), .B(in128[25]), .C(n_60339), .Z(n_1526100831
		));
	notech_ao3 i_12778916(.A(n_60820), .B(in128[27]), .C(n_60339), .Z(n_1527100832
		));
	notech_ao3 i_22278827(.A(n_60820), .B(in128[41]), .C(n_60339), .Z(n_1528100833
		));
	notech_ao3 i_18078864(.A(n_60820), .B(in128[107]), .C(n_60339), .Z(n_1529100834
		));
	notech_ao3 i_17978865(.A(n_60820), .B(in128[108]), .C(n_60339), .Z(n_1530100835
		));
	notech_ao3 i_17878866(.A(n_60820), .B(in128[109]), .C(n_60339), .Z(n_1531100836
		));
	notech_ao3 i_16378881(.A(n_60820), .B(in128[124]), .C(n_60339), .Z(n_1532100837
		));
	notech_ao3 i_16178883(.A(n_60820), .B(in128[126]), .C(n_60339), .Z(n_1533100838
		));
	notech_and2 i_3299(.A(ififo_rvect3[0]), .B(n_1554100859), .Z(n_1534100839
		));
	notech_and2 i_3304(.A(ififo_rvect3[1]), .B(n_1554100859), .Z(n_1535100840
		));
	notech_and2 i_3305(.A(ififo_rvect3[2]), .B(n_1554100859), .Z(n_1536100841
		));
	notech_and2 i_3306(.A(ififo_rvect3[3]), .B(n_1554100859), .Z(n_1537100842
		));
	notech_and2 i_3307(.A(ififo_rvect3[4]), .B(n_1554100859), .Z(n_1538100843
		));
	notech_and2 i_3308(.A(ififo_rvect3[5]), .B(n_1554100859), .Z(n_1539100844
		));
	notech_and2 i_3309(.A(ififo_rvect3[6]), .B(n_1554100859), .Z(n_1540100845
		));
	notech_and2 i_3310(.A(ififo_rvect3[7]), .B(n_1554100859), .Z(n_1541100846
		));
	notech_ao3 i_3312(.A(n_60820), .B(udeco[0]), .C(n_60337), .Z(n_1542100847
		));
	notech_ao3 i_3317(.A(n_60820), .B(udeco[5]), .C(n_60348), .Z(n_1543100848
		));
	notech_ao3 i_3319(.A(n_60820), .B(udeco[7]), .C(n_60348), .Z(n_1544100849
		));
	notech_ao3 i_3320(.A(n_60820), .B(udeco[8]), .C(n_60348), .Z(n_1545100850
		));
	notech_ao3 i_3353(.A(n_60820), .B(udeco[41]), .C(n_60337), .Z(n_1546100851
		));
	notech_ao3 i_3354(.A(n_60820), .B(udeco[42]), .C(n_60337), .Z(n_1547100852
		));
	notech_ao3 i_3355(.A(n_60825), .B(udeco[43]), .C(n_60348), .Z(n_1548100853
		));
	notech_ao3 i_3356(.A(n_60831), .B(udeco[44]), .C(n_60348), .Z(n_1549100854
		));
	notech_ao3 i_3357(.A(n_60831), .B(udeco[45]), .C(n_60348), .Z(n_1550100855
		));
	notech_and3 i_3686(.A(db67), .B(n_41609), .C(n_1241100548), .Z(n_1551100856
		));
	notech_nao3 i_77378276(.A(n_42556), .B(n_42548), .C(n_2850), .Z(n_1552100857
		));
	notech_nand3 i_77478275(.A(n_1477100783), .B(\to_acu2_0[0] ), .C(\to_acu2_0[1] 
		), .Z(n_1553100858));
	notech_nand2 i_211439(.A(trig_it), .B(n_43377), .Z(n_1554100859));
	notech_ao3 i_627193(.A(n_60831), .B(\nbus_12406[5] ), .C(n_60348), .Z(n_1559100864
		));
	notech_mux2 i_70586(.S(adz), .A(n_41609), .B(n_1714), .Z(n_46118));
	notech_ao4 i_2727750(.A(n_59185), .B(n_42703), .C(n_2603), .D(n_60232), 
		.Z(n_45809));
	notech_xor2 i_110098249(.A(int_excl[3]), .B(n_1755), .Z(n_1563100868));
	notech_nand3 i_327178(.A(n_3029), .B(start), .C(n_1597100902), .Z(n_49863
		));
	notech_xor2 i_110598252(.A(int_excl[1]), .B(int_excl[0]), .Z(n_1566100871
		));
	notech_and4 i_111398256(.A(n_1600100905), .B(adz), .C(n_44684), .D(n_1602100907
		), .Z(n_1570100875));
	notech_xor2 i_110898257(.A(opz[2]), .B(opz[1]), .Z(n_1571100876));
	notech_and3 i_111198258(.A(\to_acu2_0[16] ), .B(twobyte), .C(n_41609), .Z
		(n_1572100877));
	notech_and4 i_111498259(.A(n_41609), .B(n_42551), .C(n_1571100876), .D(n_42550
		), .Z(n_1573100878));
	notech_and4 i_111298260(.A(opz[2]), .B(n_1599100904), .C(n_1744), .D(n_1878
		), .Z(n_1574100879));
	notech_or4 i_323162(.A(n_1574100879), .B(n_1572100877), .C(n_1570100875)
		, .D(n_1573100878), .Z(n_41813));
	notech_and4 i_112598261(.A(n_1600100905), .B(n_1602100907), .C(n_44684),
		 .D(n_44760), .Z(n_1575100880));
	notech_ao3 i_112298262(.A(\to_acu2_0[50] ), .B(n_41609), .C(n_42553), .Z
		(n_1576100881));
	notech_and4 i_112398263(.A(n_41609), .B(n_42550), .C(n_42551), .D(n_44524
		), .Z(n_1577100882));
	notech_and4 i_112498264(.A(n_1599100904), .B(n_1744), .C(n_1878), .D(opz
		[1]), .Z(n_1578100883));
	notech_or4 i_223161(.A(n_1578100883), .B(n_1577100882), .C(n_1576100881)
		, .D(n_1575100880), .Z(n_41807));
	notech_nand3 i_113598265(.A(n_44684), .B(n_1600100905), .C(\to_acu2_0[74] 
		), .Z(n_1579100884));
	notech_ao3 i_113398266(.A(n_44683), .B(n_44682), .C(n_1744), .Z(n_1580100885
		));
	notech_nao3 i_113498267(.A(n_60825), .B(n_1724), .C(n_2994), .Z(n_1581100886
		));
	notech_or4 i_113698268(.A(n_44523), .B(n_1580100885), .C(n_43465), .D(n_1598100903
		), .Z(n_1582100887));
	notech_nand3 i_123160(.A(n_1579100884), .B(n_1582100887), .C(n_1581100886
		), .Z(n_41801));
	notech_xor2 i_123698269(.A(pfx_sz[4]), .B(n_1619100924), .Z(n_1583100888
		));
	notech_xor2 i_123998272(.A(pfx_sz[3]), .B(n_1618100923), .Z(n_1586100891
		));
	notech_xor2 i_124298275(.A(pfx_sz[2]), .B(n_1617100922), .Z(n_1589100894
		));
	notech_ao4 i_226964(.A(n_43465), .B(n_1620100925), .C(n_1621100926), .D(n_44373
		), .Z(n_41736));
	notech_xor2 i_110398283(.A(int_excl[2]), .B(n_1734), .Z(n_1597100902));
	notech_or2 i_110798284(.A(n_42553), .B(\to_acu2_0[50] ), .Z(n_1598100903
		));
	notech_ao3 i_7498285(.A(n_60831), .B(n_42550), .C(n_2994), .Z(n_1599100904
		));
	notech_and4 i_11198286(.A(n_44683), .B(n_44682), .C(n_41609), .D(n_42550
		), .Z(n_1600100905));
	notech_and3 i_19498288(.A(n_2967), .B(n_2964), .C(n_44685), .Z(n_1602100907
		));
	notech_and2 i_299498303(.A(pfx_sz[0]), .B(pfx_sz[1]), .Z(n_1617100922)
		);
	notech_and3 i_2398304(.A(pfx_sz[0]), .B(pfx_sz[2]), .C(pfx_sz[1]), .Z(n_1618100923
		));
	notech_and4 i_123598305(.A(pfx_sz[1]), .B(pfx_sz[0]), .C(pfx_sz[2]), .D(pfx_sz
		[3]), .Z(n_1619100924));
	notech_nand2 i_124798306(.A(pfx_sz[0]), .B(n_44373), .Z(n_1620100925));
	notech_nand2 i_72186(.A(n_5765), .B(n_1098100406), .Z(\nbus_13545[1] )
		);
	notech_nand2 i_73153(.A(n_5765), .B(n_1097100405), .Z(n_46115));
	notech_nand2 i_70836(.A(n_5765), .B(n_17054783), .Z(\nbus_13538[0] ));
	notech_mux2 i_122073(.S(n_62050), .A(lenpc[0]), .B(lenpc1[0]), .Z(lenpc_out
		[0]));
	notech_mux2 i_222074(.S(n_62050), .A(lenpc[1]), .B(lenpc1[1]), .Z(lenpc_out
		[1]));
	notech_mux2 i_322075(.S(n_62050), .A(lenpc[2]), .B(lenpc1[2]), .Z(lenpc_out
		[2]));
	notech_mux2 i_422076(.S(n_62044), .A(lenpc[3]), .B(lenpc1[3]), .Z(lenpc_out
		[3]));
	notech_mux2 i_522077(.S(n_62044), .A(lenpc[4]), .B(lenpc1[4]), .Z(lenpc_out
		[4]));
	notech_mux2 i_622078(.S(n_62044), .A(lenpc[5]), .B(lenpc1[5]), .Z(lenpc_out
		[5]));
	notech_mux2 i_722079(.S(n_62050), .A(lenpc[6]), .B(lenpc1[6]), .Z(lenpc_out
		[6]));
	notech_mux2 i_822080(.S(n_62050), .A(lenpc[7]), .B(lenpc1[7]), .Z(lenpc_out
		[7]));
	notech_mux2 i_922081(.S(n_62050), .A(lenpc[8]), .B(lenpc1[8]), .Z(lenpc_out
		[8]));
	notech_mux2 i_1022082(.S(n_62050), .A(lenpc[9]), .B(lenpc1[9]), .Z(lenpc_out
		[9]));
	notech_mux2 i_1122083(.S(n_62050), .A(lenpc[10]), .B(lenpc1[10]), .Z(lenpc_out
		[10]));
	notech_mux2 i_1222084(.S(n_62050), .A(lenpc[11]), .B(lenpc1[11]), .Z(lenpc_out
		[11]));
	notech_mux2 i_1322085(.S(n_62050), .A(lenpc[12]), .B(lenpc1[12]), .Z(lenpc_out
		[12]));
	notech_mux2 i_1422086(.S(n_62044), .A(lenpc[13]), .B(lenpc1[13]), .Z(lenpc_out
		[13]));
	notech_mux2 i_1522087(.S(n_62044), .A(lenpc[14]), .B(lenpc1[14]), .Z(lenpc_out
		[14]));
	notech_mux2 i_1622088(.S(n_62044), .A(lenpc[15]), .B(lenpc1[15]), .Z(lenpc_out
		[15]));
	notech_mux2 i_1722089(.S(n_62044), .A(lenpc[16]), .B(lenpc1[16]), .Z(lenpc_out
		[16]));
	notech_mux2 i_1822090(.S(n_62044), .A(lenpc[17]), .B(lenpc1[17]), .Z(lenpc_out
		[17]));
	notech_mux2 i_1922091(.S(n_62044), .A(lenpc[18]), .B(lenpc1[18]), .Z(lenpc_out
		[18]));
	notech_mux2 i_2022092(.S(n_62044), .A(lenpc[19]), .B(lenpc1[19]), .Z(lenpc_out
		[19]));
	notech_mux2 i_2122093(.S(n_62044), .A(lenpc[20]), .B(lenpc1[20]), .Z(lenpc_out
		[20]));
	notech_mux2 i_2222094(.S(n_62044), .A(lenpc[21]), .B(lenpc1[21]), .Z(lenpc_out
		[21]));
	notech_mux2 i_2322095(.S(n_62044), .A(lenpc[22]), .B(lenpc1[22]), .Z(lenpc_out
		[22]));
	notech_mux2 i_2422096(.S(n_62044), .A(lenpc[23]), .B(lenpc1[23]), .Z(lenpc_out
		[23]));
	notech_mux2 i_2522097(.S(n_62044), .A(lenpc[24]), .B(lenpc1[24]), .Z(lenpc_out
		[24]));
	notech_mux2 i_2622098(.S(n_62044), .A(lenpc[25]), .B(lenpc1[25]), .Z(lenpc_out
		[25]));
	notech_mux2 i_2722099(.S(n_62050), .A(lenpc[26]), .B(lenpc1[26]), .Z(lenpc_out
		[26]));
	notech_mux2 i_2822100(.S(n_62055), .A(lenpc[27]), .B(lenpc1[27]), .Z(lenpc_out
		[27]));
	notech_mux2 i_2922101(.S(n_62055), .A(lenpc[28]), .B(lenpc1[28]), .Z(lenpc_out
		[28]));
	notech_mux2 i_3022102(.S(n_62055), .A(lenpc[29]), .B(lenpc1[29]), .Z(lenpc_out
		[29]));
	notech_mux2 i_3122103(.S(n_62055), .A(lenpc[30]), .B(lenpc1[30]), .Z(lenpc_out
		[30]));
	notech_mux2 i_3222104(.S(n_62055), .A(lenpc[31]), .B(lenpc1[31]), .Z(lenpc_out
		[31]));
	notech_mux2 i_123106(.S(n_62055), .A(reps0[0]), .B(reps1[0]), .Z(reps[0]
		));
	notech_mux2 i_223107(.S(n_62056), .A(reps0[1]), .B(reps1[1]), .Z(reps[1]
		));
	notech_mux2 i_323108(.S(n_62056), .A(reps0[2]), .B(reps1[2]), .Z(reps[2]
		));
	notech_mux2 i_123109(.S(n_62056), .A(opz0[0]), .B(opz1[0]), .Z(operand_size
		[0]));
	notech_mux2 i_223110(.S(n_62056), .A(opz0[1]), .B(opz1[1]), .Z(operand_size
		[1]));
	notech_mux2 i_323111(.S(n_62056), .A(opz0[2]), .B(opz1[2]), .Z(operand_size
		[2]));
	notech_mux2 i_125127(.S(n_62056), .A(inst_deco[0]), .B(inst_deco1[0]), .Z
		(to_vliw[0]));
	notech_mux2 i_225128(.S(n_62056), .A(inst_deco[1]), .B(inst_deco1[1]), .Z
		(to_vliw[1]));
	notech_mux2 i_325129(.S(n_62055), .A(inst_deco[2]), .B(inst_deco1[2]), .Z
		(to_vliw[2]));
	notech_mux2 i_425130(.S(n_62055), .A(inst_deco[3]), .B(inst_deco1[3]), .Z
		(to_vliw[3]));
	notech_mux2 i_525131(.S(n_62055), .A(inst_deco[4]), .B(inst_deco1[4]), .Z
		(to_vliw[4]));
	notech_mux2 i_625132(.S(n_62050), .A(inst_deco[5]), .B(inst_deco1[5]), .Z
		(to_vliw[5]));
	notech_mux2 i_725133(.S(n_62055), .A(inst_deco[6]), .B(inst_deco1[6]), .Z
		(to_vliw[6]));
	notech_mux2 i_825134(.S(n_62055), .A(inst_deco[7]), .B(inst_deco1[7]), .Z
		(to_vliw[7]));
	notech_mux2 i_925135(.S(n_62055), .A(inst_deco[8]), .B(inst_deco1[8]), .Z
		(to_vliw[8]));
	notech_mux2 i_1025136(.S(n_62055), .A(inst_deco[9]), .B(inst_deco1[9]), 
		.Z(to_vliw[9]));
	notech_mux2 i_1125137(.S(n_62055), .A(inst_deco[10]), .B(inst_deco1[10])
		, .Z(to_vliw[10]));
	notech_mux2 i_1225138(.S(n_62055), .A(inst_deco[11]), .B(inst_deco1[11])
		, .Z(to_vliw[11]));
	notech_mux2 i_1325139(.S(n_62055), .A(inst_deco[12]), .B(inst_deco1[12])
		, .Z(to_vliw[12]));
	notech_mux2 i_1425140(.S(n_62055), .A(inst_deco[13]), .B(inst_deco1[13])
		, .Z(to_vliw[13]));
	notech_mux2 i_1525141(.S(n_62055), .A(inst_deco[14]), .B(inst_deco1[14])
		, .Z(to_vliw[14]));
	notech_mux2 i_1625142(.S(n_62044), .A(inst_deco[15]), .B(inst_deco1[15])
		, .Z(to_vliw[15]));
	notech_mux2 i_1725143(.S(n_62033), .A(inst_deco[16]), .B(inst_deco1[16])
		, .Z(to_vliw[16]));
	notech_mux2 i_1825144(.S(n_62033), .A(inst_deco[17]), .B(inst_deco1[17])
		, .Z(to_vliw[17]));
	notech_mux2 i_1925145(.S(n_62033), .A(inst_deco[18]), .B(inst_deco1[18])
		, .Z(to_vliw[18]));
	notech_mux2 i_2025146(.S(n_62033), .A(inst_deco[19]), .B(inst_deco1[19])
		, .Z(to_vliw[19]));
	notech_mux2 i_2125147(.S(n_62033), .A(inst_deco[20]), .B(inst_deco1[20])
		, .Z(to_vliw[20]));
	notech_mux2 i_2225148(.S(n_62033), .A(inst_deco[21]), .B(inst_deco1[21])
		, .Z(to_vliw[21]));
	notech_mux2 i_2325149(.S(n_62033), .A(inst_deco[22]), .B(inst_deco1[22])
		, .Z(to_vliw[22]));
	notech_mux2 i_2425150(.S(n_62038), .A(inst_deco[23]), .B(inst_deco1[23])
		, .Z(to_vliw[23]));
	notech_mux2 i_2525151(.S(n_62038), .A(inst_deco[24]), .B(inst_deco1[24])
		, .Z(to_vliw[24]));
	notech_mux2 i_2625152(.S(n_62038), .A(inst_deco[25]), .B(inst_deco1[25])
		, .Z(to_vliw[25]));
	notech_mux2 i_2725153(.S(n_62033), .A(inst_deco[26]), .B(inst_deco1[26])
		, .Z(to_vliw[26]));
	notech_mux2 i_2825154(.S(n_62033), .A(inst_deco[27]), .B(inst_deco1[27])
		, .Z(to_vliw[27]));
	notech_mux2 i_2925155(.S(n_62038), .A(inst_deco[28]), .B(inst_deco1[28])
		, .Z(to_vliw[28]));
	notech_mux2 i_3025156(.S(n_62032), .A(inst_deco[29]), .B(inst_deco1[29])
		, .Z(to_vliw[29]));
	notech_mux2 i_3125157(.S(n_62033), .A(inst_deco[30]), .B(inst_deco1[30])
		, .Z(to_vliw[30]));
	notech_mux2 i_3225158(.S(n_62033), .A(inst_deco[31]), .B(inst_deco1[31])
		, .Z(to_vliw[31]));
	notech_mux2 i_3325159(.S(n_62032), .A(inst_deco[32]), .B(inst_deco1[32])
		, .Z(to_vliw[32]));
	notech_mux2 i_3425160(.S(n_62032), .A(inst_deco[33]), .B(inst_deco1[33])
		, .Z(to_vliw[33]));
	notech_mux2 i_3525161(.S(n_62032), .A(inst_deco[34]), .B(inst_deco1[34])
		, .Z(to_vliw[34]));
	notech_mux2 i_3625162(.S(n_62033), .A(inst_deco[35]), .B(inst_deco1[35])
		, .Z(to_vliw[35]));
	notech_mux2 i_3725163(.S(n_62033), .A(inst_deco[36]), .B(inst_deco1[36])
		, .Z(to_vliw[36]));
	notech_mux2 i_3825164(.S(n_62033), .A(inst_deco[37]), .B(inst_deco1[37])
		, .Z(to_vliw[37]));
	notech_mux2 i_3925165(.S(n_62033), .A(inst_deco[38]), .B(inst_deco1[38])
		, .Z(to_vliw[38]));
	notech_mux2 i_4025166(.S(n_62033), .A(inst_deco[39]), .B(inst_deco1[39])
		, .Z(to_vliw[39]));
	notech_mux2 i_4125167(.S(n_62033), .A(inst_deco[40]), .B(inst_deco1[40])
		, .Z(to_vliw[40]));
	notech_mux2 i_4225168(.S(n_62033), .A(inst_deco[41]), .B(inst_deco1[41])
		, .Z(to_vliw[41]));
	notech_mux2 i_4325169(.S(n_62038), .A(inst_deco[42]), .B(inst_deco1[42])
		, .Z(to_vliw[42]));
	notech_mux2 i_4425170(.S(n_62043), .A(inst_deco[43]), .B(inst_deco1[43])
		, .Z(to_vliw[43]));
	notech_mux2 i_4525171(.S(n_62043), .A(inst_deco[44]), .B(inst_deco1[44])
		, .Z(to_vliw[44]));
	notech_mux2 i_4625172(.S(n_62043), .A(inst_deco[45]), .B(inst_deco1[45])
		, .Z(to_vliw[45]));
	notech_mux2 i_4725173(.S(n_62043), .A(inst_deco[46]), .B(inst_deco1[46])
		, .Z(to_vliw[46]));
	notech_mux2 i_4825174(.S(n_62043), .A(inst_deco[47]), .B(inst_deco1[47])
		, .Z(to_vliw[47]));
	notech_mux2 i_4925175(.S(n_62043), .A(inst_deco[48]), .B(inst_deco1[48])
		, .Z(to_vliw[48]));
	notech_mux2 i_5025176(.S(n_62043), .A(inst_deco[49]), .B(inst_deco1[49])
		, .Z(to_vliw[49]));
	notech_mux2 i_5125177(.S(n_62043), .A(inst_deco[50]), .B(inst_deco1[50])
		, .Z(to_vliw[50]));
	notech_mux2 i_5225178(.S(n_62043), .A(inst_deco[51]), .B(inst_deco1[51])
		, .Z(to_vliw[51]));
	notech_mux2 i_5325179(.S(n_62044), .A(inst_deco[52]), .B(inst_deco1[52])
		, .Z(to_vliw[52]));
	notech_mux2 i_5425180(.S(n_62043), .A(inst_deco[53]), .B(inst_deco1[53])
		, .Z(to_vliw[53]));
	notech_mux2 i_5525181(.S(n_62043), .A(inst_deco[54]), .B(inst_deco1[54])
		, .Z(to_vliw[54]));
	notech_mux2 i_5625182(.S(n_62043), .A(inst_deco[55]), .B(inst_deco1[55])
		, .Z(to_vliw[55]));
	notech_mux2 i_5725183(.S(n_62038), .A(inst_deco[56]), .B(inst_deco1[56])
		, .Z(to_vliw[56]));
	notech_mux2 i_5825184(.S(n_62038), .A(inst_deco[57]), .B(inst_deco1[57])
		, .Z(to_vliw[57]));
	notech_mux2 i_5925185(.S(n_62038), .A(inst_deco[58]), .B(inst_deco1[58])
		, .Z(to_vliw[58]));
	notech_mux2 i_6025186(.S(n_62038), .A(inst_deco[59]), .B(inst_deco1[59])
		, .Z(to_vliw[59]));
	notech_mux2 i_6125187(.S(n_62038), .A(inst_deco[60]), .B(inst_deco1[60])
		, .Z(to_vliw[60]));
	notech_mux2 i_6225188(.S(n_62038), .A(inst_deco[61]), .B(inst_deco1[61])
		, .Z(to_vliw[61]));
	notech_mux2 i_6325189(.S(n_62038), .A(inst_deco[62]), .B(inst_deco1[62])
		, .Z(to_vliw[62]));
	notech_mux2 i_6425190(.S(n_62043), .A(inst_deco[63]), .B(inst_deco1[63])
		, .Z(to_vliw[63]));
	notech_mux2 i_6525191(.S(n_62043), .A(inst_deco[64]), .B(inst_deco1[64])
		, .Z(to_vliw[64]));
	notech_mux2 i_6625192(.S(n_62043), .A(inst_deco[65]), .B(inst_deco1[65])
		, .Z(to_vliw[65]));
	notech_mux2 i_6725193(.S(n_62043), .A(inst_deco[66]), .B(inst_deco1[66])
		, .Z(to_vliw[66]));
	notech_mux2 i_6825194(.S(n_62043), .A(inst_deco[67]), .B(inst_deco1[67])
		, .Z(to_vliw[67]));
	notech_mux2 i_6925195(.S(n_62043), .A(inst_deco[68]), .B(inst_deco1[68])
		, .Z(to_vliw[68]));
	notech_mux2 i_7025196(.S(n_62072), .A(inst_deco[69]), .B(inst_deco1[69])
		, .Z(to_vliw[69]));
	notech_mux2 i_7125197(.S(n_62077), .A(inst_deco[70]), .B(inst_deco1[70])
		, .Z(to_vliw[70]));
	notech_mux2 i_7225198(.S(n_62077), .A(inst_deco[71]), .B(inst_deco1[71])
		, .Z(to_vliw[71]));
	notech_mux2 i_7325199(.S(n_62072), .A(inst_deco[72]), .B(inst_deco1[72])
		, .Z(to_vliw[72]));
	notech_mux2 i_7425200(.S(n_62072), .A(inst_deco[73]), .B(inst_deco1[73])
		, .Z(to_vliw[73]));
	notech_mux2 i_7525201(.S(n_62072), .A(inst_deco[74]), .B(inst_deco1[74])
		, .Z(to_vliw[74]));
	notech_mux2 i_7625202(.S(n_62077), .A(inst_deco[75]), .B(inst_deco1[75])
		, .Z(to_vliw[75]));
	notech_mux2 i_7725203(.S(n_62077), .A(inst_deco[76]), .B(inst_deco1[76])
		, .Z(to_vliw[76]));
	notech_mux2 i_7825204(.S(n_62077), .A(inst_deco[77]), .B(inst_deco1[77])
		, .Z(to_vliw[77]));
	notech_mux2 i_7925205(.S(n_62077), .A(inst_deco[78]), .B(inst_deco1[78])
		, .Z(to_vliw[78]));
	notech_mux2 i_8025206(.S(n_62077), .A(inst_deco[79]), .B(inst_deco1[79])
		, .Z(to_vliw[79]));
	notech_mux2 i_8125207(.S(n_62077), .A(inst_deco[80]), .B(inst_deco1[80])
		, .Z(to_vliw[80]));
	notech_mux2 i_8225208(.S(n_62077), .A(inst_deco[81]), .B(inst_deco1[81])
		, .Z(to_vliw[81]));
	notech_mux2 i_8325209(.S(n_62067), .A(inst_deco[82]), .B(inst_deco1[82])
		, .Z(to_vliw[82]));
	notech_mux2 i_8425210(.S(n_62067), .A(inst_deco[83]), .B(inst_deco1[83])
		, .Z(to_vliw[83]));
	notech_mux2 i_8525211(.S(n_62072), .A(inst_deco[84]), .B(inst_deco1[84])
		, .Z(to_vliw[84]));
	notech_mux2 i_8625212(.S(n_62067), .A(inst_deco[85]), .B(inst_deco1[85])
		, .Z(to_vliw[85]));
	notech_mux2 i_8725213(.S(n_62067), .A(inst_deco[86]), .B(inst_deco1[86])
		, .Z(to_vliw[86]));
	notech_mux2 i_8825214(.S(n_62067), .A(inst_deco[87]), .B(inst_deco1[87])
		, .Z(to_vliw[87]));
	notech_mux2 i_8925215(.S(n_62072), .A(inst_deco[88]), .B(inst_deco1[88])
		, .Z(to_vliw[88]));
	notech_mux2 i_9025216(.S(n_62072), .A(inst_deco[89]), .B(inst_deco1[89])
		, .Z(to_vliw[89]));
	notech_mux2 i_9125217(.S(n_62072), .A(inst_deco[90]), .B(inst_deco1[90])
		, .Z(to_vliw[90]));
	notech_mux2 i_9225218(.S(n_62072), .A(inst_deco[91]), .B(inst_deco1[91])
		, .Z(to_vliw[91]));
	notech_mux2 i_9325219(.S(n_62072), .A(inst_deco[92]), .B(inst_deco1[92])
		, .Z(to_vliw[92]));
	notech_mux2 i_9425220(.S(n_62072), .A(inst_deco[93]), .B(inst_deco1[93])
		, .Z(to_vliw[93]));
	notech_mux2 i_9525221(.S(n_62072), .A(inst_deco[94]), .B(inst_deco1[94])
		, .Z(to_vliw[94]));
	notech_mux2 i_9625222(.S(n_62077), .A(inst_deco[95]), .B(inst_deco1[95])
		, .Z(to_vliw[95]));
	notech_mux2 i_9725223(.S(n_62078), .A(inst_deco[96]), .B(inst_deco1[96])
		, .Z(to_vliw[96]));
	notech_mux2 i_9825224(.S(n_62078), .A(inst_deco[97]), .B(inst_deco1[97])
		, .Z(to_vliw[97]));
	notech_mux2 i_9925225(.S(n_62078), .A(inst_deco[98]), .B(inst_deco1[98])
		, .Z(to_vliw[98]));
	notech_mux2 i_10025226(.S(n_62078), .A(inst_deco[99]), .B(inst_deco1[99]
		), .Z(to_vliw[99]));
	notech_mux2 i_10125227(.S(n_62078), .A(inst_deco[100]), .B(inst_deco1[
		100]), .Z(to_vliw[100]));
	notech_mux2 i_10225228(.S(n_62078), .A(inst_deco[101]), .B(inst_deco1[
		101]), .Z(to_vliw[101]));
	notech_mux2 i_10325229(.S(n_62078), .A(inst_deco[102]), .B(inst_deco1[
		102]), .Z(to_vliw[102]));
	notech_mux2 i_10425230(.S(n_62078), .A(inst_deco[103]), .B(inst_deco1[
		103]), .Z(to_vliw[103]));
	notech_mux2 i_10525231(.S(n_62078), .A(inst_deco[104]), .B(inst_deco1[
		104]), .Z(to_vliw[104]));
	notech_mux2 i_10625232(.S(n_62078), .A(inst_deco[105]), .B(inst_deco1[
		105]), .Z(to_vliw[105]));
	notech_mux2 i_10725233(.S(n_62078), .A(inst_deco[106]), .B(inst_deco1[
		106]), .Z(to_vliw[106]));
	notech_mux2 i_10825234(.S(n_62078), .A(inst_deco[107]), .B(inst_deco1[
		107]), .Z(to_vliw[107]));
	notech_mux2 i_10925235(.S(n_62078), .A(inst_deco[108]), .B(inst_deco1[
		108]), .Z(to_vliw[108]));
	notech_mux2 i_11025236(.S(n_62077), .A(inst_deco[109]), .B(inst_deco1[
		109]), .Z(to_vliw[109]));
	notech_mux2 i_11125237(.S(n_62077), .A(inst_deco[110]), .B(inst_deco1[
		110]), .Z(to_vliw[110]));
	notech_mux2 i_11225238(.S(n_62077), .A(inst_deco[111]), .B(inst_deco1[
		111]), .Z(to_vliw[111]));
	notech_mux2 i_11325239(.S(n_62077), .A(inst_deco[112]), .B(inst_deco1[
		112]), .Z(to_vliw[112]));
	notech_mux2 i_11425240(.S(n_62077), .A(inst_deco[113]), .B(inst_deco1[
		113]), .Z(to_vliw[113]));
	notech_mux2 i_11525241(.S(n_62077), .A(inst_deco[114]), .B(inst_deco1[
		114]), .Z(to_vliw[114]));
	notech_mux2 i_11625242(.S(n_62077), .A(inst_deco[115]), .B(inst_deco1[
		115]), .Z(to_vliw[115]));
	notech_mux2 i_11725243(.S(n_62078), .A(inst_deco[116]), .B(inst_deco1[
		116]), .Z(to_vliw[116]));
	notech_mux2 i_11825244(.S(n_62078), .A(inst_deco[117]), .B(inst_deco1[
		117]), .Z(to_vliw[117]));
	notech_mux2 i_11925245(.S(n_62078), .A(inst_deco[118]), .B(inst_deco1[
		118]), .Z(to_vliw[118]));
	notech_mux2 i_12025246(.S(n_62077), .A(inst_deco[119]), .B(inst_deco1[
		119]), .Z(to_vliw[119]));
	notech_mux2 i_12125247(.S(n_62078), .A(inst_deco[120]), .B(inst_deco1[
		120]), .Z(to_vliw[120]));
	notech_mux2 i_12225248(.S(n_62078), .A(inst_deco[121]), .B(inst_deco1[
		121]), .Z(to_vliw[121]));
	notech_mux2 i_12325249(.S(n_62067), .A(inst_deco[122]), .B(inst_deco1[
		122]), .Z(to_vliw[122]));
	notech_mux2 i_12425250(.S(n_62061), .A(inst_deco[123]), .B(inst_deco1[
		123]), .Z(to_vliw[123]));
	notech_mux2 i_12525251(.S(n_62061), .A(inst_deco[124]), .B(inst_deco1[
		124]), .Z(to_vliw[124]));
	notech_mux2 i_12625252(.S(n_62061), .A(inst_deco[125]), .B(inst_deco1[
		125]), .Z(to_vliw[125]));
	notech_mux2 i_12725253(.S(n_62061), .A(inst_deco[126]), .B(inst_deco1[
		126]), .Z(to_vliw[126]));
	notech_mux2 i_12825254(.S(n_62061), .A(inst_deco[127]), .B(inst_deco1[
		127]), .Z(to_vliw[127]));
	notech_mux2 i_125895(.S(n_62061), .A(to_acu0[0]), .B(to_acu1[0]), .Z(to_acu
		[0]));
	notech_mux2 i_225896(.S(n_62061), .A(to_acu0[1]), .B(to_acu1[1]), .Z(to_acu
		[1]));
	notech_mux2 i_325897(.S(n_62066), .A(to_acu0[2]), .B(to_acu1[2]), .Z(to_acu
		[2]));
	notech_mux2 i_425898(.S(n_62066), .A(to_acu0[3]), .B(to_acu1[3]), .Z(to_acu
		[3]));
	notech_mux2 i_525899(.S(n_62066), .A(to_acu0[4]), .B(to_acu1[4]), .Z(to_acu
		[4]));
	notech_mux2 i_625900(.S(n_62061), .A(to_acu0[5]), .B(to_acu1[5]), .Z(to_acu
		[5]));
	notech_mux2 i_725901(.S(n_62061), .A(to_acu0[6]), .B(to_acu1[6]), .Z(to_acu
		[6]));
	notech_mux2 i_825902(.S(n_62061), .A(to_acu0[7]), .B(to_acu1[7]), .Z(to_acu
		[7]));
	notech_mux2 i_925903(.S(n_62056), .A(to_acu0[8]), .B(to_acu1[8]), .Z(to_acu
		[8]));
	notech_mux2 i_1025904(.S(n_62056), .A(to_acu0[9]), .B(to_acu1[9]), .Z(to_acu
		[9]));
	notech_mux2 i_1125905(.S(n_62056), .A(to_acu0[10]), .B(to_acu1[10]), .Z(to_acu
		[10]));
	notech_mux2 i_1225906(.S(n_62056), .A(to_acu0[11]), .B(to_acu1[11]), .Z(to_acu
		[11]));
	notech_mux2 i_1325907(.S(n_62056), .A(to_acu0[12]), .B(to_acu1[12]), .Z(to_acu
		[12]));
	notech_mux2 i_1425908(.S(n_62056), .A(to_acu0[13]), .B(to_acu1[13]), .Z(to_acu
		[13]));
	notech_mux2 i_1525909(.S(n_62056), .A(to_acu0[14]), .B(to_acu1[14]), .Z(to_acu
		[14]));
	notech_mux2 i_1625910(.S(n_62056), .A(to_acu0[15]), .B(to_acu1[15]), .Z(to_acu
		[15]));
	notech_mux2 i_1725911(.S(n_62061), .A(to_acu0[16]), .B(to_acu1[16]), .Z(to_acu
		[16]));
	notech_mux2 i_1825912(.S(n_62061), .A(to_acu0[17]), .B(to_acu1[17]), .Z(to_acu
		[17]));
	notech_mux2 i_1925913(.S(n_62056), .A(to_acu0[18]), .B(to_acu1[18]), .Z(to_acu
		[18]));
	notech_mux2 i_2025914(.S(n_62056), .A(to_acu0[19]), .B(to_acu1[19]), .Z(to_acu
		[19]));
	notech_mux2 i_2125915(.S(n_62056), .A(to_acu0[20]), .B(to_acu1[20]), .Z(to_acu
		[20]));
	notech_mux2 i_2225916(.S(n_62066), .A(to_acu0[21]), .B(to_acu1[21]), .Z(to_acu
		[21]));
	notech_mux2 i_2325917(.S(n_62067), .A(to_acu0[22]), .B(to_acu1[22]), .Z(to_acu
		[22]));
	notech_mux2 i_2425918(.S(n_62067), .A(to_acu0[23]), .B(to_acu1[23]), .Z(to_acu
		[23]));
	notech_mux2 i_2525919(.S(n_62067), .A(to_acu0[24]), .B(to_acu1[24]), .Z(to_acu
		[24]));
	notech_mux2 i_2625920(.S(n_62066), .A(to_acu0[25]), .B(to_acu1[25]), .Z(to_acu
		[25]));
	notech_mux2 i_2725921(.S(n_62067), .A(to_acu0[26]), .B(to_acu1[26]), .Z(to_acu
		[26]));
	notech_mux2 i_2825922(.S(n_62067), .A(to_acu0[27]), .B(to_acu1[27]), .Z(to_acu
		[27]));
	notech_mux2 i_2925923(.S(n_62067), .A(to_acu0[28]), .B(to_acu1[28]), .Z(to_acu
		[28]));
	notech_mux2 i_3025924(.S(n_62067), .A(to_acu0[29]), .B(to_acu1[29]), .Z(to_acu
		[29]));
	notech_mux2 i_3125925(.S(n_62067), .A(to_acu0[30]), .B(to_acu1[30]), .Z(to_acu
		[30]));
	notech_mux2 i_3225926(.S(n_62067), .A(to_acu0[31]), .B(to_acu1[31]), .Z(to_acu
		[31]));
	notech_mux2 i_3325927(.S(n_62067), .A(to_acu0[32]), .B(to_acu1[32]), .Z(to_acu
		[32]));
	notech_mux2 i_3425928(.S(n_62067), .A(to_acu0[33]), .B(to_acu1[33]), .Z(to_acu
		[33]));
	notech_mux2 i_3525929(.S(n_62067), .A(to_acu0[34]), .B(to_acu1[34]), .Z(to_acu
		[34]));
	notech_mux2 i_3625930(.S(n_62066), .A(to_acu0[35]), .B(to_acu1[35]), .Z(to_acu
		[35]));
	notech_mux2 i_3725931(.S(n_62066), .A(to_acu0[36]), .B(to_acu1[36]), .Z(to_acu
		[36]));
	notech_mux2 i_3825932(.S(n_62066), .A(to_acu0[37]), .B(to_acu1[37]), .Z(to_acu
		[37]));
	notech_mux2 i_3925933(.S(n_62066), .A(to_acu0[38]), .B(to_acu1[38]), .Z(to_acu
		[38]));
	notech_mux2 i_4025934(.S(n_62066), .A(to_acu0[39]), .B(to_acu1[39]), .Z(to_acu
		[39]));
	notech_mux2 i_4125935(.S(n_62066), .A(to_acu0[40]), .B(to_acu1[40]), .Z(to_acu
		[40]));
	notech_mux2 i_4225936(.S(n_62066), .A(to_acu0[41]), .B(to_acu1[41]), .Z(to_acu
		[41]));
	notech_mux2 i_4325937(.S(n_62066), .A(to_acu0[42]), .B(to_acu1[42]), .Z(to_acu
		[42]));
	notech_mux2 i_4425938(.S(n_62066), .A(to_acu0[43]), .B(to_acu1[43]), .Z(to_acu
		[43]));
	notech_mux2 i_4525939(.S(n_62066), .A(to_acu0[44]), .B(to_acu1[44]), .Z(to_acu
		[44]));
	notech_mux2 i_4625940(.S(n_62066), .A(to_acu0[45]), .B(to_acu1[45]), .Z(to_acu
		[45]));
	notech_mux2 i_4725941(.S(n_62066), .A(to_acu0[46]), .B(to_acu1[46]), .Z(to_acu
		[46]));
	notech_mux2 i_4825942(.S(n_62066), .A(to_acu0[47]), .B(to_acu1[47]), .Z(to_acu
		[47]));
	notech_mux2 i_4925943(.S(n_62032), .A(to_acu0[48]), .B(to_acu1[48]), .Z(to_acu
		[48]));
	notech_mux2 i_5025944(.S(n_61998), .A(to_acu0[49]), .B(to_acu1[49]), .Z(to_acu
		[49]));
	notech_mux2 i_5125945(.S(n_61998), .A(to_acu0[50]), .B(to_acu1[50]), .Z(to_acu
		[50]));
	notech_mux2 i_5225946(.S(n_61998), .A(to_acu0[51]), .B(to_acu1[51]), .Z(to_acu
		[51]));
	notech_mux2 i_5325947(.S(n_61998), .A(to_acu0[52]), .B(to_acu1[52]), .Z(to_acu
		[52]));
	notech_mux2 i_5425948(.S(n_61998), .A(to_acu0[53]), .B(to_acu1[53]), .Z(to_acu
		[53]));
	notech_mux2 i_5525949(.S(n_61998), .A(to_acu0[54]), .B(to_acu1[54]), .Z(to_acu
		[54]));
	notech_mux2 i_5625950(.S(n_61998), .A(to_acu0[55]), .B(to_acu1[55]), .Z(to_acu
		[55]));
	notech_mux2 i_5725951(.S(n_61999), .A(to_acu0[56]), .B(to_acu1[56]), .Z(to_acu
		[56]));
	notech_mux2 i_5825952(.S(n_61999), .A(to_acu0[57]), .B(to_acu1[57]), .Z(to_acu
		[57]));
	notech_mux2 i_5925953(.S(n_61999), .A(to_acu0[58]), .B(to_acu1[58]), .Z(to_acu
		[58]));
	notech_mux2 i_6025954(.S(n_61998), .A(to_acu0[59]), .B(to_acu1[59]), .Z(to_acu
		[59]));
	notech_mux2 i_6125955(.S(n_61999), .A(to_acu0[60]), .B(to_acu1[60]), .Z(to_acu
		[60]));
	notech_mux2 i_6225956(.S(n_61999), .A(to_acu0[61]), .B(to_acu1[61]), .Z(to_acu
		[61]));
	notech_mux2 i_6325957(.S(n_61998), .A(to_acu0[62]), .B(to_acu1[62]), .Z(to_acu
		[62]));
	notech_mux2 i_6425958(.S(n_61998), .A(to_acu0[63]), .B(to_acu1[63]), .Z(to_acu
		[63]));
	notech_mux2 i_6525959(.S(n_61998), .A(to_acu0[64]), .B(to_acu1[64]), .Z(to_acu
		[64]));
	notech_mux2 i_6625960(.S(n_61993), .A(to_acu0[65]), .B(to_acu1[65]), .Z(to_acu
		[65]));
	notech_mux2 i_6725961(.S(n_61993), .A(to_acu0[66]), .B(to_acu1[66]), .Z(to_acu
		[66]));
	notech_mux2 i_6825962(.S(n_61993), .A(to_acu0[67]), .B(to_acu1[67]), .Z(to_acu
		[67]));
	notech_mux2 i_6925963(.S(n_61998), .A(to_acu0[68]), .B(to_acu1[68]), .Z(to_acu
		[68]));
	notech_mux2 i_7025964(.S(n_61998), .A(to_acu0[69]), .B(to_acu1[69]), .Z(to_acu
		[69]));
	notech_mux2 i_7125965(.S(n_61998), .A(to_acu0[70]), .B(to_acu1[70]), .Z(to_acu
		[70]));
	notech_mux2 i_7225966(.S(n_61998), .A(to_acu0[71]), .B(to_acu1[71]), .Z(to_acu
		[71]));
	notech_mux2 i_7325967(.S(n_61998), .A(to_acu0[72]), .B(to_acu1[72]), .Z(to_acu
		[72]));
	notech_mux2 i_7425968(.S(n_61998), .A(to_acu0[73]), .B(to_acu1[73]), .Z(to_acu
		[73]));
	notech_mux2 i_7525969(.S(n_61998), .A(to_acu0[74]), .B(to_acu1[74]), .Z(to_acu
		[74]));
	notech_mux2 i_7625970(.S(n_61999), .A(to_acu0[75]), .B(to_acu1[75]), .Z(to_acu
		[75]));
	notech_mux2 i_7725971(.S(n_62004), .A(to_acu0[76]), .B(to_acu1[76]), .Z(to_acu
		[76]));
	notech_mux2 i_7825972(.S(n_62004), .A(to_acu0[77]), .B(to_acu1[77]), .Z(to_acu
		[77]));
	notech_mux2 i_7925973(.S(n_62004), .A(to_acu0[78]), .B(to_acu1[78]), .Z(to_acu
		[78]));
	notech_mux2 i_8025974(.S(n_62004), .A(to_acu0[79]), .B(to_acu1[79]), .Z(to_acu
		[79]));
	notech_mux2 i_8125975(.S(n_62004), .A(to_acu0[80]), .B(to_acu1[80]), .Z(to_acu
		[80]));
	notech_mux2 i_8225976(.S(n_62004), .A(to_acu0[81]), .B(to_acu1[81]), .Z(to_acu
		[81]));
	notech_mux2 i_8325977(.S(n_62004), .A(to_acu0[82]), .B(to_acu1[82]), .Z(to_acu
		[82]));
	notech_mux2 i_8425978(.S(n_62004), .A(to_acu0[83]), .B(to_acu1[83]), .Z(to_acu
		[83]));
	notech_mux2 i_8525979(.S(n_62009), .A(to_acu0[84]), .B(to_acu1[84]), .Z(to_acu
		[84]));
	notech_mux2 i_8625980(.S(n_62009), .A(to_acu0[85]), .B(to_acu1[85]), .Z(to_acu
		[85]));
	notech_mux2 i_8725981(.S(n_62004), .A(to_acu0[86]), .B(to_acu1[86]), .Z(to_acu
		[86]));
	notech_mux2 i_8825982(.S(n_62004), .A(to_acu0[87]), .B(to_acu1[87]), .Z(to_acu
		[87]));
	notech_mux2 i_8925983(.S(n_62004), .A(to_acu0[88]), .B(to_acu1[88]), .Z(to_acu
		[88]));
	notech_mux2 i_9025984(.S(n_61999), .A(to_acu0[89]), .B(to_acu1[89]), .Z(to_acu
		[89]));
	notech_mux2 i_9125985(.S(n_61999), .A(to_acu0[90]), .B(to_acu1[90]), .Z(to_acu
		[90]));
	notech_mux2 i_9225986(.S(n_61999), .A(to_acu0[91]), .B(to_acu1[91]), .Z(to_acu
		[91]));
	notech_mux2 i_9325987(.S(n_61999), .A(to_acu0[92]), .B(to_acu1[92]), .Z(to_acu
		[92]));
	notech_mux2 i_9425988(.S(n_61999), .A(to_acu0[93]), .B(to_acu1[93]), .Z(to_acu
		[93]));
	notech_mux2 i_9525989(.S(n_61999), .A(to_acu0[94]), .B(to_acu1[94]), .Z(to_acu
		[94]));
	notech_mux2 i_9625990(.S(n_61999), .A(to_acu0[95]), .B(to_acu1[95]), .Z(to_acu
		[95]));
	notech_mux2 i_9725991(.S(n_61999), .A(to_acu0[96]), .B(to_acu1[96]), .Z(to_acu
		[96]));
	notech_mux2 i_9825992(.S(n_61999), .A(to_acu0[97]), .B(to_acu1[97]), .Z(to_acu
		[97]));
	notech_mux2 i_9925993(.S(n_62004), .A(to_acu0[98]), .B(to_acu1[98]), .Z(to_acu
		[98]));
	notech_mux2 i_10025994(.S(n_61999), .A(to_acu0[99]), .B(to_acu1[99]), .Z
		(to_acu[99]));
	notech_mux2 i_10125995(.S(n_61999), .A(to_acu0[100]), .B(to_acu1[100]), 
		.Z(to_acu[100]));
	notech_mux2 i_10225996(.S(n_61999), .A(to_acu0[101]), .B(to_acu1[101]), 
		.Z(to_acu[101]));
	notech_mux2 i_10325997(.S(n_61993), .A(to_acu0[102]), .B(to_acu1[102]), 
		.Z(to_acu[102]));
	notech_mux2 i_10425998(.S(n_61987), .A(to_acu0[103]), .B(to_acu1[103]), 
		.Z(to_acu[103]));
	notech_mux2 i_10525999(.S(n_61987), .A(to_acu0[104]), .B(to_acu1[104]), 
		.Z(to_acu[104]));
	notech_mux2 i_10626000(.S(n_61987), .A(to_acu0[105]), .B(to_acu1[105]), 
		.Z(to_acu[105]));
	notech_mux2 i_10726001(.S(n_61987), .A(to_acu0[106]), .B(to_acu1[106]), 
		.Z(to_acu[106]));
	notech_mux2 i_10826002(.S(n_61987), .A(to_acu0[107]), .B(to_acu1[107]), 
		.Z(to_acu[107]));
	notech_mux2 i_10926003(.S(n_61987), .A(to_acu0[108]), .B(to_acu1[108]), 
		.Z(to_acu[108]));
	notech_mux2 i_11026004(.S(n_61987), .A(to_acu0[109]), .B(to_acu1[109]), 
		.Z(to_acu[109]));
	notech_mux2 i_11126005(.S(n_61987), .A(to_acu0[110]), .B(to_acu1[110]), 
		.Z(to_acu[110]));
	notech_mux2 i_11226006(.S(n_61987), .A(to_acu0[111]), .B(to_acu1[111]), 
		.Z(to_acu[111]));
	notech_mux2 i_11326007(.S(n_61987), .A(to_acu0[112]), .B(to_acu1[112]), 
		.Z(to_acu[112]));
	notech_mux2 i_11426008(.S(n_61987), .A(to_acu0[113]), .B(to_acu1[113]), 
		.Z(to_acu[113]));
	notech_mux2 i_11526009(.S(n_61987), .A(to_acu0[114]), .B(to_acu1[114]), 
		.Z(to_acu[114]));
	notech_mux2 i_11626010(.S(n_61987), .A(to_acu0[115]), .B(to_acu1[115]), 
		.Z(to_acu[115]));
	notech_mux2 i_11726011(.S(n_61982), .A(to_acu0[116]), .B(to_acu1[116]), 
		.Z(to_acu[116]));
	notech_mux2 i_11826012(.S(n_61982), .A(to_acu0[117]), .B(to_acu1[117]), 
		.Z(to_acu[117]));
	notech_mux2 i_11926013(.S(n_61982), .A(to_acu0[118]), .B(to_acu1[118]), 
		.Z(to_acu[118]));
	notech_mux2 i_12026014(.S(n_61982), .A(to_acu0[119]), .B(to_acu1[119]), 
		.Z(to_acu[119]));
	notech_mux2 i_12126015(.S(n_61982), .A(to_acu0[120]), .B(to_acu1[120]), 
		.Z(to_acu[120]));
	notech_mux2 i_12226016(.S(n_61982), .A(to_acu0[121]), .B(to_acu1[121]), 
		.Z(to_acu[121]));
	notech_mux2 i_12326017(.S(n_61982), .A(to_acu0[122]), .B(to_acu1[122]), 
		.Z(to_acu[122]));
	notech_mux2 i_12426018(.S(n_61987), .A(to_acu0[123]), .B(to_acu1[123]), 
		.Z(to_acu[123]));
	notech_mux2 i_12526019(.S(n_61987), .A(to_acu0[124]), .B(to_acu1[124]), 
		.Z(to_acu[124]));
	notech_mux2 i_12626020(.S(n_61987), .A(to_acu0[125]), .B(to_acu1[125]), 
		.Z(to_acu[125]));
	notech_mux2 i_12726021(.S(n_61982), .A(to_acu0[126]), .B(to_acu1[126]), 
		.Z(to_acu[126]));
	notech_mux2 i_12826022(.S(n_61982), .A(to_acu0[127]), .B(to_acu1[127]), 
		.Z(to_acu[127]));
	notech_mux2 i_12926023(.S(n_61982), .A(to_acu0[128]), .B(to_acu1[128]), 
		.Z(to_acu[128]));
	notech_mux2 i_13026024(.S(n_61987), .A(to_acu0[129]), .B(to_acu1[129]), 
		.Z(to_acu[129]));
	notech_mux2 i_13126025(.S(n_61988), .A(to_acu0[130]), .B(to_acu1[130]), 
		.Z(to_acu[130]));
	notech_mux2 i_13226026(.S(n_61988), .A(to_acu0[131]), .B(to_acu1[131]), 
		.Z(to_acu[131]));
	notech_mux2 i_13326027(.S(n_61993), .A(to_acu0[132]), .B(to_acu1[132]), 
		.Z(to_acu[132]));
	notech_mux2 i_13426028(.S(n_61988), .A(to_acu0[133]), .B(to_acu1[133]), 
		.Z(to_acu[133]));
	notech_mux2 i_13526029(.S(n_61988), .A(to_acu0[134]), .B(to_acu1[134]), 
		.Z(to_acu[134]));
	notech_mux2 i_13626030(.S(n_61988), .A(to_acu0[135]), .B(to_acu1[135]), 
		.Z(to_acu[135]));
	notech_mux2 i_13726031(.S(n_61993), .A(to_acu0[136]), .B(to_acu1[136]), 
		.Z(to_acu[136]));
	notech_mux2 i_13826032(.S(n_61993), .A(to_acu0[137]), .B(to_acu1[137]), 
		.Z(to_acu[137]));
	notech_mux2 i_13926033(.S(n_61993), .A(to_acu0[138]), .B(to_acu1[138]), 
		.Z(to_acu[138]));
	notech_mux2 i_14026034(.S(n_61993), .A(to_acu0[139]), .B(to_acu1[139]), 
		.Z(to_acu[139]));
	notech_mux2 i_14126035(.S(n_61993), .A(to_acu0[140]), .B(to_acu1[140]), 
		.Z(to_acu[140]));
	notech_mux2 i_14226036(.S(n_61993), .A(to_acu0[141]), .B(to_acu1[141]), 
		.Z(to_acu[141]));
	notech_mux2 i_14326037(.S(n_61993), .A(to_acu0[142]), .B(to_acu1[142]), 
		.Z(to_acu[142]));
	notech_mux2 i_14426038(.S(n_61988), .A(to_acu0[143]), .B(to_acu1[143]), 
		.Z(to_acu[143]));
	notech_mux2 i_14526039(.S(n_61988), .A(to_acu0[144]), .B(to_acu1[144]), 
		.Z(to_acu[144]));
	notech_mux2 i_14626040(.S(n_61988), .A(to_acu0[145]), .B(to_acu1[145]), 
		.Z(to_acu[145]));
	notech_mux2 i_14726041(.S(n_61988), .A(to_acu0[146]), .B(to_acu1[146]), 
		.Z(to_acu[146]));
	notech_mux2 i_14826042(.S(n_61988), .A(to_acu0[147]), .B(to_acu1[147]), 
		.Z(to_acu[147]));
	notech_mux2 i_14926043(.S(n_61988), .A(to_acu0[148]), .B(to_acu1[148]), 
		.Z(to_acu[148]));
	notech_mux2 i_15026044(.S(n_61988), .A(to_acu0[149]), .B(to_acu1[149]), 
		.Z(to_acu[149]));
	notech_mux2 i_15126045(.S(n_61988), .A(to_acu0[150]), .B(to_acu1[150]), 
		.Z(to_acu[150]));
	notech_mux2 i_15226046(.S(n_61988), .A(to_acu0[151]), .B(to_acu1[151]), 
		.Z(to_acu[151]));
	notech_mux2 i_15326047(.S(n_61988), .A(to_acu0[152]), .B(to_acu1[152]), 
		.Z(to_acu[152]));
	notech_mux2 i_15426048(.S(n_61988), .A(to_acu0[153]), .B(to_acu1[153]), 
		.Z(to_acu[153]));
	notech_mux2 i_15526049(.S(n_61988), .A(to_acu0[154]), .B(to_acu1[154]), 
		.Z(to_acu[154]));
	notech_mux2 i_15626050(.S(n_61988), .A(to_acu0[155]), .B(to_acu1[155]), 
		.Z(to_acu[155]));
	notech_mux2 i_15726051(.S(n_62022), .A(to_acu0[156]), .B(to_acu1[156]), 
		.Z(to_acu[156]));
	notech_mux2 i_15826052(.S(n_62022), .A(to_acu0[157]), .B(to_acu1[157]), 
		.Z(to_acu[157]));
	notech_mux2 i_15926053(.S(n_62022), .A(to_acu0[158]), .B(to_acu1[158]), 
		.Z(to_acu[158]));
	notech_mux2 i_16026054(.S(n_62022), .A(to_acu0[159]), .B(to_acu1[159]), 
		.Z(to_acu[159]));
	notech_mux2 i_16126055(.S(n_62022), .A(to_acu0[160]), .B(to_acu1[160]), 
		.Z(to_acu[160]));
	notech_mux2 i_16226056(.S(n_62022), .A(to_acu0[161]), .B(to_acu1[161]), 
		.Z(to_acu[161]));
	notech_mux2 i_16326057(.S(n_62022), .A(to_acu0[162]), .B(to_acu1[162]), 
		.Z(to_acu[162]));
	notech_mux2 i_16426058(.S(n_62022), .A(to_acu0[163]), .B(to_acu1[163]), 
		.Z(to_acu[163]));
	notech_mux2 i_16526059(.S(n_62022), .A(to_acu0[164]), .B(to_acu1[164]), 
		.Z(to_acu[164]));
	notech_mux2 i_16626060(.S(n_62022), .A(to_acu0[165]), .B(to_acu1[165]), 
		.Z(to_acu[165]));
	notech_mux2 i_16726061(.S(n_62022), .A(to_acu0[166]), .B(to_acu1[166]), 
		.Z(to_acu[166]));
	notech_mux2 i_16826062(.S(n_62022), .A(to_acu0[167]), .B(to_acu1[167]), 
		.Z(to_acu[167]));
	notech_mux2 i_16926063(.S(n_62022), .A(to_acu0[168]), .B(to_acu1[168]), 
		.Z(to_acu[168]));
	notech_mux2 i_17026064(.S(n_62021), .A(to_acu0[169]), .B(to_acu1[169]), 
		.Z(to_acu[169]));
	notech_mux2 i_17126065(.S(n_62021), .A(to_acu0[170]), .B(to_acu1[170]), 
		.Z(to_acu[170]));
	notech_mux2 i_17226066(.S(n_62021), .A(to_acu0[171]), .B(to_acu1[171]), 
		.Z(to_acu[171]));
	notech_mux2 i_17326067(.S(n_62021), .A(to_acu0[172]), .B(to_acu1[172]), 
		.Z(to_acu[172]));
	notech_mux2 i_17426068(.S(n_62021), .A(to_acu0[173]), .B(to_acu1[173]), 
		.Z(to_acu[173]));
	notech_mux2 i_17526069(.S(n_62021), .A(to_acu0[174]), .B(to_acu1[174]), 
		.Z(to_acu[174]));
	notech_mux2 i_17626070(.S(n_62021), .A(to_acu0[175]), .B(to_acu1[175]), 
		.Z(to_acu[175]));
	notech_mux2 i_17726071(.S(n_62022), .A(to_acu0[176]), .B(to_acu1[176]), 
		.Z(to_acu[176]));
	notech_mux2 i_17826072(.S(n_62022), .A(to_acu0[177]), .B(to_acu1[177]), 
		.Z(to_acu[177]));
	notech_mux2 i_17926073(.S(n_62022), .A(to_acu0[178]), .B(to_acu1[178]), 
		.Z(to_acu[178]));
	notech_mux2 i_18026074(.S(n_62021), .A(to_acu0[179]), .B(to_acu1[179]), 
		.Z(to_acu[179]));
	notech_mux2 i_18126075(.S(n_62021), .A(to_acu0[180]), .B(to_acu1[180]), 
		.Z(to_acu[180]));
	notech_mux2 i_18226076(.S(n_62021), .A(to_acu0[181]), .B(to_acu1[181]), 
		.Z(to_acu[181]));
	notech_mux2 i_18326077(.S(n_62022), .A(to_acu0[182]), .B(to_acu1[182]), 
		.Z(to_acu[182]));
	notech_mux2 i_18426078(.S(n_62032), .A(to_acu0[183]), .B(to_acu1[183]), 
		.Z(to_acu[183]));
	notech_mux2 i_18526079(.S(n_62032), .A(to_acu0[184]), .B(to_acu1[184]), 
		.Z(to_acu[184]));
	notech_mux2 i_18626080(.S(n_62032), .A(to_acu0[185]), .B(to_acu1[185]), 
		.Z(to_acu[185]));
	notech_mux2 i_18726081(.S(n_62032), .A(to_acu0[186]), .B(to_acu1[186]), 
		.Z(to_acu[186]));
	notech_mux2 i_18826082(.S(n_62032), .A(to_acu0[187]), .B(to_acu1[187]), 
		.Z(to_acu[187]));
	notech_mux2 i_18926083(.S(n_62032), .A(to_acu0[188]), .B(to_acu1[188]), 
		.Z(to_acu[188]));
	notech_mux2 i_19026084(.S(n_62032), .A(to_acu0[189]), .B(to_acu1[189]), 
		.Z(to_acu[189]));
	notech_mux2 i_19126085(.S(n_62032), .A(to_acu0[190]), .B(to_acu1[190]), 
		.Z(to_acu[190]));
	notech_mux2 i_19226086(.S(n_62032), .A(to_acu0[191]), .B(to_acu1[191]), 
		.Z(to_acu[191]));
	notech_mux2 i_19326087(.S(n_62032), .A(to_acu0[192]), .B(to_acu1[192]), 
		.Z(to_acu[192]));
	notech_mux2 i_19426088(.S(n_62032), .A(to_acu0[193]), .B(to_acu1[193]), 
		.Z(to_acu[193]));
	notech_mux2 i_19526089(.S(n_62032), .A(to_acu0[194]), .B(to_acu1[194]), 
		.Z(to_acu[194]));
	notech_mux2 i_19626090(.S(n_62032), .A(to_acu0[195]), .B(to_acu1[195]), 
		.Z(to_acu[195]));
	notech_mux2 i_19726091(.S(n_62027), .A(to_acu0[196]), .B(to_acu1[196]), 
		.Z(to_acu[196]));
	notech_mux2 i_19826092(.S(n_62027), .A(to_acu0[197]), .B(to_acu1[197]), 
		.Z(to_acu[197]));
	notech_mux2 i_19926093(.S(n_62027), .A(to_acu0[198]), .B(to_acu1[198]), 
		.Z(to_acu[198]));
	notech_mux2 i_20026094(.S(n_62022), .A(to_acu0[199]), .B(to_acu1[199]), 
		.Z(to_acu[199]));
	notech_mux2 i_20126095(.S(n_62027), .A(to_acu0[200]), .B(to_acu1[200]), 
		.Z(to_acu[200]));
	notech_mux2 i_20226096(.S(n_62027), .A(to_acu0[201]), .B(to_acu1[201]), 
		.Z(to_acu[201]));
	notech_mux2 i_20326097(.S(n_62027), .A(to_acu0[202]), .B(to_acu1[202]), 
		.Z(to_acu[202]));
	notech_mux2 i_20426098(.S(n_62027), .A(to_acu0[203]), .B(to_acu1[203]), 
		.Z(to_acu[203]));
	notech_mux2 i_20526099(.S(n_62027), .A(to_acu0[204]), .B(to_acu1[204]), 
		.Z(to_acu[204]));
	notech_mux2 i_20626100(.S(n_62027), .A(to_acu0[205]), .B(to_acu1[205]), 
		.Z(to_acu[205]));
	notech_mux2 i_20726101(.S(n_62027), .A(to_acu0[206]), .B(to_acu1[206]), 
		.Z(to_acu[206]));
	notech_mux2 i_20826102(.S(n_62027), .A(to_acu0[207]), .B(to_acu1[207]), 
		.Z(to_acu[207]));
	notech_mux2 i_20926103(.S(n_62027), .A(to_acu0[208]), .B(to_acu1[208]), 
		.Z(to_acu[208]));
	notech_mux2 i_21026104(.S(n_62021), .A(to_acu0[209]), .B(to_acu1[209]), 
		.Z(to_acu[209]));
	notech_mux2 i_21126105(.S(n_62010), .A(to_acu0[210]), .B(to_acu1[210]), 
		.Z(to_acu[210]));
	notech_mux2 i_627199(.S(n_62010), .A(\over_seg0[5] ), .B(\over_seg1[5] )
		, .Z(over_seg[5]));
	notech_mux2 i_127596(.S(n_62010), .A(\imm0[0] ), .B(\imm1[0] ), .Z(immediate
		[0]));
	notech_mux2 i_227597(.S(n_62009), .A(\imm0[1] ), .B(\imm1[1] ), .Z(immediate
		[1]));
	notech_mux2 i_327598(.S(n_62009), .A(\imm0[2] ), .B(\imm1[2] ), .Z(immediate
		[2]));
	notech_mux2 i_427599(.S(n_62009), .A(\imm0[3] ), .B(\imm1[3] ), .Z(immediate
		[3]));
	notech_mux2 i_527600(.S(n_62010), .A(\imm0[4] ), .B(\imm1[4] ), .Z(immediate
		[4]));
	notech_mux2 i_627601(.S(n_62010), .A(\imm0[5] ), .B(\imm1[5] ), .Z(immediate
		[5]));
	notech_mux2 i_727602(.S(n_62010), .A(\imm0[6] ), .B(\imm1[6] ), .Z(immediate
		[6]));
	notech_mux2 i_827603(.S(n_62010), .A(\imm0[7] ), .B(\imm1[7] ), .Z(immediate
		[7]));
	notech_mux2 i_927604(.S(n_62010), .A(\imm0[8] ), .B(\imm1[8] ), .Z(immediate
		[8]));
	notech_mux2 i_1027605(.S(n_62010), .A(\imm0[9] ), .B(\imm1[9] ), .Z(immediate
		[9]));
	notech_mux2 i_1127606(.S(n_62010), .A(\imm0[10] ), .B(\imm1[10] ), .Z(immediate
		[10]));
	notech_mux2 i_1227607(.S(n_62009), .A(\imm0[11] ), .B(\imm1[11] ), .Z(immediate
		[11]));
	notech_mux2 i_1327608(.S(n_62009), .A(\imm0[12] ), .B(\imm1[12] ), .Z(immediate
		[12]));
	notech_mux2 i_1427609(.S(n_62009), .A(\imm0[13] ), .B(\imm1[13] ), .Z(immediate
		[13]));
	notech_mux2 i_1527610(.S(n_62009), .A(\imm0[14] ), .B(\imm1[14] ), .Z(immediate
		[14]));
	notech_mux2 i_1627611(.S(n_62009), .A(\imm0[15] ), .B(\imm1[15] ), .Z(immediate
		[15]));
	notech_mux2 i_1727612(.S(n_62009), .A(\imm0[16] ), .B(\imm1[16] ), .Z(immediate
		[16]));
	notech_mux2 i_1827613(.S(n_62009), .A(\imm0[17] ), .B(\imm1[17] ), .Z(immediate
		[17]));
	notech_mux2 i_1927614(.S(n_62009), .A(\imm0[18] ), .B(\imm1[18] ), .Z(immediate
		[18]));
	notech_mux2 i_2027615(.S(n_62009), .A(\imm0[19] ), .B(\imm1[19] ), .Z(immediate
		[19]));
	notech_mux2 i_2127616(.S(n_62009), .A(\imm0[20] ), .B(\imm1[20] ), .Z(immediate
		[20]));
	notech_mux2 i_2227617(.S(n_62009), .A(\imm0[21] ), .B(\imm1[21] ), .Z(immediate
		[21]));
	notech_mux2 i_2327618(.S(n_62009), .A(\imm0[22] ), .B(\imm1[22] ), .Z(immediate
		[22]));
	notech_mux2 i_2427619(.S(n_62009), .A(\imm0[23] ), .B(\imm1[23] ), .Z(immediate
		[23]));
	notech_mux2 i_2527620(.S(n_62010), .A(\imm0[24] ), .B(\imm1[24] ), .Z(immediate
		[24]));
	notech_mux2 i_2627621(.S(n_62016), .A(\imm0[25] ), .B(\imm1[25] ), .Z(immediate
		[25]));
	notech_mux2 i_2727622(.S(n_62016), .A(\imm0[26] ), .B(\imm1[26] ), .Z(immediate
		[26]));
	notech_mux2 i_2827623(.S(n_62016), .A(\imm0[27] ), .B(\imm1[27] ), .Z(immediate
		[27]));
	notech_mux2 i_2927624(.S(n_62016), .A(\imm0[28] ), .B(\imm1[28] ), .Z(immediate
		[28]));
	notech_mux2 i_3027625(.S(n_62016), .A(\imm0[29] ), .B(\imm1[29] ), .Z(immediate
		[29]));
	notech_mux2 i_3127626(.S(n_62016), .A(\imm0[30] ), .B(\imm1[30] ), .Z(immediate
		[30]));
	notech_mux2 i_3227627(.S(n_62021), .A(\imm0[31] ), .B(\imm1[31] ), .Z(immediate
		[31]));
	notech_mux2 i_3327628(.S(n_62021), .A(\imm0[32] ), .B(\imm1[32] ), .Z(immediate
		[32]));
	notech_mux2 i_3427629(.S(n_62021), .A(\imm0[33] ), .B(\imm1[33] ), .Z(immediate
		[33]));
	notech_mux2 i_3527630(.S(n_62021), .A(\imm0[34] ), .B(\imm1[34] ), .Z(immediate
		[34]));
	notech_mux2 i_3627631(.S(n_62021), .A(\imm0[35] ), .B(\imm1[35] ), .Z(immediate
		[35]));
	notech_mux2 i_3727632(.S(n_62021), .A(\imm0[36] ), .B(\imm1[36] ), .Z(immediate
		[36]));
	notech_mux2 i_3827633(.S(n_62021), .A(\imm0[37] ), .B(\imm1[37] ), .Z(immediate
		[37]));
	notech_mux2 i_3927634(.S(n_62010), .A(\imm0[38] ), .B(\imm1[38] ), .Z(immediate
		[38]));
	notech_mux2 i_4027635(.S(n_62010), .A(\imm0[39] ), .B(\imm1[39] ), .Z(immediate
		[39]));
	notech_mux2 i_4127636(.S(n_62010), .A(\imm0[40] ), .B(\imm1[40] ), .Z(immediate
		[40]));
	notech_mux2 i_4227637(.S(n_62010), .A(\imm0[41] ), .B(\imm1[41] ), .Z(immediate
		[41]));
	notech_mux2 i_4327638(.S(n_62010), .A(\imm0[42] ), .B(\imm1[42] ), .Z(immediate
		[42]));
	notech_mux2 i_4427639(.S(n_62010), .A(\imm0[43] ), .B(\imm1[43] ), .Z(immediate
		[43]));
	notech_mux2 i_4527640(.S(n_62010), .A(\imm0[44] ), .B(\imm1[44] ), .Z(immediate
		[44]));
	notech_mux2 i_4627641(.S(n_62016), .A(\imm0[45] ), .B(\imm1[45] ), .Z(immediate
		[45]));
	notech_mux2 i_4727642(.S(n_62016), .A(\imm0[46] ), .B(\imm1[46] ), .Z(immediate
		[46]));
	notech_mux2 i_4827643(.S(n_62016), .A(\imm0[47] ), .B(\imm1[47] ), .Z(immediate
		[47]));
	notech_nand3 i_6580661(.A(n_60932), .B(n_194199020), .C(n_16799552), .Z(\nbus_13544[0] 
		));
	notech_nand2 i_12580659(.A(n_5765), .B(n_16599551), .Z(n_42755));
	notech_nand2 i_430232(.A(cpl[0]), .B(cpl[1]), .Z(n_160356214));
	notech_ao4 i_69071(.A(n_1913), .B(n_44171), .C(n_60348), .D(n_44739), .Z
		(n_46130));
	notech_ao4 i_69075(.A(n_1913), .B(n_44174), .C(n_60348), .D(n_44761), .Z
		(n_46136));
	notech_ao4 i_69079(.A(n_1913), .B(n_44176), .C(n_60337), .D(n_44762), .Z
		(n_46142));
	notech_ao4 i_69083(.A(n_1913), .B(n_44179), .C(n_60337), .D(n_44763), .Z
		(n_46148));
	notech_ao4 i_69087(.A(n_1913), .B(n_44181), .C(n_60337), .D(n_44764), .Z
		(n_46154));
	notech_ao4 i_69091(.A(n_1913), .B(n_44183), .C(n_60337), .D(n_44765), .Z
		(n_46160));
	notech_ao4 i_1126116(.A(n_59197), .B(n_43491), .C(n_60232), .D(n_44752),
		 .Z(n_48498));
	notech_nand3 i_11425752(.A(n_1198100506), .B(n_12254735), .C(n_1178100486
		), .Z(n_45447));
	notech_nand3 i_7525713(.A(n_60932), .B(n_59129), .C(n_1200100508), .Z(n_45213
		));
	notech_nand3 i_6525703(.A(n_60932), .B(n_59129), .C(n_1201100509), .Z(n_45153
		));
	notech_nand2 i_6425702(.A(n_60932), .B(n_1202100510), .Z(n_45147));
	notech_nand3 i_6325701(.A(n_158456195), .B(n_60932), .C(n_1204100511), .Z
		(n_45141));
	notech_nand3 i_6225700(.A(n_59157), .B(n_60932), .C(n_1205100512), .Z(n_45135
		));
	notech_nand2 i_6125699(.A(n_60932), .B(n_1206100513), .Z(n_45129));
	notech_nand2 i_6025698(.A(n_60932), .B(n_1207100514), .Z(n_45123));
	notech_nand2 i_5825696(.A(n_60932), .B(n_1208100515), .Z(n_45111));
	notech_nao3 i_5725695(.A(n_60932), .B(n_1209100516), .C(n_1538), .Z(n_45105
		));
	notech_nand3 i_5525693(.A(n_60932), .B(n_1210100517), .C(n_59157), .Z(n_45093
		));
	notech_nao3 i_5425692(.A(n_60932), .B(n_1211100518), .C(n_1538), .Z(n_45087
		));
	notech_nand2 i_5325691(.A(n_60932), .B(n_1212100519), .Z(n_45081));
	notech_nand2 i_5225690(.A(n_60937), .B(n_1213100520), .Z(n_45075));
	notech_nand2 i_5025688(.A(n_60939), .B(n_1214100521), .Z(n_45063));
	notech_nand2 i_4925687(.A(n_60939), .B(n_1215100522), .Z(n_45057));
	notech_nand3 i_4625684(.A(n_60939), .B(n_59129), .C(n_1216100523), .Z(n_45039
		));
	notech_nand2 i_4525683(.A(n_60939), .B(n_1217100524), .Z(n_45033));
	notech_nao3 i_4325681(.A(n_60939), .B(n_1218100525), .C(n_1538), .Z(n_45021
		));
	notech_nand2 i_4225680(.A(n_60939), .B(n_1219100526), .Z(n_45015));
	notech_nand2 i_4125679(.A(n_60939), .B(n_1220100527), .Z(n_45009));
	notech_nand2 i_4025678(.A(n_60939), .B(n_1221100528), .Z(n_45003));
	notech_nand3 i_3925677(.A(n_60939), .B(n_59129), .C(n_1222100529), .Z(n_44997
		));
	notech_nand2 i_3725675(.A(n_60939), .B(n_1223100530), .Z(n_44985));
	notech_nand2 i_3625674(.A(n_60939), .B(n_1224100531), .Z(n_44979));
	notech_nand3 i_3525673(.A(n_60939), .B(n_59129), .C(n_1225100532), .Z(n_44973
		));
	notech_nand3 i_3425672(.A(n_60939), .B(n_1226100533), .C(n_59129), .Z(n_44967
		));
	notech_nand2 i_3225670(.A(n_60939), .B(n_1227100534), .Z(n_44955));
	notech_nand2 i_2425662(.A(n_60939), .B(n_1228100535), .Z(n_44907));
	notech_nand2 i_2325661(.A(n_60939), .B(n_1229100536), .Z(n_44901));
	notech_nand2 i_2025658(.A(n_60937), .B(n_1230100537), .Z(n_44883));
	notech_nand2 i_1925657(.A(n_60937), .B(n_1231100538), .Z(n_44877));
	notech_nand2 i_1725655(.A(n_60937), .B(n_1232100539), .Z(n_44865));
	notech_nand2 i_1525653(.A(n_60937), .B(n_1233100540), .Z(n_44853));
	notech_nand2 i_1425652(.A(n_60937), .B(n_1234100541), .Z(n_44847));
	notech_nand2 i_1325651(.A(n_60937), .B(n_1235100542), .Z(n_44841));
	notech_nand2 i_1225650(.A(n_60937), .B(n_1236100543), .Z(n_44835));
	notech_nand2 i_1125649(.A(n_60937), .B(n_1237100544), .Z(n_44829));
	notech_nand2 i_1025648(.A(n_60937), .B(n_1238100545), .Z(n_44823));
	notech_nand2 i_925647(.A(n_1239100546), .B(n_60937), .Z(n_44817));
	notech_ao4 i_18326499(.A(n_60232), .B(n_44624), .C(n_59197), .D(n_44108)
		, .Z(n_43864));
	notech_ao4 i_18226498(.A(n_60232), .B(n_44623), .C(n_59197), .D(n_44107)
		, .Z(n_43858));
	notech_ao4 i_18126497(.A(n_60232), .B(n_44622), .C(n_59197), .D(n_44104)
		, .Z(n_43852));
	notech_ao4 i_18026496(.A(n_60230), .B(n_44620), .C(n_59197), .D(n_44103)
		, .Z(n_43846));
	notech_ao4 i_17926495(.A(n_60227), .B(n_44619), .C(n_59197), .D(n_44102)
		, .Z(n_43840));
	notech_ao4 i_1926335(.A(n_60227), .B(n_44714), .C(n_59197), .D(n_43860),
		 .Z(n_42880));
	notech_ao4 i_1826334(.A(n_60227), .B(n_44715), .C(n_59197), .D(n_43859),
		 .Z(n_42874));
	notech_ao4 i_1726333(.A(n_60230), .B(n_44718), .C(n_59197), .D(n_43856),
		 .Z(n_42868));
	notech_ao4 i_1626332(.A(n_60230), .B(n_44711), .C(n_59197), .D(n_43854),
		 .Z(n_42862));
	notech_ao4 i_1526331(.A(n_60227), .B(n_44712), .C(n_59201), .D(n_43853),
		 .Z(n_42856));
	notech_ao4 i_1426330(.A(n_60227), .B(n_44713), .C(n_59201), .D(n_43850),
		 .Z(n_42850));
	notech_ao4 i_1326329(.A(n_60227), .B(n_44716), .C(n_59201), .D(n_43848),
		 .Z(n_42844));
	notech_ao4 i_1226328(.A(n_60227), .B(n_44727), .C(n_59201), .D(n_43847),
		 .Z(n_42838));
	notech_ao4 i_1126327(.A(n_59201), .B(n_43844), .C(n_60227), .D(n_44752),
		 .Z(n_42832));
	notech_ao4 i_1026326(.A(n_60230), .B(n_44728), .C(n_59197), .D(n_43842),
		 .Z(n_42826));
	notech_ao4 i_926325(.A(n_60230), .B(n_44726), .C(n_59197), .D(n_43839), 
		.Z(n_42820));
	notech_ao4 i_826324(.A(n_60230), .B(n_44759), .C(n_59197), .D(n_43837), 
		.Z(n_42814));
	notech_and2 i_780638(.A(n_1912), .B(n_44744), .Z(n_158456195));
	notech_ao4 i_502(.A(n_44157), .B(n_44710), .C(n_3078), .D(n_44557), .Z(n_3095
		));
	notech_and2 i_497(.A(n_3092), .B(n_2451), .Z(n_3093));
	notech_ao4 i_496(.A(n_3072), .B(n_44576), .C(n_3069), .D(n_44566), .Z(n_3092
		));
	notech_ao4 i_489(.A(n_44157), .B(n_44720), .C(n_3078), .D(n_44556), .Z(n_3090
		));
	notech_and2 i_484(.A(n_3087), .B(n_2443), .Z(n_3088));
	notech_ao4 i_483(.A(n_3072), .B(n_44575), .C(n_3069), .D(n_44565), .Z(n_3087
		));
	notech_ao4 i_476(.A(n_44157), .B(n_44723), .C(n_3078), .D(n_44554), .Z(n_3085
		));
	notech_and2 i_471(.A(n_3082), .B(n_2435), .Z(n_3083));
	notech_ao4 i_470(.A(n_3072), .B(n_44574), .C(n_3069), .D(n_44564), .Z(n_3082
		));
	notech_ao4 i_463(.A(n_44722), .B(n_44157), .C(n_44553), .D(n_3078), .Z(n_3080
		));
	notech_and2 i_21(.A(n_3060), .B(n_3077), .Z(n_3079));
	notech_or2 i_32(.A(n_3060), .B(n_44158), .Z(n_3078));
	notech_ao3 i_448(.A(n_3062), .B(n_44161), .C(n_3057), .Z(n_3077));
	notech_and4 i_18(.A(n_3062), .B(n_3057), .C(n_3060), .D(n_44161), .Z(n_3076
		));
	notech_nand2 i_75040(.A(n_1554100859), .B(n_2695), .Z(\nbus_13566[0] )
		);
	notech_nand3 i_6479049(.A(n_60937), .B(n_1481100787), .C(n_194199020), .Z
		(\nbus_13540[0] ));
	notech_nand2 i_9379048(.A(n_1554100859), .B(n_1240100547), .Z(\nbus_13546[0] 
		));
	notech_ao4 i_4625428(.A(n_60230), .B(n_44428), .C(n_59201), .D(n_42927),
		 .Z(n_50165));
	notech_ao4 i_4525427(.A(n_60230), .B(n_44427), .C(n_59201), .D(n_42925),
		 .Z(n_50159));
	notech_ao4 i_4425426(.A(n_60230), .B(n_44426), .C(n_59197), .D(n_42923),
		 .Z(n_50153));
	notech_ao4 i_4325425(.A(n_60230), .B(n_44425), .C(n_59195), .D(n_42920),
		 .Z(n_50147));
	notech_ao4 i_4225424(.A(n_60230), .B(n_44424), .C(n_59191), .D(n_42918),
		 .Z(n_50141));
	notech_ao4 i_925391(.A(n_60230), .B(n_44384), .C(n_59195), .D(n_42858), 
		.Z(n_49943));
	notech_ao4 i_825390(.A(n_60230), .B(n_44383), .C(n_59195), .D(n_42855), 
		.Z(n_49937));
	notech_ao4 i_625388(.A(n_60208), .B(n_44380), .C(n_59195), .D(n_42851), 
		.Z(n_49925));
	notech_ao4 i_125383(.A(n_60208), .B(n_44374), .C(n_59191), .D(n_42841), 
		.Z(n_49895));
	notech_mux2 i_828067(.S(n_1554100859), .A(ififo_rvect4[7]), .B(ififo_rvect2
		[7]), .Z(n_46080));
	notech_mux2 i_728066(.S(n_1554100859), .A(ififo_rvect4[6]), .B(ififo_rvect2
		[6]), .Z(n_46074));
	notech_mux2 i_628065(.S(n_1554100859), .A(ififo_rvect4[5]), .B(ififo_rvect2
		[5]), .Z(n_46068));
	notech_mux2 i_528064(.S(n_1554100859), .A(ififo_rvect4[4]), .B(ififo_rvect2
		[4]), .Z(n_46062));
	notech_mux2 i_428063(.S(n_1554100859), .A(ififo_rvect4[3]), .B(ififo_rvect2
		[3]), .Z(n_46056));
	notech_mux2 i_328062(.S(n_1554100859), .A(ififo_rvect4[2]), .B(ififo_rvect2
		[2]), .Z(n_46050));
	notech_mux2 i_228061(.S(n_1554100859), .A(ififo_rvect4[1]), .B(ififo_rvect2
		[1]), .Z(n_46044));
	notech_mux2 i_128060(.S(n_56813), .A(ififo_rvect4[0]), .B(ififo_rvect2[0
		]), .Z(n_46038));
	notech_mux2 i_828027(.S(n_56813), .A(ififo_rvect3[7]), .B(ififo_rvect1[7
		]), .Z(n_48403));
	notech_mux2 i_728026(.S(n_56813), .A(ififo_rvect3[6]), .B(ififo_rvect1[6
		]), .Z(n_48397));
	notech_mux2 i_628025(.S(n_56813), .A(ififo_rvect3[5]), .B(ififo_rvect1[5
		]), .Z(n_48391));
	notech_mux2 i_528024(.S(n_56813), .A(ififo_rvect3[4]), .B(ififo_rvect1[4
		]), .Z(n_48385));
	notech_mux2 i_428023(.S(n_56813), .A(ififo_rvect3[3]), .B(ififo_rvect1[3
		]), .Z(n_48379));
	notech_mux2 i_328022(.S(n_56813), .A(ififo_rvect3[2]), .B(ififo_rvect1[2
		]), .Z(n_48373));
	notech_mux2 i_228021(.S(n_56813), .A(ififo_rvect3[1]), .B(ififo_rvect1[1
		]), .Z(n_48367));
	notech_mux2 i_128020(.S(n_56813), .A(ififo_rvect3[0]), .B(ififo_rvect1[0
		]), .Z(n_48361));
	notech_mux2 i_828035(.S(n_56813), .A(ififo_rvect2[7]), .B(ivect[7]), .Z(n_44334
		));
	notech_mux2 i_728034(.S(n_56813), .A(ififo_rvect2[6]), .B(ivect[6]), .Z(n_44328
		));
	notech_mux2 i_628033(.S(n_1554100859), .A(ififo_rvect2[5]), .B(ivect[5])
		, .Z(n_44322));
	notech_mux2 i_528032(.S(n_56813), .A(ififo_rvect2[4]), .B(ivect[4]), .Z(n_44316
		));
	notech_mux2 i_428031(.S(n_56813), .A(ififo_rvect2[3]), .B(ivect[3]), .Z(n_44310
		));
	notech_mux2 i_328030(.S(n_56813), .A(ififo_rvect2[2]), .B(ivect[2]), .Z(n_44304
		));
	notech_mux2 i_228029(.S(n_56813), .A(ififo_rvect2[1]), .B(ivect[1]), .Z(n_44298
		));
	notech_mux2 i_128028(.S(n_56813), .A(ififo_rvect2[0]), .B(ivect[0]), .Z(n_44292
		));
	notech_ao4 i_21026315(.A(n_60208), .B(n_44656), .C(n_59191), .D(n_43824)
		, .Z(n_49692));
	notech_ao4 i_20826313(.A(n_60209), .B(n_44654), .C(n_59191), .D(n_43821)
		, .Z(n_49680));
	notech_ao4 i_19326298(.A(n_60208), .B(n_44636), .C(n_59191), .D(n_43801)
		, .Z(n_49590));
	notech_ao4 i_19226297(.A(n_60208), .B(n_44635), .C(n_59191), .D(n_43800)
		, .Z(n_49584));
	notech_ao4 i_19126296(.A(n_60208), .B(n_44634), .C(n_59195), .D(n_43799)
		, .Z(n_49578));
	notech_ao4 i_12526230(.A(n_60208), .B(n_44554), .C(n_59195), .D(n_43664)
		, .Z(n_49182));
	notech_ao4 i_12326228(.A(n_60208), .B(n_44552), .C(n_59195), .D(n_43659)
		, .Z(n_49170));
	notech_ao4 i_12226227(.A(n_60208), .B(n_44551), .C(n_59195), .D(n_43657)
		, .Z(n_49164));
	notech_ao4 i_12126226(.A(n_60209), .B(n_44550), .C(n_59195), .D(n_43655)
		, .Z(n_49158));
	notech_ao4 i_12026225(.A(n_60209), .B(n_44548), .C(n_59195), .D(n_43652)
		, .Z(n_49152));
	notech_ao4 i_11926224(.A(n_60209), .B(n_44547), .C(n_59195), .D(n_43650)
		, .Z(n_49146));
	notech_ao4 i_11826223(.A(n_60209), .B(n_44546), .C(n_59195), .D(n_43647)
		, .Z(n_49140));
	notech_ao4 i_11726222(.A(n_60209), .B(n_44545), .C(n_59195), .D(n_43645)
		, .Z(n_49134));
	notech_ao4 i_11626221(.A(n_60209), .B(n_44544), .C(n_59195), .D(n_43643)
		, .Z(n_49128));
	notech_ao4 i_11526220(.A(n_60209), .B(n_44542), .C(n_59184), .D(n_43640)
		, .Z(n_49122));
	notech_ao4 i_11326218(.A(n_60209), .B(n_44540), .C(n_59173), .D(n_43635)
		, .Z(n_49110));
	notech_ao4 i_11226217(.A(n_60209), .B(n_44539), .C(n_59173), .D(n_43633)
		, .Z(n_49104));
	notech_ao4 i_11126216(.A(n_60209), .B(n_44538), .C(n_59173), .D(n_43631)
		, .Z(n_49098));
	notech_ao4 i_11026215(.A(n_60208), .B(n_44536), .C(n_59174), .D(n_43628)
		, .Z(n_49092));
	notech_ao4 i_10926214(.A(n_60203), .B(n_44535), .C(n_59173), .D(n_43626)
		, .Z(n_49086));
	notech_ao4 i_10826213(.A(n_60203), .B(n_44534), .C(n_59174), .D(n_43625)
		, .Z(n_49080));
	notech_ao4 i_10626211(.A(n_60203), .B(n_44532), .C(n_59174), .D(n_43622)
		, .Z(n_49068));
	notech_ao4 i_10426209(.A(n_60203), .B(n_44529), .C(n_59174), .D(n_43620)
		, .Z(n_49056));
	notech_ao4 i_10326208(.A(n_60203), .B(n_44528), .C(n_59173), .D(n_43619)
		, .Z(n_49050));
	notech_ao4 i_10126206(.A(n_60203), .B(n_44526), .C(n_59173), .D(n_43616)
		, .Z(n_49038));
	notech_ao4 i_10026205(.A(n_60203), .B(n_44525), .C(n_59173), .D(n_43615)
		, .Z(n_49032));
	notech_ao4 i_4626151(.A(n_60203), .B(n_44750), .C(n_59174), .D(n_43549),
		 .Z(n_48708));
	notech_ao4 i_4226147(.A(n_60203), .B(n_44749), .C(n_59173), .D(n_43544),
		 .Z(n_48684));
	notech_ao4 i_3126136(.A(n_60203), .B(n_44767), .C(n_59173), .D(n_43531),
		 .Z(n_48618));
	notech_ao4 i_3026135(.A(n_60208), .B(n_44766), .C(n_59173), .D(n_43529),
		 .Z(n_48612));
	notech_ao4 i_2926134(.A(n_60208), .B(n_44757), .C(n_59174), .D(n_43527),
		 .Z(n_48606));
	notech_ao4 i_2826133(.A(n_60208), .B(n_44746), .C(n_59174), .D(n_43526),
		 .Z(n_48600));
	notech_ao4 i_2726132(.A(n_60208), .B(n_44743), .C(n_59174), .D(n_43525),
		 .Z(n_48594));
	notech_ao4 i_2626131(.A(n_60208), .B(n_44755), .C(n_59174), .D(n_43523),
		 .Z(n_48588));
	notech_ao4 i_2526130(.A(n_60203), .B(n_44756), .C(n_59174), .D(n_43520),
		 .Z(n_48582));
	notech_ao4 i_2426129(.A(n_60203), .B(n_44741), .C(n_59174), .D(n_43518),
		 .Z(n_48576));
	notech_ao4 i_2326128(.A(n_60208), .B(n_44740), .C(n_59168), .D(n_43515),
		 .Z(n_48570));
	notech_ao4 i_2226127(.A(n_60208), .B(n_44742), .C(n_59168), .D(n_43513),
		 .Z(n_48564));
	notech_ao4 i_2126126(.A(n_60208), .B(n_44754), .C(n_59168), .D(n_43511),
		 .Z(n_48558));
	notech_ao4 i_2026125(.A(n_60209), .B(n_44753), .C(n_59168), .D(n_43508),
		 .Z(n_48552));
	notech_ao4 i_622110(.A(n_60216), .B(n_44765), .C(n_59168), .D(n_44156), 
		.Z(n_44088));
	notech_ao4 i_522109(.A(n_60216), .B(n_44764), .C(n_59168), .D(n_44155), 
		.Z(n_44082));
	notech_ao4 i_422108(.A(n_60216), .B(n_44763), .C(n_59168), .D(n_44153), 
		.Z(n_44076));
	notech_ao4 i_322107(.A(n_60216), .B(n_44762), .C(n_59168), .D(n_44152), 
		.Z(n_44070));
	notech_ao4 i_222106(.A(n_60216), .B(n_44761), .C(n_59168), .D(n_44151), 
		.Z(n_44064));
	notech_ao4 i_21026526(.A(n_60216), .B(n_44656), .C(n_59168), .D(n_44146)
		, .Z(n_44026));
	notech_ao4 i_20926525(.A(n_60216), .B(n_44655), .C(n_59174), .D(n_44144)
		, .Z(n_44020));
	notech_ao4 i_20826524(.A(n_60216), .B(n_44654), .C(n_59174), .D(n_44143)
		, .Z(n_44014));
	notech_ao4 i_20726523(.A(n_60216), .B(n_44653), .C(n_59174), .D(n_44140)
		, .Z(n_44008));
	notech_ao4 i_20626522(.A(n_60216), .B(n_44652), .C(n_59174), .D(n_44139)
		, .Z(n_44002));
	notech_ao4 i_20526521(.A(n_60219), .B(n_44650), .C(n_59174), .D(n_44138)
		, .Z(n_43996));
	notech_ao4 i_20426520(.A(n_60219), .B(n_44649), .C(n_59168), .D(n_44137)
		, .Z(n_43990));
	notech_ao4 i_20326519(.A(n_60219), .B(n_44648), .C(n_59168), .D(n_44135)
		, .Z(n_43984));
	notech_ao4 i_20226518(.A(n_60219), .B(n_44647), .C(n_59174), .D(n_44134)
		, .Z(n_43978));
	notech_ao4 i_20126517(.A(n_60219), .B(n_44646), .C(n_59174), .D(n_44133)
		, .Z(n_43972));
	notech_ao4 i_20026516(.A(n_60216), .B(n_44644), .C(n_59174), .D(n_44132)
		, .Z(n_43966));
	notech_ao4 i_19926515(.A(n_60216), .B(n_44643), .C(n_59180), .D(n_44131)
		, .Z(n_43960));
	notech_ao4 i_19826514(.A(n_60216), .B(n_44642), .C(n_59180), .D(n_44129)
		, .Z(n_43954));
	notech_ao4 i_19726513(.A(n_60219), .B(n_44641), .C(n_59180), .D(n_44128)
		, .Z(n_43948));
	notech_ao4 i_19626512(.A(n_60216), .B(n_44640), .C(n_59180), .D(n_44127)
		, .Z(n_43942));
	notech_ao4 i_19526511(.A(n_60214), .B(n_44638), .C(n_59180), .D(n_44126)
		, .Z(n_43936));
	notech_ao4 i_19426510(.A(n_60209), .B(n_44637), .C(n_59180), .D(n_44125)
		, .Z(n_43930));
	notech_ao4 i_19326509(.A(n_60209), .B(n_44636), .C(n_59180), .D(n_44123)
		, .Z(n_43924));
	notech_ao4 i_19226508(.A(n_60214), .B(n_44635), .C(n_59180), .D(n_44121)
		, .Z(n_43918));
	notech_ao4 i_19126507(.A(n_60214), .B(n_44634), .C(n_59180), .D(n_44119)
		, .Z(n_43912));
	notech_ao4 i_19026506(.A(n_60214), .B(n_44632), .C(n_59180), .D(n_44116)
		, .Z(n_43906));
	notech_ao4 i_18926505(.A(n_60209), .B(n_44631), .C(n_59184), .D(n_44115)
		, .Z(n_43900));
	notech_ao4 i_18826504(.A(n_60209), .B(n_44630), .C(n_59184), .D(n_44114)
		, .Z(n_43894));
	notech_ao4 i_18726503(.A(n_60209), .B(n_44629), .C(n_59184), .D(n_44113)
		, .Z(n_43888));
	notech_ao4 i_18626502(.A(n_60209), .B(n_44628), .C(n_59184), .D(n_44111)
		, .Z(n_43882));
	notech_ao4 i_18526501(.A(n_60209), .B(n_44626), .C(n_59184), .D(n_44110)
		, .Z(n_43876));
	notech_ao4 i_18426500(.A(n_60214), .B(n_44625), .C(n_59184), .D(n_44109)
		, .Z(n_43870));
	notech_ao4 i_17826494(.A(n_60214), .B(n_44618), .C(n_59184), .D(n_44101)
		, .Z(n_43834));
	notech_ao4 i_17726493(.A(n_60214), .B(n_44617), .C(n_59184), .D(n_44099)
		, .Z(n_43828));
	notech_ao4 i_17626492(.A(n_60214), .B(n_44616), .C(n_59184), .D(n_44098)
		, .Z(n_43822));
	notech_ao4 i_17526491(.A(n_60214), .B(n_44614), .C(n_59184), .D(n_44097)
		, .Z(n_43816));
	notech_ao4 i_17426490(.A(n_60214), .B(n_44613), .C(n_59180), .D(n_44096)
		, .Z(n_43810));
	notech_ao4 i_17326489(.A(n_60214), .B(n_44612), .C(n_59173), .D(n_44095)
		, .Z(n_43804));
	notech_ao4 i_17226488(.A(n_60214), .B(n_44611), .C(n_59173), .D(n_44093)
		, .Z(n_43798));
	notech_ao4 i_17126487(.A(n_60214), .B(n_44610), .C(n_59173), .D(n_44092)
		, .Z(n_43792));
	notech_ao4 i_17026486(.A(n_60214), .B(n_44608), .C(n_59173), .D(n_44091)
		, .Z(n_43786));
	notech_ao4 i_16926485(.A(n_60259), .B(n_44607), .C(n_59173), .D(n_44090)
		, .Z(n_43780));
	notech_ao4 i_16826484(.A(n_60259), .B(n_44606), .C(n_59173), .D(n_44089)
		, .Z(n_43774));
	notech_ao4 i_16726483(.A(n_60259), .B(n_44605), .C(n_59173), .D(n_44087)
		, .Z(n_43768));
	notech_ao4 i_16626482(.A(n_60259), .B(n_44604), .C(n_59173), .D(n_44086)
		, .Z(n_43762));
	notech_ao4 i_16526481(.A(n_60259), .B(n_44602), .C(n_59173), .D(n_44085)
		, .Z(n_43756));
	notech_ao4 i_16426480(.A(n_60255), .B(n_44601), .C(n_59173), .D(n_44084)
		, .Z(n_43750));
	notech_ao4 i_16326479(.A(n_60255), .B(n_44600), .C(n_59168), .D(n_44083)
		, .Z(n_43744));
	notech_ao4 i_16226478(.A(n_60255), .B(n_44599), .C(n_59168), .D(n_44081)
		, .Z(n_43738));
	notech_ao4 i_16126477(.A(n_60259), .B(n_44598), .C(n_59180), .D(n_44080)
		, .Z(n_43732));
	notech_ao4 i_16026476(.A(n_60259), .B(n_44596), .C(n_59180), .D(n_44079)
		, .Z(n_43726));
	notech_ao4 i_15926475(.A(n_60259), .B(n_44595), .C(n_59180), .D(n_44078)
		, .Z(n_43720));
	notech_ao4 i_15826474(.A(n_60259), .B(n_44594), .C(n_59168), .D(n_44077)
		, .Z(n_43714));
	notech_ao4 i_15726473(.A(n_60261), .B(n_44593), .C(n_59168), .D(n_44075)
		, .Z(n_43708));
	notech_ao4 i_15626472(.A(n_60261), .B(n_44592), .C(n_59168), .D(n_44074)
		, .Z(n_43702));
	notech_ao4 i_15526471(.A(n_60261), .B(n_44590), .C(n_59168), .D(n_44073)
		, .Z(n_43696));
	notech_ao4 i_15426470(.A(n_60259), .B(n_44589), .C(n_59168), .D(n_44072)
		, .Z(n_43690));
	notech_ao4 i_15326469(.A(n_60259), .B(n_44588), .C(n_59201), .D(n_44071)
		, .Z(n_43684));
	notech_ao4 i_15226468(.A(n_60259), .B(n_44587), .C(n_59224), .D(n_44069)
		, .Z(n_43678));
	notech_ao4 i_15126467(.A(n_60259), .B(n_44586), .C(n_59224), .D(n_44068)
		, .Z(n_43672));
	notech_ao4 i_15026466(.A(n_60259), .B(n_44584), .C(n_59224), .D(n_44067)
		, .Z(n_43666));
	notech_ao4 i_14926465(.A(n_60255), .B(n_44583), .C(n_59224), .D(n_44066)
		, .Z(n_43660));
	notech_ao4 i_14826464(.A(n_60253), .B(n_44582), .C(n_59224), .D(n_44065)
		, .Z(n_43654));
	notech_ao4 i_14726463(.A(n_60253), .B(n_44581), .C(n_59224), .D(n_44063)
		, .Z(n_43648));
	notech_ao4 i_14626462(.A(n_60253), .B(n_44580), .C(n_59224), .D(n_44062)
		, .Z(n_43642));
	notech_ao4 i_14526461(.A(n_60253), .B(n_44578), .C(n_59224), .D(n_44061)
		, .Z(n_43636));
	notech_ao4 i_14426460(.A(n_60253), .B(n_44577), .C(n_59224), .D(n_44060)
		, .Z(n_43630));
	notech_ao4 i_14326459(.A(n_60253), .B(n_44576), .C(n_59224), .D(n_44059)
		, .Z(n_43624));
	notech_ao4 i_14226458(.A(n_60253), .B(n_44575), .C(n_59226), .D(n_44057)
		, .Z(n_43618));
	notech_ao4 i_14126457(.A(n_60253), .B(n_44574), .C(n_59226), .D(n_44056)
		, .Z(n_43612));
	notech_ao4 i_14026456(.A(n_60253), .B(n_44572), .C(n_59226), .D(n_44055)
		, .Z(n_43606));
	notech_ao4 i_13926455(.A(n_60253), .B(n_44571), .C(n_59226), .D(n_44054)
		, .Z(n_43600));
	notech_ao4 i_13826454(.A(n_60255), .B(n_44570), .C(n_59226), .D(n_44053)
		, .Z(n_43594));
	notech_ao4 i_13726453(.A(n_60255), .B(n_44569), .C(n_59224), .D(n_44052)
		, .Z(n_43588));
	notech_ao4 i_13626452(.A(n_60255), .B(n_44568), .C(n_59224), .D(n_44051)
		, .Z(n_43582));
	notech_ao4 i_13426450(.A(n_60255), .B(n_44565), .C(n_59224), .D(n_44049)
		, .Z(n_43570));
	notech_ao4 i_13326449(.A(n_60255), .B(n_44564), .C(n_59226), .D(n_44048)
		, .Z(n_43564));
	notech_ao4 i_13226448(.A(n_60255), .B(n_44563), .C(n_59224), .D(n_44047)
		, .Z(n_43558));
	notech_ao4 i_13126447(.A(n_60255), .B(n_44562), .C(n_59220), .D(n_44046)
		, .Z(n_43552));
	notech_ao4 i_13026446(.A(n_60255), .B(n_44560), .C(n_59218), .D(n_44045)
		, .Z(n_43546));
	notech_ao4 i_12926445(.A(n_60255), .B(n_44559), .C(n_59218), .D(n_44043)
		, .Z(n_43540));
	notech_ao4 i_12826444(.A(n_60255), .B(n_44558), .C(n_59220), .D(n_44042)
		, .Z(n_43534));
	notech_ao4 i_12726443(.A(n_60261), .B(n_44557), .C(n_59220), .D(n_44040)
		, .Z(n_43528));
	notech_ao4 i_12626442(.A(n_60266), .B(n_44556), .C(n_59220), .D(n_44039)
		, .Z(n_43522));
	notech_ao4 i_12526441(.A(n_60266), .B(n_44554), .C(n_59218), .D(n_44038)
		, .Z(n_43516));
	notech_ao4 i_11126427(.A(n_60266), .B(n_44538), .C(n_59218), .D(n_44007)
		, .Z(n_43432));
	notech_ao4 i_10926425(.A(n_60266), .B(n_44535), .C(n_59218), .D(n_44003)
		, .Z(n_43420));
	notech_ao4 i_10726423(.A(n_60266), .B(n_44533), .C(n_59218), .D(n_43998)
		, .Z(n_43408));
	notech_ao4 i_10026416(.A(n_60264), .B(n_44525), .C(n_59218), .D(n_43985)
		, .Z(n_43366));
	notech_ao4 i_9926415(.A(n_60264), .B(n_44719), .C(n_59220), .D(n_43982),
		 .Z(n_43360));
	notech_ao4 i_9826414(.A(n_60264), .B(n_44721), .C(n_59220), .D(n_43981),
		 .Z(n_43354));
	notech_ao4 i_9226408(.A(n_60266), .B(n_44722), .C(n_59220), .D(n_43974),
		 .Z(n_43318));
	notech_ao4 i_9126407(.A(n_60266), .B(n_44674), .C(n_59220), .D(n_43973),
		 .Z(n_43312));
	notech_ao4 i_9026406(.A(n_60266), .B(n_44675), .C(n_59220), .D(n_43971),
		 .Z(n_43306));
	notech_ao4 i_8926405(.A(n_60266), .B(n_44676), .C(n_59220), .D(n_43970),
		 .Z(n_43300));
	notech_ao4 i_8826404(.A(n_60270), .B(n_44677), .C(n_59220), .D(n_43969),
		 .Z(n_43294));
	notech_ao4 i_8726403(.A(n_60270), .B(n_44678), .C(n_59220), .D(n_43968),
		 .Z(n_43288));
	notech_ao4 i_8626402(.A(n_60270), .B(n_44737), .C(n_59220), .D(n_43967),
		 .Z(n_43282));
	notech_ao4 i_8426400(.A(n_60266), .B(n_44659), .C(n_59220), .D(n_43964),
		 .Z(n_43270));
	notech_ao4 i_8326399(.A(n_60266), .B(n_44731), .C(n_59231), .D(n_43963),
		 .Z(n_43264));
	notech_ao4 i_8226398(.A(n_60266), .B(n_44730), .C(n_59231), .D(n_43962),
		 .Z(n_43258));
	notech_ao4 i_8126397(.A(n_60266), .B(n_44679), .C(n_59231), .D(n_43961),
		 .Z(n_43252));
	notech_ao4 i_8026396(.A(n_60266), .B(n_44705), .C(n_59231), .D(n_43959),
		 .Z(n_43246));
	notech_ao4 i_7926395(.A(n_60264), .B(n_44707), .C(n_59231), .D(n_43958),
		 .Z(n_43240));
	notech_ao4 i_7826394(.A(n_60261), .B(n_44660), .C(n_59231), .D(n_43957),
		 .Z(n_43234));
	notech_ao4 i_7726393(.A(n_60261), .B(n_44682), .C(n_59229), .D(n_43956),
		 .Z(n_43228));
	notech_ao4 i_7626392(.A(n_60261), .B(n_44673), .C(n_59231), .D(n_43955),
		 .Z(n_43222));
	notech_ao4 i_7526391(.A(n_60261), .B(n_44685), .C(n_59231), .D(n_43953),
		 .Z(n_43216));
	notech_ao4 i_7426390(.A(n_60261), .B(n_44684), .C(n_59231), .D(n_43952),
		 .Z(n_43210));
	notech_ao4 i_7326389(.A(n_60261), .B(n_44683), .C(n_59235), .D(n_43951),
		 .Z(n_43204));
	notech_ao4 i_7226388(.A(n_60261), .B(n_44671), .C(n_59235), .D(n_43950),
		 .Z(n_43198));
	notech_ao4 i_7126387(.A(n_60261), .B(n_44672), .C(n_59235), .D(n_43949),
		 .Z(n_43192));
	notech_ao4 i_7026386(.A(n_60261), .B(n_44725), .C(n_59235), .D(n_43947),
		 .Z(n_43186));
	notech_ao4 i_6926385(.A(n_60261), .B(n_44717), .C(n_59235), .D(n_43946),
		 .Z(n_43180));
	notech_ao4 i_6826384(.A(n_60264), .B(n_44661), .C(n_59231), .D(n_43945),
		 .Z(n_43174));
	notech_ao4 i_6626382(.A(n_60264), .B(n_44662), .C(n_59231), .D(n_43943),
		 .Z(n_43162));
	notech_ao4 i_6526381(.A(n_60264), .B(n_44663), .C(n_59231), .D(n_43941),
		 .Z(n_43156));
	notech_ao4 i_6326379(.A(n_60264), .B(n_44724), .C(n_59231), .D(n_43939),
		 .Z(n_43144));
	notech_ao4 i_6026376(.A(n_60264), .B(n_44692), .C(n_59231), .D(n_43935),
		 .Z(n_43126));
	notech_ao4 i_5926375(.A(n_60264), .B(n_44686), .C(n_59229), .D(n_43934),
		 .Z(n_43120));
	notech_ao4 i_5426370(.A(n_60264), .B(n_44690), .C(n_59226), .D(n_43928),
		 .Z(n_43090));
	notech_ao4 i_4926365(.A(n_60264), .B(n_44693), .C(n_59226), .D(n_43922),
		 .Z(n_43060));
	notech_ao4 i_4826364(.A(n_60264), .B(n_44704), .C(n_59226), .D(n_43921),
		 .Z(n_43054));
	notech_ao4 i_4726363(.A(n_60264), .B(n_44703), .C(n_59229), .D(n_43920),
		 .Z(n_43048));
	notech_ao4 i_4626362(.A(n_60241), .B(n_44750), .C(n_59229), .D(n_43919),
		 .Z(n_43042));
	notech_ao4 i_4526361(.A(n_60241), .B(n_44702), .C(n_59226), .D(n_43916),
		 .Z(n_43036));
	notech_ao4 i_4426360(.A(n_60241), .B(n_44700), .C(n_59226), .D(n_43915),
		 .Z(n_43030));
	notech_ao4 i_4326359(.A(n_60241), .B(n_44701), .C(n_59226), .D(n_43914),
		 .Z(n_43024));
	notech_ao4 i_3926355(.A(n_60241), .B(n_44699), .C(n_59226), .D(n_43908),
		 .Z(n_43000));
	notech_ao4 i_3826354(.A(n_60238), .B(n_44696), .C(n_59226), .D(n_43907),
		 .Z(n_42994));
	notech_ao4 i_3726353(.A(n_60238), .B(n_44697), .C(n_59229), .D(n_43904),
		 .Z(n_42988));
	notech_ao4 i_3626352(.A(n_60241), .B(n_44694), .C(n_59229), .D(n_43902),
		 .Z(n_42982));
	notech_ao4 i_3326349(.A(n_60241), .B(n_44664), .C(n_59229), .D(n_43896),
		 .Z(n_42964));
	notech_ao4 i_3226348(.A(n_60241), .B(n_44665), .C(n_59229), .D(n_43895),
		 .Z(n_42958));
	notech_ao4 i_3126347(.A(n_60243), .B(n_44767), .C(n_59229), .D(n_43892),
		 .Z(n_42952));
	notech_ao4 i_3026346(.A(n_60241), .B(n_44766), .C(n_59229), .D(n_43890),
		 .Z(n_42946));
	notech_ao4 i_2126337(.A(n_60243), .B(n_44754), .C(n_59229), .D(n_43866),
		 .Z(n_42892));
	notech_ao3 i_3579006(.A(n_60831), .B(in128[37]), .C(n_60337), .Z(n_83054515
		));
	notech_ao3 i_3679005(.A(n_60836), .B(in128[33]), .C(n_60337), .Z(n_82954514
		));
	notech_ao3 i_3779004(.A(n_60836), .B(in128[81]), .C(n_60337), .Z(n_82854513
		));
	notech_ao3 i_3879003(.A(n_60836), .B(in128[65]), .C(n_60337), .Z(n_82754512
		));
	notech_ao3 i_3979002(.A(n_60836), .B(in128[29]), .C(n_60337), .Z(n_82654511
		));
	notech_ao3 i_4079001(.A(n_60836), .B(in128[77]), .C(n_60337), .Z(n_82554510
		));
	notech_ao3 i_4179000(.A(n_60836), .B(in128[61]), .C(n_60337), .Z(n_82454509
		));
	notech_ao3 i_4278999(.A(n_60825), .B(in128[30]), .C(n_60372), .Z(n_82354508
		));
	notech_ao3 i_4378998(.A(n_60825), .B(in128[38]), .C(n_60372), .Z(n_82254507
		));
	notech_ao3 i_4478997(.A(n_60825), .B(in128[62]), .C(n_60372), .Z(n_82154506
		));
	notech_ao3 i_4578996(.A(n_60825), .B(in128[70]), .C(n_60372), .Z(n_82054505
		));
	notech_ao3 i_4678995(.A(n_60825), .B(in128[46]), .C(n_60372), .Z(n_81954504
		));
	notech_ao3 i_4778994(.A(n_60825), .B(in128[54]), .C(n_60372), .Z(n_81854503
		));
	notech_ao3 i_4878993(.A(n_60825), .B(in128[22]), .C(n_60376), .Z(n_81754502
		));
	notech_ao3 i_4978992(.A(n_60825), .B(in128[21]), .C(n_60376), .Z(n_81654501
		));
	notech_ao3 i_5178990(.A(n_60825), .B(in128[17]), .C(n_60376), .Z(n_81454499
		));
	notech_ao3 i_5378988(.A(n_60825), .B(in128[82]), .C(n_60376), .Z(n_81254497
		));
	notech_ao3 i_5678985(.A(n_60825), .B(in128[83]), .C(n_60376), .Z(n_80954494
		));
	notech_ao3 i_5978982(.A(n_60825), .B(\to_acu2_0[26] ), .C(n_60372), .Z(n_80654491
		));
	notech_ao3 i_6078981(.A(n_60825), .B(in128[23]), .C(n_60372), .Z(n_80554490
		));
	notech_ao3 i_6278979(.A(n_60847), .B(in128[86]), .C(n_60371), .Z(n_80354488
		));
	notech_ao3 i_6378978(.A(n_60860), .B(in128[84]), .C(n_60371), .Z(n_80254487
		));
	notech_ao3 i_6578977(.A(n_60860), .B(in128[80]), .C(n_60371), .Z(n_80154486
		));
	notech_ao3 i_6678976(.A(n_60865), .B(in128[79]), .C(n_60372), .Z(n_80054485
		));
	notech_ao3 i_6778975(.A(n_60860), .B(in128[75]), .C(n_60372), .Z(n_79954484
		));
	notech_ao3 i_7178971(.A(n_60860), .B(in128[19]), .C(n_60372), .Z(n_79554480
		));
	notech_ao3 i_7378969(.A(n_60860), .B(in128[66]), .C(n_60372), .Z(n_79354478
		));
	notech_ao3 i_7478968(.A(n_60865), .B(in128[67]), .C(n_60372), .Z(n_79254477
		));
	notech_ao3 i_7578967(.A(n_60865), .B(in128[24]), .C(n_60372), .Z(n_79154476
		));
	notech_ao3 i_7978963(.A(n_60865), .B(in128[87]), .C(n_60376), .Z(n_78754472
		));
	notech_ao3 i_8078962(.A(n_60865), .B(in128[85]), .C(n_60380), .Z(n_78654471
		));
	notech_ao3 i_8278960(.A(n_60865), .B(in128[58]), .C(n_60380), .Z(n_78454469
		));
	notech_ao3 i_8378959(.A(n_60865), .B(in128[52]), .C(n_60380), .Z(n_78354468
		));
	notech_ao3 i_8678956(.A(n_60860), .B(in128[72]), .C(n_60380), .Z(n_78054465
		));
	notech_ao3 i_8978953(.A(n_60860), .B(in128[71]), .C(n_60380), .Z(n_77754462
		));
	notech_ao3 i_9178951(.A(n_60860), .B(in128[18]), .C(n_60380), .Z(n_77554460
		));
	notech_ao3 i_9278950(.A(n_60860), .B(in128[26]), .C(n_60380), .Z(n_77454459
		));
	notech_ao3 i_9478949(.A(n_60860), .B(in128[47]), .C(n_60380), .Z(n_77354458
		));
	notech_ao3 i_9578948(.A(n_60860), .B(in128[64]), .C(n_60380), .Z(n_77254457
		));
	notech_ao3 i_9678947(.A(n_60860), .B(in128[55]), .C(n_60380), .Z(n_77154456
		));
	notech_ao3 i_9978944(.A(n_60860), .B(in128[20]), .C(n_60380), .Z(n_76854453
		));
	notech_ao3 i_10078943(.A(n_60860), .B(in128[78]), .C(n_60376), .Z(n_76754452
		));
	notech_ao3 i_10278941(.A(n_60860), .B(in128[39]), .C(n_60376), .Z(n_76554450
		));
	notech_ao3 i_10378940(.A(n_60860), .B(in128[44]), .C(n_60376), .Z(n_76454449
		));
	notech_ao3 i_10478939(.A(n_60860), .B(in128[31]), .C(n_60376), .Z(n_76354448
		));
	notech_ao3 i_10578938(.A(n_60860), .B(in128[56]), .C(n_60376), .Z(n_76254447
		));
	notech_ao3 i_10678937(.A(n_60865), .B(in128[59]), .C(n_60376), .Z(n_76154446
		));
	notech_ao3 i_10778936(.A(n_60870), .B(in128[60]), .C(n_60380), .Z(n_76054445
		));
	notech_ao3 i_10878935(.A(n_60870), .B(in128[63]), .C(n_60380), .Z(n_75954444
		));
	notech_ao3 i_10978934(.A(n_60870), .B(in128[35]), .C(n_60380), .Z(n_75854443
		));
	notech_ao3 i_11078933(.A(n_60870), .B(in128[51]), .C(n_60376), .Z(n_75754442
		));
	notech_ao3 i_11178932(.A(n_60870), .B(in128[42]), .C(n_60376), .Z(n_75654441
		));
	notech_ao3 i_11278931(.A(n_60870), .B(in128[76]), .C(n_60371), .Z(n_75554440
		));
	notech_ao3 i_11378930(.A(n_60871), .B(in128[50]), .C(n_60362), .Z(n_75454439
		));
	notech_ao3 i_11478929(.A(n_60871), .B(in128[36]), .C(n_60362), .Z(n_75354438
		));
	notech_ao3 i_11578928(.A(n_60871), .B(in128[43]), .C(n_60362), .Z(n_75254437
		));
	notech_ao3 i_11678927(.A(n_60870), .B(in128[74]), .C(n_60362), .Z(n_75154436
		));
	notech_ao3 i_11878925(.A(n_60870), .B(in128[32]), .C(n_60362), .Z(n_74954434
		));
	notech_ao3 i_11978924(.A(n_60870), .B(in128[34]), .C(n_60362), .Z(n_74854433
		));
	notech_ao3 i_12278921(.A(n_60870), .B(in128[48]), .C(n_60362), .Z(n_74554430
		));
	notech_ao3 i_12378920(.A(n_60865), .B(in128[40]), .C(n_60367), .Z(n_74454429
		));
	notech_ao3 i_12478919(.A(n_60870), .B(in128[68]), .C(n_60362), .Z(n_74354428
		));
	notech_ao3 i_12678917(.A(n_60870), .B(in128[28]), .C(n_60362), .Z(n_74154426
		));
	notech_ao3 i_12878915(.A(n_60865), .B(\to_acu2_0[19] ), .C(n_60362), .Z(n_73954424
		));
	notech_ao3 i_13078913(.A(n_60865), .B(\to_acu2_0[24] ), .C(n_60361), .Z(n_73754422
		));
	notech_ao3 i_13178912(.A(n_60865), .B(\to_acu2_0[25] ), .C(n_60361), .Z(n_73654421
		));
	notech_ao3 i_13278911(.A(n_60870), .B(\to_acu2_0[27] ), .C(n_60361), .Z(n_73554420
		));
	notech_ao3 i_13378910(.A(n_60870), .B(\to_acu2_0[28] ), .C(n_60361), .Z(n_73454419
		));
	notech_ao3 i_14678897(.A(n_60870), .B(\to_acu2_0[21] ), .C(n_60361), .Z(n_72154406
		));
	notech_ao3 i_14778896(.A(n_60870), .B(\to_acu2_0[22] ), .C(n_60361), .Z(n_72054405
		));
	notech_ao3 i_14878895(.A(n_60870), .B(\to_acu2_0[23] ), .C(n_60362), .Z(n_71954404
		));
	notech_ao3 i_17778867(.A(n_60870), .B(in128[110]), .C(n_60362), .Z(n_69154376
		));
	notech_ao3 i_18178863(.A(n_60859), .B(in128[106]), .C(n_60362), .Z(n_68754372
		));
	notech_ao3 i_18278862(.A(n_60848), .B(in128[105]), .C(n_60361), .Z(n_68654371
		));
	notech_ao3 i_18378861(.A(n_60848), .B(in128[104]), .C(n_60362), .Z(n_68554370
		));
	notech_ao3 i_18478860(.A(n_60848), .B(in128[103]), .C(n_60367), .Z(n_68454369
		));
	notech_ao3 i_18578859(.A(n_60848), .B(in128[102]), .C(n_60371), .Z(n_68354368
		));
	notech_ao3 i_18678858(.A(n_60848), .B(in128[101]), .C(n_60371), .Z(n_68254367
		));
	notech_ao3 i_18778857(.A(n_60848), .B(in128[100]), .C(n_60371), .Z(n_68154366
		));
	notech_ao3 i_18878856(.A(n_60854), .B(in128[94]), .C(n_60367), .Z(n_68054365
		));
	notech_ao3 i_18978855(.A(n_60854), .B(in128[92]), .C(n_60371), .Z(n_67954364
		));
	notech_ao3 i_19078854(.A(n_60854), .B(in128[91]), .C(n_60371), .Z(n_67854363
		));
	notech_ao3 i_19178853(.A(n_60848), .B(in128[90]), .C(n_60371), .Z(n_67654362
		));
	notech_ao3 i_19278852(.A(n_60848), .B(in128[89]), .C(n_60371), .Z(n_67554361
		));
	notech_ao3 i_19378851(.A(n_60848), .B(in128[88]), .C(n_60371), .Z(n_67454360
		));
	notech_ao3 i_21578832(.A(n_60848), .B(\to_acu2_0[41] ), .C(n_60371), .Z(n_65554341
		));
	notech_ao3 i_21778831(.A(n_60847), .B(in128[57]), .C(n_60371), .Z(n_65454340
		));
	notech_ao3 i_21878830(.A(n_60847), .B(in128[45]), .C(n_60367), .Z(n_65354339
		));
	notech_ao3 i_21978829(.A(n_60847), .B(in128[69]), .C(n_60367), .Z(n_65254338
		));
	notech_ao3 i_22178828(.A(n_60847), .B(in128[53]), .C(n_60367), .Z(n_65154337
		));
	notech_ao3 i_22378826(.A(n_60847), .B(in128[49]), .C(n_60367), .Z(n_64954335
		));
	notech_ao3 i_22478825(.A(n_60847), .B(in128[73]), .C(n_60367), .Z(n_64854334
		));
	notech_and2 i_458(.A(n_3073), .B(n_2427), .Z(n_3074));
	notech_ao4 i_457(.A(n_3072), .B(n_44572), .C(n_44563), .D(n_3069), .Z(n_3073
		));
	notech_or4 i_36(.A(n_3057), .B(n_3062), .C(n_3060), .D(n_2423), .Z(n_3072
		));
	notech_or2 i_35(.A(n_3060), .B(n_3068), .Z(n_3069));
	notech_nand3 i_450(.A(n_3062), .B(n_3057), .C(n_44161), .Z(n_3068));
	notech_nand2 i_34(.A(n_3057), .B(n_44162), .Z(n_3065));
	notech_or4 i_19(.A(n_2418), .B(n_2417), .C(n_3062), .D(n_2423), .Z(n_3064
		));
	notech_xor2 i_2230105(.A(displc[1]), .B(n_3058), .Z(n_3062));
	notech_or2 i_442(.A(imm_sz[1]), .B(imm_sz[2]), .Z(n_3061));
	notech_nor2 i_2330106(.A(n_2418), .B(n_2417), .Z(n_3060));
	notech_nand2 i_435(.A(displc[1]), .B(n_44163), .Z(n_3059));
	notech_ao4 i_2732(.A(n_2416), .B(n_44370), .C(n_44731), .D(n_44730), .Z(n_3058
		));
	notech_or2 i_2130104(.A(n_2420), .B(n_2419), .Z(n_3057));
	notech_xor2 i_121(.A(n_44731), .B(sib_dec), .Z(n_3056));
	notech_and3 i_316(.A(\fpu_indrm[7] ), .B(\fpu_modrm[2] ), .C(\fpu_indrm[0] 
		), .Z(n_3052));
	notech_and4 i_308(.A(n_44718), .B(n_44757), .C(n_44755), .D(n_44756), .Z
		(n_3046));
	notech_and4 i_299(.A(n_44718), .B(n_44754), .C(n_44753), .D(n_44716), .Z
		(n_3041));
	notech_ao3 i_271(.A(ie), .B(n_44744), .C(ipg_fault), .Z(n_3037));
	notech_nand2 i_265(.A(n_43405), .B(n_43403), .Z(n_3033));
	notech_or4 i_267(.A(ififo_rvect1[5]), .B(ififo_rvect1[4]), .C(ififo_rvect1
		[7]), .D(ififo_rvect1[6]), .Z(n_3032));
	notech_or2 i_2235(.A(int_excl[5]), .B(n_1730), .Z(n_3029));
	notech_nand2 i_260(.A(n_62016), .B(term_f), .Z(n_3028));
	notech_nand3 i_257(.A(n_2395), .B(n_43434), .C(n_43431), .Z(n_3027));
	notech_nand2 i_6274(.A(n_43434), .B(n_43431), .Z(n_3026));
	notech_or2 i_327(.A(n_2975), .B(pc_req), .Z(n_3025));
	notech_and4 i_247(.A(n_60937), .B(n_2385), .C(n_44164), .D(n_2384), .Z(n_3022
		));
	notech_nand3 i_76(.A(n_1676), .B(n_44167), .C(n_44165), .Z(n_3020));
	notech_nao3 i_65839(.A(fsm[0]), .B(n_43437), .C(n_2970), .Z(n_3017));
	notech_nand2 i_22(.A(n_3014), .B(n_44729), .Z(n_3015));
	notech_and3 i_17(.A(n_1676), .B(n_44167), .C(n_44165), .Z(n_3014));
	notech_ao3 i_6243(.A(n_44729), .B(\to_acu2_0[62] ), .C(twobyte), .Z(n_3012
		));
	notech_ao3 i_20(.A(n_44729), .B(\to_acu2_0[69] ), .C(twobyte), .Z(n_3009
		));
	notech_or4 i_1130086(.A(in128[8]), .B(in128[14]), .C(n_44723), .D(n_3004
		), .Z(n_3007));
	notech_nand2 i_180(.A(n_44719), .B(n_59489), .Z(n_3004));
	notech_ao3 i_25(.A(n_2336), .B(n_42549), .C(ipg_fault), .Z(n_2999));
	notech_nor2 i_24(.A(ipg_fault), .B(n_2997), .Z(n_2998));
	notech_and2 i_6228(.A(n_62016), .B(n_42622), .Z(n_2997));
	notech_ao3 i_3779(.A(n_60848), .B(n_44744), .C(n_2994), .Z(n_2996));
	notech_and2 i_5(.A(n_60848), .B(n_44744), .Z(n_2995));
	notech_or4 i_65845(.A(fsm[2]), .B(fsm[1]), .C(fsm[0]), .D(n_2969), .Z(n_2994
		));
	notech_ao4 i_160(.A(n_2989), .B(n_44186), .C(valid_len[4]), .D(n_2980), 
		.Z(n_2990));
	notech_or2 i_14(.A(valid_len[2]), .B(valid_len[3]), .Z(n_2989));
	notech_xor2 i_6239(.A(n_2977), .B(n_2984), .Z(n_2985));
	notech_xor2 i_119(.A(imm_sz[1]), .B(i_ptr[1]), .Z(n_2984));
	notech_xor2 i_6238(.A(n_2978), .B(n_2982), .Z(n_2983));
	notech_xor2 i_29(.A(imm_sz[2]), .B(i_ptr[2]), .Z(n_2982));
	notech_xor2 i_6237(.A(i_ptr[3]), .B(n_2979), .Z(n_2981));
	notech_nand2 i_6235(.A(i_ptr[3]), .B(n_44187), .Z(n_2980));
	notech_ao4 i_6236(.A(n_2362), .B(n_44188), .C(n_44372), .D(n_43428), .Z(n_2979
		));
	notech_ao4 i_2130186(.A(n_2977), .B(n_2352), .C(imm_sz[1]), .D(i_ptr[1])
		, .Z(n_2978));
	notech_and2 i_6234(.A(i_ptr[0]), .B(imm_sz[0]), .Z(n_2977));
	notech_nand2 i_187(.A(fsm[0]), .B(fsm[1]), .Z(n_2976));
	notech_or4 i_6246(.A(fsm[3]), .B(fsm[0]), .C(fsm[1]), .D(n_2972), .Z(n_2975
		));
	notech_nand2 i_185(.A(fsm[2]), .B(n_43441), .Z(n_2972));
	notech_or2 i_72(.A(fsm[2]), .B(n_2969), .Z(n_2970));
	notech_or2 i_165(.A(fsm[4]), .B(fsm[3]), .Z(n_2969));
	notech_and4 i_47(.A(n_2338), .B(n_44732), .C(n_44691), .D(n_44690), .Z(n_2967
		));
	notech_and4 i_45(.A(n_44689), .B(n_44688), .C(n_44687), .D(n_44686), .Z(n_2964
		));
	notech_ao4 i_116(.A(n_42553), .B(n_2347), .C(n_2345), .D(n_44745), .Z(n_2960
		));
	notech_and4 i_54(.A(n_2954), .B(n_2951), .C(n_2948), .D(n_44745), .Z(n_2957
		));
	notech_nand3 i_65693(.A(n_2954), .B(n_2951), .C(n_2948), .Z(n_2956));
	notech_and4 i_95(.A(n_44705), .B(n_44704), .C(n_44750), .D(n_44703), .Z(n_2954
		));
	notech_and4 i_93(.A(n_44702), .B(n_44701), .C(n_44700), .D(n_44749), .Z(n_2951
		));
	notech_and4 i_97(.A(n_44695), .B(n_44694), .C(n_2340), .D(n_2947), .Z(n_2948
		));
	notech_and4 i_79(.A(n_44699), .B(n_44698), .C(n_44697), .D(n_44696), .Z(n_2947
		));
	notech_and3 i_61(.A(n_3014), .B(n_2379), .C(n_44729), .Z(n_2942));
	notech_ao4 i_123139(.A(n_59229), .B(n_43459), .C(n_44737), .D(n_43596), 
		.Z(n_2941));
	notech_ao4 i_223140(.A(n_59229), .B(n_43461), .C(n_60243), .D(n_43445), 
		.Z(n_2939));
	notech_ao4 i_323141(.A(n_59229), .B(n_43464), .C(n_43446), .D(n_43032), 
		.Z(n_2937));
	notech_ao4 i_123136(.A(n_59218), .B(n_44197), .C(n_60243), .D(n_44523), 
		.Z(n_2935));
	notech_ao4 i_223137(.A(n_59206), .B(n_44198), .C(n_60241), .D(n_44524), 
		.Z(n_2933));
	notech_nand3 i_323138(.A(n_2891), .B(n_60848), .C(n_2930), .Z(n_2931));
	notech_nand3 i_1288(.A(n_60921), .B(opz1[2]), .C(n_60848), .Z(n_2930));
	notech_ao4 i_126317(.A(n_59206), .B(n_43826), .C(n_60241), .D(n_44758), 
		.Z(n_2929));
	notech_ao4 i_226318(.A(n_59206), .B(n_43829), .C(n_60241), .D(n_44735), 
		.Z(n_2927));
	notech_ao4 i_326319(.A(n_59206), .B(n_43830), .C(n_60241), .D(n_44748), 
		.Z(n_2925));
	notech_ao4 i_426320(.A(n_59206), .B(n_43831), .C(n_60241), .D(n_44747), 
		.Z(n_2923));
	notech_ao4 i_526321(.A(n_59206), .B(n_43833), .C(n_60238), .D(n_44751), 
		.Z(n_2921));
	notech_ao4 i_626322(.A(n_59206), .B(n_43835), .C(n_60236), .D(n_44734), 
		.Z(n_2919));
	notech_ao4 i_726323(.A(n_59206), .B(n_43836), .C(n_60236), .D(n_44733), 
		.Z(n_2917));
	notech_ao4 i_5526371(.A(n_59206), .B(n_43929), .C(n_60236), .D(n_44732),
		 .Z(n_2915));
	notech_or2 i_299098324(.A(n_43465), .B(pfx_sz[0]), .Z(n_1621100926));
	notech_and2 i_294598325(.A(lenpc1[19]), .B(n_59405), .Z(n_1622100927));
	notech_nand3 i_1825656(.A(n_60937), .B(n_2912), .C(n_2910), .Z(n_2913)
		);
	notech_ao3 i_299298327(.A(n_60848), .B(n_1589100894), .C(n_2994), .Z(n_1623100928
		));
	notech_ao3 i_299398328(.A(n_60848), .B(n_1586100891), .C(n_2994), .Z(n_1624100929
		));
	notech_ao3 i_299598329(.A(n_1583100888), .B(n_60854), .C(n_2994), .Z(n_1625100930
		));
	notech_ao3 i_3216(.A(n_60859), .B(in128[0]), .C(n_2994), .Z(n_1626100931
		));
	notech_ao3 i_3289(.A(n_1676), .B(n_60859), .C(n_2994), .Z(n_1627100932)
		);
	notech_ao3 i_3290(.A(n_3029), .B(start), .C(int_excl[0]), .Z(n_1628100933
		));
	notech_ao3 i_3291(.A(n_3029), .B(start), .C(n_1566100871), .Z(n_1629100934
		));
	notech_ao3 i_3292(.A(n_3029), .B(n_1563100868), .C(n_1915), .Z(n_1630100935
		));
	notech_ao3 i_3293(.A(int_excl[5]), .B(n_1730), .C(n_1915), .Z(n_1631100936
		));
	notech_or4 i_3311(.A(n_2975), .B(n_42549), .C(n_42611), .D(pc_req), .Z(n_1632100937
		));
	notech_ao3 i_3666(.A(n_60859), .B(n_44729), .C(n_2994), .Z(n_1633100938)
		);
	notech_or4 i_3682(.A(n_3256), .B(n_1733), .C(\to_acu2_0[4] ), .D(n_1892)
		, .Z(n_1634100939));
	notech_ao3 i_3694(.A(n_60859), .B(in128[16]), .C(n_57724), .Z(n_1635100940
		));
	notech_ao3 i_3695(.A(n_60859), .B(in128[17]), .C(n_57724), .Z(n_1636100941
		));
	notech_ao3 i_3696(.A(n_60859), .B(in128[18]), .C(n_57724), .Z(n_1637100942
		));
	notech_ao3 i_3697(.A(n_60859), .B(\to_acu2_0[0] ), .C(n_57724), .Z(n_1638100943
		));
	notech_ao3 i_3700(.A(n_60859), .B(\to_acu2_0[2] ), .C(n_57724), .Z(n_1639100944
		));
	notech_ao3 i_3701(.A(n_60859), .B(\to_acu2_0[3] ), .C(n_57724), .Z(n_1640100945
		));
	notech_ao3 i_3702(.A(n_60859), .B(\to_acu2_0[4] ), .C(n_57724), .Z(n_1641100946
		));
	notech_ao3 i_3703(.A(n_60859), .B(\to_acu2_0[7] ), .C(n_2994), .Z(n_1642100947
		));
	notech_ao3 i_3704(.A(opz[2]), .B(n_60859), .C(n_57724), .Z(n_1643100948)
		);
	notech_nand3 i_1269(.A(inst_deco1[17]), .B(n_59405), .C(n_2995), .Z(n_2912
		));
	notech_nand2 i_10(.A(n_44744), .B(pc_req), .Z(n_2911));
	notech_or4 i_1268(.A(n_60367), .B(pc_req), .C(pg_fault), .D(n_44395), .Z
		(n_2910));
	notech_nand3 i_2225660(.A(n_60937), .B(n_2908), .C(n_2907), .Z(n_2909)
		);
	notech_reg term_f_reg(.CP(n_63217), .D(n_62016), .CD(n_62619), .Q(term_f
		));
	notech_reg twobyte_reg(.CP(n_63217), .D(n_34252), .CD(n_62619), .Q(twobyte
		));
	notech_mux2 i_36022(.S(n_3292), .A(n_41609), .B(twobyte), .Z(n_34252));
	notech_nand3 i_1263(.A(n_2995), .B(inst_deco1[21]), .C(n_59405), .Z(n_2908
		));
	notech_reg opz_reg_0(.CP(n_63217), .D(n_34261), .CD(n_62619), .Q(opz[0])
		);
	notech_and2 i_36032(.A(n_5765), .B(opz[0]), .Z(n_34261));
	notech_or4 i_1262(.A(n_60367), .B(pc_req), .C(pg_fault), .D(n_44400), .Z
		(n_2907));
	notech_reg opz_reg_1(.CP(n_63217), .D(n_34264), .CD(n_62619), .Q(opz[1])
		);
	notech_mux2 i_36038(.S(\nbus_13545[1] ), .A(opz[1]), .B(n_1643100948), .Z
		(n_34264));
	notech_nand3 i_323135(.A(n_2891), .B(n_60859), .C(n_2905), .Z(n_2906));
	notech_reg_set opz_reg_2(.CP(n_63217), .D(n_34270), .SD(n_62619), .Q(opz
		[2]));
	notech_mux2 i_36046(.S(\nbus_13545[1] ), .A(opz[2]), .B(n_42683), .Z(n_34270
		));
	notech_nand3 i_1260(.A(n_60921), .B(opz2[2]), .C(n_60854), .Z(n_2905));
	notech_reg db67_reg(.CP(n_63217), .D(n_34276), .CD(n_62619), .Q(db67));
	notech_mux2 i_36054(.S(n_46115), .A(db67), .B(n_46118), .Z(n_34276));
	notech_ao4 i_122105(.A(n_59206), .B(n_44150), .C(n_60238), .D(n_44739), 
		.Z(n_2904));
	notech_reg_set fpu_indrm_reg_0(.CP(n_63217), .D(n_34282), .SD(1'b1), .Q(\fpu_indrm[0] 
		));
	notech_mux2 i_36062(.S(n_3293), .A(n_1638100943), .B(\fpu_indrm[0] ), .Z
		(n_34282));
	notech_reg_set fpu_indrm_reg_2(.CP(n_63217), .D(n_34288), .SD(1'b1), .Q(\fpu_indrm[2] 
		));
	notech_mux2 i_36070(.S(n_3293), .A(n_1639100944), .B(\fpu_indrm[2] ), .Z
		(n_34288));
	notech_ao4 i_3927826(.A(n_59208), .B(n_42817), .C(n_55701), .D(n_43832),
		 .Z(n_2902));
	notech_reg_set fpu_indrm_reg_3(.CP(n_63217), .D(n_34294), .SD(1'b1), .Q(\fpu_indrm[3] 
		));
	notech_mux2 i_36078(.S(n_3293), .A(n_1640100945), .B(\fpu_indrm[3] ), .Z
		(n_34294));
	notech_reg_set fpu_indrm_reg_4(.CP(n_63217), .D(n_34300), .SD(1'b1), .Q(\fpu_indrm[4] 
		));
	notech_mux2 i_36086(.S(n_3293), .A(n_1641100946), .B(\fpu_indrm[4] ), .Z
		(n_34300));
	notech_ao4 i_627211(.A(n_59208), .B(n_43471), .C(n_60236), .D(n_43466), 
		.Z(n_2900));
	notech_reg_set fpu_indrm_reg_7(.CP(n_63217), .D(n_34306), .SD(1'b1), .Q(\fpu_indrm[7] 
		));
	notech_mux2 i_36094(.S(n_3293), .A(n_1642100947), .B(\fpu_indrm[7] ), .Z
		(n_34306));
	notech_reg_set fpu_modrm_reg_0(.CP(n_63215), .D(n_34312), .SD(1'b1), .Q(\fpu_modrm[0] 
		));
	notech_mux2 i_36102(.S(n_3293), .A(n_1635100940), .B(\fpu_modrm[0] ), .Z
		(n_34312));
	notech_ao4 i_17726282(.A(n_60236), .B(n_44617), .C(n_59208), .D(n_43779)
		, .Z(n_2898));
	notech_reg_set fpu_modrm_reg_1(.CP(n_63215), .D(n_34318), .SD(1'b1), .Q(\fpu_modrm[1] 
		));
	notech_mux2 i_36110(.S(n_3293), .A(n_1636100941), .B(\fpu_modrm[1] ), .Z
		(n_34318));
	notech_reg_set fpu_modrm_reg_2(.CP(n_63215), .D(n_34324), .SD(1'b1), .Q(\fpu_modrm[2] 
		));
	notech_mux2 i_36118(.S(n_3293), .A(n_1637100942), .B(\fpu_modrm[2] ), .Z
		(n_34324));
	notech_ao4 i_627205(.A(n_59208), .B(n_43469), .C(n_60236), .D(n_43466), 
		.Z(n_2896));
	notech_reg displc_reg_0(.CP(n_63215), .D(n_34330), .CD(n_62619), .Q(displc
		[0]));
	notech_mux2 i_36126(.S(n_3294), .A(n_2704), .B(displc[0]), .Z(n_34330)
		);
	notech_reg displc_reg_1(.CP(n_63215), .D(n_34336), .CD(n_62619), .Q(displc
		[1]));
	notech_mux2 i_36134(.S(n_3294), .A(n_42616), .B(displc[1]), .Z(n_34336)
		);
	notech_ao4 i_323132(.A(n_59208), .B(n_43457), .C(n_43446), .D(n_43032), 
		.Z(n_2894));
	notech_reg displc_reg_2(.CP(n_63217), .D(n_34342), .CD(n_62619), .Q(displc
		[2]));
	notech_mux2 i_36142(.S(n_3294), .A(n_1551100856), .B(displc[2]), .Z(n_34342
		));
	notech_reg sib_dec_reg(.CP(n_63217), .D(n_34348), .CD(n_62619), .Q(sib_dec
		));
	notech_mux2 i_36150(.S(n_3295), .A(n_41609), .B(sib_dec), .Z(n_34348));
	notech_nand2 i_108(.A(n_2891), .B(n_60854), .Z(n_2892));
	notech_reg mod_dec_reg(.CP(n_63215), .D(n_34354), .CD(n_62619), .Q(mod_dec
		));
	notech_mux2 i_36158(.S(n_3296), .A(n_1633100938), .B(mod_dec), .Z(n_34354
		));
	notech_nao3 i_1227(.A(opz[2]), .B(n_60854), .C(n_60367), .Z(n_2891));
	notech_reg imm2_reg_0(.CP(n_63215), .D(n_34360), .CD(n_62617), .Q(\imm2[0] 
		));
	notech_mux2 i_36166(.S(n_56516), .A(\imm2[0] ), .B(n_44375), .Z(n_34360)
		);
	notech_ao4 i_123097(.A(n_3289), .B(n_43465), .C(n_42549), .D(n_2882), .Z
		(n_2890));
	notech_reg imm2_reg_1(.CP(n_63215), .D(n_34366), .CD(n_62617), .Q(\imm2[1] 
		));
	notech_mux2 i_36174(.S(n_56516), .A(\imm2[1] ), .B(n_44381), .Z(n_34366)
		);
	notech_reg imm2_reg_2(.CP(n_63220), .D(n_34372), .CD(n_62617), .Q(\imm2[2] 
		));
	notech_mux2 i_36182(.S(n_56516), .A(\imm2[2] ), .B(n_44387), .Z(n_34372)
		);
	notech_ao4 i_223098(.A(n_43465), .B(n_2887), .C(n_42549), .D(n_2882), .Z
		(n_2888));
	notech_reg imm2_reg_3(.CP(n_63220), .D(n_34378), .CD(n_62617), .Q(\imm2[3] 
		));
	notech_mux2 i_36190(.S(n_56510), .A(\imm2[3] ), .B(n_44393), .Z(n_34378)
		);
	notech_nor2 i_1220(.A(ipg_fault), .B(n_2885), .Z(n_2887));
	notech_reg imm2_reg_4(.CP(n_63220), .D(n_34384), .CD(n_62617), .Q(\imm2[4] 
		));
	notech_mux2 i_36198(.S(n_56510), .A(\imm2[4] ), .B(n_44399), .Z(n_34384)
		);
	notech_reg imm2_reg_5(.CP(n_63220), .D(n_34390), .CD(n_62619), .Q(\imm2[5] 
		));
	notech_mux2 i_36206(.S(n_56510), .A(\imm2[5] ), .B(n_44405), .Z(n_34390)
		);
	notech_and3 i_1221(.A(n_2336), .B(n_2998), .C(n_3014), .Z(n_2885));
	notech_reg imm2_reg_6(.CP(n_63220), .D(n_34396), .CD(n_62619), .Q(\imm2[6] 
		));
	notech_mux2 i_36214(.S(n_56516), .A(\imm2[6] ), .B(n_44411), .Z(n_34396)
		);
	notech_reg imm2_reg_7(.CP(n_63220), .D(n_34402), .CD(n_62619), .Q(\imm2[7] 
		));
	notech_mux2 i_36222(.S(n_56516), .A(\imm2[7] ), .B(n_44417), .Z(n_34402)
		);
	notech_reg imm2_reg_8(.CP(n_63220), .D(n_34408), .CD(n_62617), .Q(\imm2[8] 
		));
	notech_mux2 i_36230(.S(n_56516), .A(\imm2[8] ), .B(n_44423), .Z(n_34408)
		);
	notech_and2 i_1218(.A(n_60236), .B(n_3288), .Z(n_2882));
	notech_reg imm2_reg_9(.CP(n_63220), .D(n_34414), .CD(n_62619), .Q(\imm2[9] 
		));
	notech_mux2 i_36238(.S(n_56516), .A(\imm2[9] ), .B(n_3470), .Z(n_34414)
		);
	notech_ao4 i_323099(.A(n_2880), .B(n_2336), .C(n_3025), .D(n_42611), .Z(n_2881
		));
	notech_reg imm2_reg_10(.CP(n_63220), .D(n_34420), .CD(n_62622), .Q(\imm2[10] 
		));
	notech_mux2 i_36246(.S(n_56516), .A(\imm2[10] ), .B(n_44435), .Z(n_34420
		));
	notech_ao4 i_1210(.A(n_43465), .B(n_44168), .C(n_60236), .D(n_2997), .Z(n_2880
		));
	notech_reg imm2_reg_11(.CP(n_63220), .D(n_34426), .CD(n_62622), .Q(\imm2[11] 
		));
	notech_mux2 i_36254(.S(n_56516), .A(\imm2[11] ), .B(n_44441), .Z(n_34426
		));
	notech_reg imm2_reg_12(.CP(n_63220), .D(n_34432), .CD(n_62622), .Q(\imm2[12] 
		));
	notech_mux2 i_36262(.S(n_56516), .A(\imm2[12] ), .B(n_44447), .Z(n_34432
		));
	notech_reg imm2_reg_13(.CP(n_63217), .D(n_34438), .CD(n_62622), .Q(\imm2[13] 
		));
	notech_mux2 i_36270(.S(n_56510), .A(\imm2[13] ), .B(n_3471), .Z(n_34438)
		);
	notech_reg imm2_reg_14(.CP(n_63217), .D(n_34444), .CD(n_62622), .Q(\imm2[14] 
		));
	notech_mux2 i_36278(.S(n_56510), .A(\imm2[14] ), .B(n_3472), .Z(n_34444)
		);
	notech_reg imm2_reg_15(.CP(n_63217), .D(n_34450), .CD(n_62622), .Q(\imm2[15] 
		));
	notech_mux2 i_36286(.S(n_56510), .A(\imm2[15] ), .B(n_44465), .Z(n_34450
		));
	notech_nand3 i_222689(.A(n_1912), .B(n_2874), .C(n_2872), .Z(n_2875));
	notech_reg imm2_reg_16(.CP(n_63217), .D(n_34456), .CD(n_62622), .Q(\imm2[16] 
		));
	notech_mux2 i_36294(.S(n_56510), .A(\imm2[16] ), .B(n_44471), .Z(n_34456
		));
	notech_or4 i_1206(.A(pg_fault), .B(n_2336), .C(pc_req), .D(n_1913), .Z(n_2874
		));
	notech_reg imm2_reg_17(.CP(n_63217), .D(n_34462), .CD(n_62622), .Q(\imm2[17] 
		));
	notech_mux2 i_36302(.S(n_56510), .A(\imm2[17] ), .B(n_44477), .Z(n_34462
		));
	notech_xor2 i_1205(.A(n_43434), .B(idx_deco[0]), .Z(n_2873));
	notech_reg imm2_reg_18(.CP(n_63220), .D(n_34468), .CD(n_62622), .Q(\imm2[18] 
		));
	notech_mux2 i_36310(.S(n_56510), .A(\imm2[18] ), .B(n_44483), .Z(n_34468
		));
	notech_or4 i_1207(.A(n_60367), .B(pc_req), .C(pg_fault), .D(n_2873), .Z(n_2872
		));
	notech_reg imm2_reg_19(.CP(n_63220), .D(n_34474), .CD(n_62622), .Q(\imm2[19] 
		));
	notech_mux2 i_36318(.S(n_56510), .A(\imm2[19] ), .B(n_44489), .Z(n_34474
		));
	notech_and4 i_123214(.A(n_43797), .B(n_3284), .C(n_2870), .D(n_3280), .Z
		(n_2871));
	notech_reg imm2_reg_20(.CP(n_63220), .D(n_34480), .CD(n_62622), .Q(\imm2[20] 
		));
	notech_mux2 i_36326(.S(n_56510), .A(\imm2[20] ), .B(n_44495), .Z(n_34480
		));
	notech_or4 i_1179(.A(\to_acu2_0[3] ), .B(\to_acu2_0[2] ), .C(n_44751), .D
		(n_43814), .Z(n_2870));
	notech_reg imm2_reg_21(.CP(n_63217), .D(n_34486), .CD(n_62619), .Q(\imm2[21] 
		));
	notech_mux2 i_36334(.S(n_56510), .A(\imm2[21] ), .B(n_3473), .Z(n_34486)
		);
	notech_reg imm2_reg_22(.CP(n_63217), .D(n_34492), .CD(n_62619), .Q(\imm2[22] 
		));
	notech_mux2 i_36342(.S(n_56510), .A(\imm2[22] ), .B(n_44507), .Z(n_34492
		));
	notech_reg imm2_reg_23(.CP(n_63215), .D(n_34498), .CD(n_62619), .Q(\imm2[23] 
		));
	notech_mux2 i_36350(.S(n_56510), .A(\imm2[23] ), .B(n_44513), .Z(n_34498
		));
	notech_nao3 i_39(.A(n_44747), .B(n_44748), .C(n_2413), .Z(n_2867));
	notech_reg imm2_reg_24(.CP(n_63210), .D(n_34504), .CD(n_62619), .Q(\imm2[24] 
		));
	notech_mux2 i_36358(.S(n_56510), .A(\imm2[24] ), .B(n_44519), .Z(n_34504
		));
	notech_ao4 i_1173(.A(n_3283), .B(n_5721), .C(n_1733), .D(n_3256), .Z(n_2866
		));
	notech_reg imm2_reg_25(.CP(n_63210), .D(n_34510), .CD(n_62619), .Q(\imm2[25] 
		));
	notech_mux2 i_36366(.S(n_56510), .A(\imm2[25] ), .B(n_3474), .Z(n_34510)
		);
	notech_and4 i_1171(.A(n_1676), .B(n_44167), .C(n_44165), .D(n_2862), .Z(n_2865
		));
	notech_reg imm2_reg_26(.CP(n_63210), .D(n_34516), .CD(n_62622), .Q(\imm2[26] 
		));
	notech_mux2 i_36374(.S(n_56516), .A(\imm2[26] ), .B(n_44531), .Z(n_34516
		));
	notech_reg imm2_reg_27(.CP(n_63210), .D(n_34522), .CD(n_62622), .Q(\imm2[27] 
		));
	notech_mux2 i_36382(.S(n_56521), .A(\imm2[27] ), .B(n_44537), .Z(n_34522
		));
	notech_reg imm2_reg_28(.CP(n_63210), .D(n_34528), .CD(n_62622), .Q(\imm2[28] 
		));
	notech_mux2 i_36390(.S(n_56521), .A(\imm2[28] ), .B(n_44543), .Z(n_34528
		));
	notech_nao3 i_1172(.A(n_3014), .B(n_44729), .C(n_2859), .Z(n_2862));
	notech_reg imm2_reg_29(.CP(n_63210), .D(n_34534), .CD(n_62622), .Q(\imm2[29] 
		));
	notech_mux2 i_36398(.S(n_56521), .A(\imm2[29] ), .B(n_44549), .Z(n_34534
		));
	notech_or4 i_223215(.A(n_2701), .B(n_2860), .C(n_3281), .D(n_3270), .Z(n_2861
		));
	notech_reg imm2_reg_30(.CP(n_63210), .D(n_34540), .CD(n_62622), .Q(\imm2[30] 
		));
	notech_mux2 i_36406(.S(n_56521), .A(\imm2[30] ), .B(n_44555), .Z(n_34540
		));
	notech_ao3 i_1165(.A(n_3007), .B(n_2859), .C(n_3263), .Z(n_2860));
	notech_reg imm2_reg_31(.CP(n_63210), .D(n_34546), .CD(n_62612), .Q(\imm2[31] 
		));
	notech_mux2 i_36414(.S(n_56521), .A(\imm2[31] ), .B(n_44561), .Z(n_34546
		));
	notech_or2 i_428(.A(n_2411), .B(n_2409), .Z(n_2859));
	notech_reg imm2_reg_32(.CP(n_63210), .D(n_34552), .CD(n_62612), .Q(\imm2[32] 
		));
	notech_mux2 i_36422(.S(n_56521), .A(\imm2[32] ), .B(n_44567), .Z(n_34552
		));
	notech_ao4 i_96(.A(n_5721), .B(n_3258), .C(db67), .D(n_43465), .Z(n_2858
		));
	notech_reg imm2_reg_33(.CP(n_63210), .D(n_34558), .CD(n_62612), .Q(\imm2[33] 
		));
	notech_mux2 i_36430(.S(n_56522), .A(\imm2[33] ), .B(n_44573), .Z(n_34558
		));
	notech_reg imm2_reg_34(.CP(n_63208), .D(n_34564), .CD(n_62612), .Q(\imm2[34] 
		));
	notech_mux2 i_36438(.S(n_56522), .A(\imm2[34] ), .B(n_44579), .Z(n_34564
		));
	notech_reg imm2_reg_35(.CP(n_63208), .D(n_34570), .CD(n_62612), .Q(\imm2[35] 
		));
	notech_mux2 i_36446(.S(n_56522), .A(\imm2[35] ), .B(n_44585), .Z(n_34570
		));
	notech_or4 i_323216(.A(n_2851), .B(n_2845), .C(n_2846), .D(n_43820), .Z(n_2855
		));
	notech_reg imm2_reg_36(.CP(n_63208), .D(n_34576), .CD(n_62612), .Q(\imm2[36] 
		));
	notech_mux2 i_36454(.S(n_56522), .A(\imm2[36] ), .B(n_44591), .Z(n_34576
		));
	notech_reg imm2_reg_37(.CP(n_63208), .D(n_34582), .CD(n_62612), .Q(\imm2[37] 
		));
	notech_mux2 i_36462(.S(n_56522), .A(\imm2[37] ), .B(n_44597), .Z(n_34582
		));
	notech_reg imm2_reg_38(.CP(n_63208), .D(n_34588), .CD(n_62612), .Q(\imm2[38] 
		));
	notech_mux2 i_36470(.S(n_56522), .A(\imm2[38] ), .B(n_44603), .Z(n_34588
		));
	notech_reg imm2_reg_39(.CP(n_63208), .D(n_34594), .CD(n_62612), .Q(\imm2[39] 
		));
	notech_mux2 i_36478(.S(n_56522), .A(\imm2[39] ), .B(n_44609), .Z(n_34594
		));
	notech_ao4 i_1151(.A(n_2848), .B(n_44199), .C(n_2411), .D(n_2409), .Z(n_2851
		));
	notech_reg imm2_reg_40(.CP(n_63208), .D(n_34600), .CD(n_62612), .Q(\imm2[40] 
		));
	notech_mux2 i_36486(.S(n_56521), .A(\imm2[40] ), .B(n_44615), .Z(n_34600
		));
	notech_and2 i_113(.A(n_44747), .B(n_44748), .Z(n_2850));
	notech_reg imm2_reg_41(.CP(n_63208), .D(n_34606), .CD(n_62612), .Q(\imm2[41] 
		));
	notech_mux2 i_36494(.S(n_56521), .A(\imm2[41] ), .B(n_44621), .Z(n_34606
		));
	notech_or4 i_1148(.A(n_3256), .B(n_3015), .C(\to_acu2_0[4] ), .D(n_44747
		), .Z(n_2849));
	notech_reg imm2_reg_42(.CP(n_63208), .D(n_34612), .CD(n_62610), .Q(\imm2[42] 
		));
	notech_mux2 i_36502(.S(n_56521), .A(\imm2[42] ), .B(n_44627), .Z(n_34612
		));
	notech_nor2 i_1147(.A(n_3007), .B(n_3263), .Z(n_2848));
	notech_reg imm2_reg_43(.CP(n_63208), .D(n_34618), .CD(n_62610), .Q(\imm2[43] 
		));
	notech_mux2 i_36510(.S(n_56516), .A(\imm2[43] ), .B(n_44633), .Z(n_34618
		));
	notech_nao3 i_71(.A(n_42641), .B(n_42638), .C(n_2412), .Z(n_2847));
	notech_reg imm2_reg_44(.CP(n_63208), .D(n_34624), .CD(n_62610), .Q(\imm2[44] 
		));
	notech_mux2 i_36518(.S(n_56521), .A(\imm2[44] ), .B(n_44639), .Z(n_34624
		));
	notech_and4 i_1141(.A(n_2859), .B(n_5712), .C(n_2867), .D(n_3266), .Z(n_2846
		));
	notech_reg imm2_reg_45(.CP(n_63215), .D(n_34630), .CD(n_62610), .Q(\imm2[45] 
		));
	notech_mux2 i_36526(.S(n_56521), .A(\imm2[45] ), .B(n_44645), .Z(n_34630
		));
	notech_and4 i_1140(.A(db67), .B(n_41609), .C(n_2847), .D(fpu), .Z(n_2845
		));
	notech_reg imm2_reg_46(.CP(n_63215), .D(n_34636), .CD(n_62610), .Q(\imm2[46] 
		));
	notech_mux2 i_36534(.S(n_56521), .A(\imm2[46] ), .B(n_44651), .Z(n_34636
		));
	notech_nao3 i_527180(.A(n_1730), .B(n_2843), .C(n_2695), .Z(n_2844));
	notech_reg imm2_reg_47(.CP(n_63215), .D(n_34642), .CD(n_62612), .Q(\imm2[47] 
		));
	notech_mux2 i_36542(.S(n_56521), .A(\imm2[47] ), .B(n_44657), .Z(n_34642
		));
	notech_nand2 i_1097(.A(n_1754), .B(int_excl[4]), .Z(n_2843));
	notech_reg imm1_reg_0(.CP(n_63215), .D(n_34648), .CD(n_62612), .Q(\imm1[0] 
		));
	notech_mux2 i_36550(.S(n_59372), .A(\imm1[0] ), .B(n_42621), .Z(n_34648)
		);
	notech_ao4 i_8625468(.A(n_59206), .B(n_42999), .C(n_60236), .D(n_44473),
		 .Z(n_2842));
	notech_reg imm1_reg_1(.CP(n_63215), .D(n_34654), .CD(n_62610), .Q(\imm1[1] 
		));
	notech_mux2 i_36558(.S(n_59372), .A(\imm1[1] ), .B(n_42623), .Z(n_34654)
		);
	notech_reg imm1_reg_2(.CP(n_63215), .D(n_34660), .CD(n_62610), .Q(\imm1[2] 
		));
	notech_mux2 i_36566(.S(n_59372), .A(\imm1[2] ), .B(n_42625), .Z(n_34660)
		);
	notech_ao4 i_8725469(.A(n_59206), .B(n_43001), .C(n_60238), .D(n_44474),
		 .Z(n_2840));
	notech_reg imm1_reg_3(.CP(n_63215), .D(n_34666), .CD(n_62610), .Q(\imm1[3] 
		));
	notech_mux2 i_36574(.S(n_59366), .A(\imm1[3] ), .B(n_42626), .Z(n_34666)
		);
	notech_reg imm1_reg_4(.CP(n_63215), .D(n_34672), .CD(n_62617), .Q(\imm1[4] 
		));
	notech_mux2 i_36582(.S(n_59366), .A(\imm1[4] ), .B(n_42627), .Z(n_34672)
		);
	notech_ao4 i_8825470(.A(n_59206), .B(n_43003), .C(n_60238), .D(n_44475),
		 .Z(n_2838));
	notech_reg imm1_reg_5(.CP(n_63215), .D(n_34678), .CD(n_62617), .Q(\imm1[5] 
		));
	notech_mux2 i_36590(.S(n_59366), .A(\imm1[5] ), .B(n_42628), .Z(n_34678)
		);
	notech_reg imm1_reg_6(.CP(n_63215), .D(n_34684), .CD(n_62617), .Q(\imm1[6] 
		));
	notech_mux2 i_36598(.S(n_59372), .A(\imm1[6] ), .B(n_42629), .Z(n_34684)
		);
	notech_ao4 i_8925471(.A(n_59208), .B(n_43004), .C(n_60238), .D(n_44476),
		 .Z(n_2836));
	notech_reg imm1_reg_7(.CP(n_63215), .D(n_34690), .CD(n_62617), .Q(\imm1[7] 
		));
	notech_mux2 i_36606(.S(n_59372), .A(\imm1[7] ), .B(n_42631), .Z(n_34690)
		);
	notech_reg imm1_reg_8(.CP(n_63210), .D(n_34696), .CD(n_62617), .Q(\imm1[8] 
		));
	notech_mux2 i_36614(.S(n_59372), .A(\imm1[8] ), .B(n_42632), .Z(n_34696)
		);
	notech_ao4 i_9025472(.A(n_59208), .B(n_43007), .C(n_60238), .D(n_44478),
		 .Z(n_2834));
	notech_reg imm1_reg_9(.CP(n_63210), .D(n_34702), .CD(n_62617), .Q(\imm1[9] 
		));
	notech_mux2 i_36622(.S(n_59372), .A(\imm1[9] ), .B(n_42633), .Z(n_34702)
		);
	notech_reg imm1_reg_10(.CP(n_63210), .D(n_34708), .CD(n_62617), .Q(\imm1[10] 
		));
	notech_mux2 i_36630(.S(n_59372), .A(\imm1[10] ), .B(n_42634), .Z(n_34708
		));
	notech_ao4 i_9125473(.A(n_59206), .B(n_43008), .C(n_60238), .D(n_44479),
		 .Z(n_2832));
	notech_reg imm1_reg_11(.CP(n_63210), .D(n_34714), .CD(n_62617), .Q(\imm1[11] 
		));
	notech_mux2 i_36638(.S(n_59372), .A(\imm1[11] ), .B(n_42635), .Z(n_34714
		));
	notech_reg imm1_reg_12(.CP(n_63210), .D(n_34720), .CD(n_62617), .Q(\imm1[12] 
		));
	notech_mux2 i_36646(.S(n_59372), .A(\imm1[12] ), .B(n_42637), .Z(n_34720
		));
	notech_ao4 i_9225474(.A(n_59203), .B(n_43010), .C(n_60238), .D(n_44480),
		 .Z(n_2830));
	notech_reg imm1_reg_13(.CP(n_63210), .D(n_34726), .CD(n_62617), .Q(\imm1[13] 
		));
	notech_mux2 i_36654(.S(n_59366), .A(\imm1[13] ), .B(n_42639), .Z(n_34726
		));
	notech_reg imm1_reg_14(.CP(n_63210), .D(n_34732), .CD(n_62617), .Q(\imm1[14] 
		));
	notech_mux2 i_36662(.S(n_59366), .A(\imm1[14] ), .B(n_42640), .Z(n_34732
		));
	notech_ao4 i_9325475(.A(n_59201), .B(n_43011), .C(n_60238), .D(n_44481),
		 .Z(n_2828));
	notech_reg imm1_reg_15(.CP(n_63210), .D(n_34738), .CD(n_62612), .Q(\imm1[15] 
		));
	notech_mux2 i_36670(.S(n_59366), .A(\imm1[15] ), .B(n_42643), .Z(n_34738
		));
	notech_reg imm1_reg_16(.CP(n_63210), .D(n_34744), .CD(n_62612), .Q(\imm1[16] 
		));
	notech_mux2 i_36678(.S(n_59366), .A(\imm1[16] ), .B(n_43519), .Z(n_34744
		));
	notech_ao4 i_9425476(.A(n_59203), .B(n_43014), .C(n_60238), .D(n_44482),
		 .Z(n_2826));
	notech_reg imm1_reg_17(.CP(n_63210), .D(n_34750), .CD(n_62612), .Q(\imm1[17] 
		));
	notech_mux2 i_36686(.S(n_59366), .A(\imm1[17] ), .B(n_42644), .Z(n_34750
		));
	notech_reg imm1_reg_18(.CP(n_63227), .D(n_34756), .CD(n_62612), .Q(\imm1[18] 
		));
	notech_mux2 i_36694(.S(n_59366), .A(\imm1[18] ), .B(n_42646), .Z(n_34756
		));
	notech_ao4 i_9525477(.A(n_59203), .B(n_43015), .C(n_60238), .D(n_44484),
		 .Z(n_2824));
	notech_reg imm1_reg_19(.CP(n_63227), .D(n_34762), .CD(n_62612), .Q(\imm1[19] 
		));
	notech_mux2 i_36702(.S(n_59366), .A(\imm1[19] ), .B(n_42647), .Z(n_34762
		));
	notech_reg imm1_reg_20(.CP(n_63227), .D(n_34768), .CD(n_62617), .Q(\imm1[20] 
		));
	notech_mux2 i_36710(.S(n_59366), .A(\imm1[20] ), .B(n_43521), .Z(n_34768
		));
	notech_ao4 i_9625478(.A(n_59203), .B(n_43017), .C(n_60238), .D(n_44485),
		 .Z(n_2822));
	notech_reg imm1_reg_21(.CP(n_63227), .D(n_34774), .CD(n_62617), .Q(\imm1[21] 
		));
	notech_mux2 i_36718(.S(n_59366), .A(\imm1[21] ), .B(n_42648), .Z(n_34774
		));
	notech_reg imm1_reg_22(.CP(n_63227), .D(n_34780), .CD(n_62617), .Q(\imm1[22] 
		));
	notech_mux2 i_36726(.S(n_59366), .A(\imm1[22] ), .B(n_42649), .Z(n_34780
		));
	notech_ao4 i_10225484(.A(n_59201), .B(n_43028), .C(n_60243), .D(n_44492)
		, .Z(n_2820));
	notech_reg imm1_reg_23(.CP(n_63227), .D(n_34786), .CD(n_62612), .Q(\imm1[23] 
		));
	notech_mux2 i_36734(.S(n_59366), .A(\imm1[23] ), .B(n_42650), .Z(n_34786
		));
	notech_reg imm1_reg_24(.CP(n_63227), .D(n_34792), .CD(n_62612), .Q(\imm1[24] 
		));
	notech_mux2 i_36742(.S(n_59366), .A(\imm1[24] ), .B(n_42651), .Z(n_34792
		));
	notech_ao4 i_10425486(.A(n_59201), .B(n_43033), .C(n_60250), .D(n_44494)
		, .Z(n_2818));
	notech_reg imm1_reg_25(.CP(n_63227), .D(n_34798), .CD(n_62622), .Q(\imm1[25] 
		));
	notech_mux2 i_36750(.S(n_59366), .A(\imm1[25] ), .B(n_42652), .Z(n_34798
		));
	notech_reg imm1_reg_26(.CP(n_63227), .D(n_34804), .CD(n_62629), .Q(\imm1[26] 
		));
	notech_mux2 i_36758(.S(n_59372), .A(\imm1[26] ), .B(n_42787), .Z(n_34804
		));
	notech_ao4 i_10825490(.A(n_59201), .B(n_43040), .C(n_60250), .D(n_44499)
		, .Z(n_2816));
	notech_reg imm1_reg_27(.CP(n_63227), .D(n_34810), .CD(n_62629), .Q(\imm1[27] 
		));
	notech_mux2 i_36766(.S(n_59377), .A(\imm1[27] ), .B(n_42653), .Z(n_34810
		));
	notech_reg imm1_reg_28(.CP(n_63227), .D(n_34816), .CD(n_62629), .Q(\imm1[28] 
		));
	notech_mux2 i_36774(.S(n_59377), .A(\imm1[28] ), .B(n_42654), .Z(n_34816
		));
	notech_ao4 i_11425496(.A(n_59201), .B(n_43051), .C(n_60250), .D(n_44505)
		, .Z(n_2814));
	notech_reg imm1_reg_29(.CP(n_63227), .D(n_34822), .CD(n_62629), .Q(\imm1[29] 
		));
	notech_mux2 i_36782(.S(n_59377), .A(\imm1[29] ), .B(n_42655), .Z(n_34822
		));
	notech_reg imm1_reg_30(.CP(n_63227), .D(n_34828), .CD(n_62629), .Q(\imm1[30] 
		));
	notech_mux2 i_36790(.S(n_59377), .A(\imm1[30] ), .B(n_42656), .Z(n_34828
		));
	notech_ao4 i_11525497(.A(n_59201), .B(n_43052), .C(n_60250), .D(n_44506)
		, .Z(n_2812));
	notech_reg imm1_reg_31(.CP(n_63225), .D(n_34834), .CD(n_62629), .Q(\imm1[31] 
		));
	notech_mux2 i_36798(.S(n_59377), .A(\imm1[31] ), .B(n_43524), .Z(n_34834
		));
	notech_reg imm1_reg_32(.CP(n_63225), .D(n_34840), .CD(n_62629), .Q(\imm1[32] 
		));
	notech_mux2 i_36806(.S(n_59377), .A(\imm1[32] ), .B(n_42657), .Z(n_34840
		));
	notech_ao4 i_11625498(.A(n_59203), .B(n_43055), .C(n_60250), .D(n_44508)
		, .Z(n_2810));
	notech_reg imm1_reg_33(.CP(n_63225), .D(n_34846), .CD(n_62629), .Q(\imm1[33] 
		));
	notech_mux2 i_36814(.S(n_59378), .A(\imm1[33] ), .B(n_42659), .Z(n_34846
		));
	notech_reg imm1_reg_34(.CP(n_63227), .D(n_34852), .CD(n_62629), .Q(\imm1[34] 
		));
	notech_mux2 i_36822(.S(n_59378), .A(\imm1[34] ), .B(n_42660), .Z(n_34852
		));
	notech_ao4 i_11925501(.A(n_59203), .B(n_43059), .C(n_60248), .D(n_44511)
		, .Z(n_2808));
	notech_reg imm1_reg_35(.CP(n_63227), .D(n_34858), .CD(n_62629), .Q(\imm1[35] 
		));
	notech_mux2 i_36830(.S(n_59378), .A(\imm1[35] ), .B(n_42661), .Z(n_34858
		));
	notech_reg imm1_reg_36(.CP(n_63227), .D(n_34864), .CD(n_62629), .Q(\imm1[36] 
		));
	notech_mux2 i_36838(.S(n_59378), .A(\imm1[36] ), .B(n_42662), .Z(n_34864
		));
	notech_ao4 i_12125503(.A(n_59203), .B(n_43063), .C(n_60248), .D(n_44514)
		, .Z(n_2806));
	notech_reg imm1_reg_37(.CP(n_63227), .D(n_34870), .CD(n_62629), .Q(\imm1[37] 
		));
	notech_mux2 i_36846(.S(n_59378), .A(\imm1[37] ), .B(n_42663), .Z(n_34870
		));
	notech_reg imm1_reg_38(.CP(n_63227), .D(n_34876), .CD(n_62629), .Q(\imm1[38] 
		));
	notech_mux2 i_36854(.S(n_59378), .A(\imm1[38] ), .B(n_42665), .Z(n_34876
		));
	notech_ao4 i_12325505(.A(n_59203), .B(n_43067), .C(n_60250), .D(n_44516)
		, .Z(n_2804));
	notech_reg imm1_reg_39(.CP(n_63231), .D(n_34882), .CD(n_62629), .Q(\imm1[39] 
		));
	notech_mux2 i_36862(.S(n_59378), .A(\imm1[39] ), .B(n_42666), .Z(n_34882
		));
	notech_reg imm1_reg_40(.CP(n_63231), .D(n_34888), .CD(n_62627), .Q(\imm1[40] 
		));
	notech_mux2 i_36870(.S(n_59377), .A(\imm1[40] ), .B(n_42667), .Z(n_34888
		));
	notech_ao4 i_12525507(.A(n_59203), .B(n_43070), .C(n_60250), .D(n_44518)
		, .Z(n_2802));
	notech_reg imm1_reg_41(.CP(n_63231), .D(n_34894), .CD(n_62629), .Q(\imm1[41] 
		));
	notech_mux2 i_36878(.S(n_59377), .A(\imm1[41] ), .B(n_42668), .Z(n_34894
		));
	notech_reg imm1_reg_42(.CP(n_63231), .D(n_34900), .CD(n_62629), .Q(\imm1[42] 
		));
	notech_mux2 i_36886(.S(n_59377), .A(\imm1[42] ), .B(n_42669), .Z(n_34900
		));
	notech_ao4 i_12725509(.A(n_59203), .B(n_43074), .C(n_60250), .D(n_44521)
		, .Z(n_2800));
	notech_reg imm1_reg_43(.CP(n_63231), .D(n_34906), .CD(n_62629), .Q(\imm1[43] 
		));
	notech_mux2 i_36894(.S(n_59372), .A(\imm1[43] ), .B(n_42672), .Z(n_34906
		));
	notech_reg imm1_reg_44(.CP(n_63231), .D(n_34912), .CD(n_62629), .Q(\imm1[44] 
		));
	notech_mux2 i_36902(.S(n_59377), .A(\imm1[44] ), .B(n_42674), .Z(n_34912
		));
	notech_ao4 i_12825510(.A(n_59203), .B(n_43076), .C(n_60253), .D(n_44522)
		, .Z(n_2798));
	notech_reg imm1_reg_45(.CP(n_63231), .D(n_34918), .CD(n_62629), .Q(\imm1[45] 
		));
	notech_mux2 i_36910(.S(n_59377), .A(\imm1[45] ), .B(n_42676), .Z(n_34918
		));
	notech_reg imm1_reg_46(.CP(n_63231), .D(n_34924), .CD(n_62629), .Q(\imm1[46] 
		));
	notech_mux2 i_36918(.S(n_59377), .A(\imm1[46] ), .B(n_42678), .Z(n_34924
		));
	notech_ao4 i_127724(.A(n_59203), .B(n_42671), .C(n_2428), .D(n_60250), .Z
		(n_2796));
	notech_reg imm1_reg_47(.CP(n_63231), .D(n_34930), .CD(n_62633), .Q(\imm1[47] 
		));
	notech_mux2 i_36926(.S(n_59377), .A(\imm1[47] ), .B(n_42680), .Z(n_34930
		));
	notech_reg inst_deco2_reg_0(.CP(n_63231), .D(n_34936), .CD(n_62633), .Q(inst_deco2
		[0]));
	notech_mux2 i_36934(.S(n_56521), .A(inst_deco2[0]), .B(n_1542100847), .Z
		(n_34936));
	notech_ao4 i_227725(.A(n_59203), .B(n_42673), .C(n_2436), .D(n_60253), .Z
		(n_2794));
	notech_reg inst_deco2_reg_1(.CP(n_63231), .D(n_34942), .CD(n_62633), .Q(inst_deco2
		[1]));
	notech_mux2 i_36942(.S(n_56521), .A(inst_deco2[1]), .B(n_41886), .Z(n_34942
		));
	notech_reg inst_deco2_reg_2(.CP(n_63231), .D(n_34948), .CD(n_62633), .Q(inst_deco2
		[2]));
	notech_mux2 i_36950(.S(n_56521), .A(inst_deco2[2]), .B(n_41892), .Z(n_34948
		));
	notech_ao4 i_327726(.A(n_59203), .B(n_42675), .C(n_2444), .D(n_60253), .Z
		(n_2792));
	notech_reg inst_deco2_reg_3(.CP(n_63231), .D(n_34954), .CD(n_62633), .Q(inst_deco2
		[3]));
	notech_mux2 i_36958(.S(n_56521), .A(inst_deco2[3]), .B(n_41898), .Z(n_34954
		));
	notech_reg inst_deco2_reg_4(.CP(n_63231), .D(n_34960), .CD(n_62633), .Q(inst_deco2
		[4]));
	notech_mux2 i_36966(.S(n_56521), .A(inst_deco2[4]), .B(n_41904), .Z(n_34960
		));
	notech_ao4 i_427727(.A(n_59215), .B(n_42677), .C(n_2452), .D(n_60253), .Z
		(n_2790));
	notech_reg inst_deco2_reg_5(.CP(n_63227), .D(n_34966), .CD(n_62635), .Q(inst_deco2
		[5]));
	notech_mux2 i_36974(.S(n_56499), .A(inst_deco2[5]), .B(n_1543100848), .Z
		(n_34966));
	notech_reg inst_deco2_reg_6(.CP(n_63227), .D(n_34972), .CD(n_62633), .Q(inst_deco2
		[6]));
	notech_mux2 i_36982(.S(n_56499), .A(inst_deco2[6]), .B(n_41916), .Z(n_34972
		));
	notech_ao4 i_527728(.A(n_59215), .B(n_42679), .C(n_2460), .D(n_60250), .Z
		(n_2788));
	notech_reg inst_deco2_reg_7(.CP(n_63231), .D(n_34978), .CD(n_62633), .Q(inst_deco2
		[7]));
	notech_mux2 i_36990(.S(n_56499), .A(inst_deco2[7]), .B(n_1544100849), .Z
		(n_34978));
	notech_reg inst_deco2_reg_8(.CP(n_63231), .D(n_34984), .CD(n_62633), .Q(inst_deco2
		[8]));
	notech_mux2 i_36998(.S(n_56499), .A(inst_deco2[8]), .B(n_1545100850), .Z
		(n_34984));
	notech_ao4 i_627729(.A(n_59215), .B(n_42681), .C(n_2468), .D(n_60250), .Z
		(n_2786));
	notech_reg inst_deco2_reg_9(.CP(n_63231), .D(n_34990), .CD(n_62633), .Q(inst_deco2
		[9]));
	notech_mux2 i_37006(.S(n_56499), .A(inst_deco2[9]), .B(n_41934), .Z(n_34990
		));
	notech_reg inst_deco2_reg_10(.CP(n_63231), .D(n_34996), .CD(n_62633), .Q
		(inst_deco2[10]));
	notech_mux2 i_37014(.S(n_56499), .A(inst_deco2[10]), .B(n_41940), .Z(n_34996
		));
	notech_ao4 i_727730(.A(n_59215), .B(n_42682), .C(n_2476), .D(n_60250), .Z
		(n_2784));
	notech_reg inst_deco2_reg_11(.CP(n_63231), .D(n_35002), .CD(n_62633), .Q
		(inst_deco2[11]));
	notech_mux2 i_37022(.S(n_56499), .A(inst_deco2[11]), .B(n_41946), .Z(n_35002
		));
	notech_reg inst_deco2_reg_12(.CP(n_63225), .D(n_35008), .CD(n_62633), .Q
		(inst_deco2[12]));
	notech_mux2 i_37030(.S(n_56504), .A(inst_deco2[12]), .B(n_41952), .Z(n_35008
		));
	notech_ao4 i_827731(.A(n_59215), .B(n_42684), .C(n_2484), .D(n_60250), .Z
		(n_2782));
	notech_reg inst_deco2_reg_13(.CP(n_63222), .D(n_35014), .CD(n_62633), .Q
		(inst_deco2[13]));
	notech_mux2 i_37038(.S(n_56504), .A(inst_deco2[13]), .B(n_41958), .Z(n_35014
		));
	notech_reg inst_deco2_reg_14(.CP(n_63222), .D(n_35020), .CD(n_62633), .Q
		(inst_deco2[14]));
	notech_mux2 i_37046(.S(n_56504), .A(inst_deco2[14]), .B(n_41964), .Z(n_35020
		));
	notech_ao4 i_927732(.A(n_59215), .B(n_42685), .C(n_2495), .D(n_60250), .Z
		(n_2780));
	notech_reg inst_deco2_reg_15(.CP(n_63222), .D(n_35026), .CD(n_62633), .Q
		(inst_deco2[15]));
	notech_mux2 i_37054(.S(n_56499), .A(inst_deco2[15]), .B(n_41970), .Z(n_35026
		));
	notech_reg inst_deco2_reg_16(.CP(n_63222), .D(n_35032), .CD(n_62633), .Q
		(inst_deco2[16]));
	notech_mux2 i_37062(.S(n_56504), .A(inst_deco2[16]), .B(n_41976), .Z(n_35032
		));
	notech_ao4 i_1027733(.A(n_225599334), .B(n_60248), .C(n_59215), .D(n_42686
		), .Z(n_2778));
	notech_reg inst_deco2_reg_17(.CP(n_63222), .D(n_35038), .CD(n_62633), .Q
		(inst_deco2[17]));
	notech_mux2 i_37070(.S(n_56504), .A(inst_deco2[17]), .B(n_41982), .Z(n_35038
		));
	notech_reg inst_deco2_reg_18(.CP(n_63222), .D(n_35044), .CD(n_62633), .Q
		(inst_deco2[18]));
	notech_mux2 i_37078(.S(n_56499), .A(inst_deco2[18]), .B(n_41988), .Z(n_35044
		));
	notech_ao4 i_1127734(.A(n_59215), .B(n_42687), .C(n_2503), .D(n_60243), 
		.Z(n_2776));
	notech_reg inst_deco2_reg_19(.CP(n_63222), .D(n_35050), .CD(n_62633), .Q
		(inst_deco2[19]));
	notech_mux2 i_37086(.S(n_56499), .A(inst_deco2[19]), .B(n_41994), .Z(n_35050
		));
	notech_reg inst_deco2_reg_20(.CP(n_63222), .D(n_35056), .CD(n_62624), .Q
		(inst_deco2[20]));
	notech_mux2 i_37094(.S(n_56499), .A(inst_deco2[20]), .B(n_42000), .Z(n_35056
		));
	notech_ao4 i_1227735(.A(n_59215), .B(n_42688), .C(n_2511), .D(n_60243), 
		.Z(n_2774));
	notech_reg inst_deco2_reg_21(.CP(n_63222), .D(n_35062), .CD(n_62624), .Q
		(inst_deco2[21]));
	notech_mux2 i_37102(.S(n_56498), .A(inst_deco2[21]), .B(n_42006), .Z(n_35062
		));
	notech_reg inst_deco2_reg_22(.CP(n_63222), .D(n_35068), .CD(n_62624), .Q
		(inst_deco2[22]));
	notech_mux2 i_37110(.S(n_56498), .A(inst_deco2[22]), .B(n_42012), .Z(n_35068
		));
	notech_ao4 i_1327736(.A(n_59215), .B(n_42689), .C(n_2519), .D(n_60243), 
		.Z(n_2772));
	notech_reg inst_deco2_reg_23(.CP(n_63222), .D(n_35074), .CD(n_62624), .Q
		(inst_deco2[23]));
	notech_mux2 i_37118(.S(n_56498), .A(inst_deco2[23]), .B(n_42018), .Z(n_35074
		));
	notech_reg inst_deco2_reg_24(.CP(n_63220), .D(n_35080), .CD(n_62624), .Q
		(inst_deco2[24]));
	notech_mux2 i_37126(.S(n_56499), .A(inst_deco2[24]), .B(n_42024), .Z(n_35080
		));
	notech_ao4 i_1427737(.A(n_225499333), .B(n_60248), .C(n_59218), .D(n_42690
		), .Z(n_2770));
	notech_reg inst_deco2_reg_25(.CP(n_63220), .D(n_35086), .CD(n_62624), .Q
		(inst_deco2[25]));
	notech_mux2 i_37134(.S(n_56499), .A(inst_deco2[25]), .B(n_42030), .Z(n_35086
		));
	notech_reg inst_deco2_reg_26(.CP(n_63220), .D(n_35092), .CD(n_62624), .Q
		(inst_deco2[26]));
	notech_mux2 i_37142(.S(n_56499), .A(inst_deco2[26]), .B(n_42036), .Z(n_35092
		));
	notech_ao4 i_1527738(.A(n_225399332), .B(n_60243), .C(n_59218), .D(n_42691
		), .Z(n_2768));
	notech_reg inst_deco2_reg_27(.CP(n_63220), .D(n_35098), .CD(n_62624), .Q
		(inst_deco2[27]));
	notech_mux2 i_37150(.S(n_56499), .A(inst_deco2[27]), .B(n_42042), .Z(n_35098
		));
	notech_reg inst_deco2_reg_28(.CP(n_63220), .D(n_35104), .CD(n_62624), .Q
		(inst_deco2[28]));
	notech_mux2 i_37158(.S(n_56499), .A(inst_deco2[28]), .B(n_42048), .Z(n_35104
		));
	notech_ao4 i_1627739(.A(n_59218), .B(n_42692), .C(n_2527), .D(n_60243), 
		.Z(n_2766));
	notech_reg inst_deco2_reg_29(.CP(n_63222), .D(n_35110), .CD(n_62624), .Q
		(inst_deco2[29]));
	notech_mux2 i_37166(.S(n_56499), .A(inst_deco2[29]), .B(n_42054), .Z(n_35110
		));
	notech_reg inst_deco2_reg_30(.CP(n_63222), .D(n_35116), .CD(n_62624), .Q
		(inst_deco2[30]));
	notech_mux2 i_37174(.S(n_56499), .A(inst_deco2[30]), .B(n_42060), .Z(n_35116
		));
	notech_ao4 i_1827741(.A(n_59218), .B(n_42694), .C(n_2545), .D(n_60243), 
		.Z(n_2764));
	notech_reg inst_deco2_reg_31(.CP(n_63222), .D(n_35122), .CD(n_62624), .Q
		(inst_deco2[31]));
	notech_mux2 i_37182(.S(n_56504), .A(inst_deco2[31]), .B(n_42066), .Z(n_35122
		));
	notech_reg inst_deco2_reg_32(.CP(n_63220), .D(n_35128), .CD(n_62624), .Q
		(inst_deco2[32]));
	notech_mux2 i_37190(.S(n_56509), .A(inst_deco2[32]), .B(n_42072), .Z(n_35128
		));
	notech_ao4 i_1927742(.A(n_59218), .B(n_42695), .C(n_2553), .D(n_60243), 
		.Z(n_2762));
	notech_reg inst_deco2_reg_33(.CP(n_63222), .D(n_35134), .CD(n_62622), .Q
		(inst_deco2[33]));
	notech_mux2 i_37198(.S(n_56509), .A(inst_deco2[33]), .B(n_42078), .Z(n_35134
		));
	notech_reg inst_deco2_reg_34(.CP(n_63225), .D(n_35140), .CD(n_62622), .Q
		(inst_deco2[34]));
	notech_mux2 i_37206(.S(n_56509), .A(inst_deco2[34]), .B(n_42084), .Z(n_35140
		));
	notech_ao4 i_2027743(.A(n_59215), .B(n_42696), .C(n_2561), .D(n_60243), 
		.Z(n_2760));
	notech_reg inst_deco2_reg_35(.CP(n_63225), .D(n_35146), .CD(n_62622), .Q
		(inst_deco2[35]));
	notech_mux2 i_37214(.S(n_56509), .A(inst_deco2[35]), .B(n_42090), .Z(n_35146
		));
	notech_reg inst_deco2_reg_36(.CP(n_63225), .D(n_35152), .CD(n_62624), .Q
		(inst_deco2[36]));
	notech_mux2 i_37222(.S(n_56509), .A(inst_deco2[36]), .B(n_42096), .Z(n_35152
		));
	notech_ao4 i_2227745(.A(n_225299331), .B(n_60243), .C(n_59215), .D(n_42698
		), .Z(n_2758));
	notech_reg inst_deco2_reg_37(.CP(n_63225), .D(n_35158), .CD(n_62624), .Q
		(inst_deco2[37]));
	notech_mux2 i_37230(.S(n_56509), .A(inst_deco2[37]), .B(n_42102), .Z(n_35158
		));
	notech_reg inst_deco2_reg_38(.CP(n_63225), .D(n_35164), .CD(n_62624), .Q
		(inst_deco2[38]));
	notech_mux2 i_37238(.S(n_56509), .A(inst_deco2[38]), .B(n_42108), .Z(n_35164
		));
	notech_ao4 i_2327746(.A(n_59215), .B(n_42699), .C(n_2577), .D(n_60248), 
		.Z(n_2756));
	notech_reg inst_deco2_reg_39(.CP(n_63225), .D(n_35170), .CD(n_62624), .Q
		(inst_deco2[39]));
	notech_mux2 i_37246(.S(n_56509), .A(inst_deco2[39]), .B(n_42114), .Z(n_35170
		));
	notech_reg inst_deco2_reg_40(.CP(n_63225), .D(n_35176), .CD(n_62624), .Q
		(inst_deco2[40]));
	notech_mux2 i_37254(.S(n_56510), .A(inst_deco2[40]), .B(n_42120), .Z(n_35176
		));
	notech_ao4 i_2427747(.A(n_59218), .B(n_42700), .C(n_2585), .D(n_60248), 
		.Z(n_2754));
	notech_reg inst_deco2_reg_41(.CP(n_63225), .D(n_35182), .CD(n_62627), .Q
		(inst_deco2[41]));
	notech_mux2 i_37262(.S(n_56510), .A(inst_deco2[41]), .B(n_1546100851), .Z
		(n_35182));
	notech_reg inst_deco2_reg_42(.CP(n_63225), .D(n_35188), .CD(n_62627), .Q
		(inst_deco2[42]));
	notech_mux2 i_37270(.S(n_56509), .A(inst_deco2[42]), .B(n_1547100852), .Z
		(n_35188));
	notech_ao4 i_2527748(.A(n_59215), .B(n_42701), .C(n_2595), .D(n_60248), 
		.Z(n_2752));
	notech_reg inst_deco2_reg_43(.CP(n_63225), .D(n_35194), .CD(n_62627), .Q
		(inst_deco2[43]));
	notech_mux2 i_37278(.S(n_56509), .A(inst_deco2[43]), .B(n_1548100853), .Z
		(n_35194));
	notech_reg inst_deco2_reg_44(.CP(n_63225), .D(n_35200), .CD(n_62627), .Q
		(inst_deco2[44]));
	notech_mux2 i_37286(.S(n_56509), .A(inst_deco2[44]), .B(n_1549100854), .Z
		(n_35200));
	notech_ao4 i_2627749(.A(n_225199330), .B(n_60248), .C(n_59213), .D(n_42702
		), .Z(n_2750));
	notech_reg inst_deco2_reg_45(.CP(n_63222), .D(n_35206), .CD(n_62627), .Q
		(inst_deco2[45]));
	notech_mux2 i_37294(.S(n_56504), .A(inst_deco2[45]), .B(n_1550100855), .Z
		(n_35206));
	notech_reg inst_deco2_reg_46(.CP(n_63222), .D(n_35212), .CD(n_62627), .Q
		(inst_deco2[46]));
	notech_mux2 i_37302(.S(n_56504), .A(inst_deco2[46]), .B(n_42156), .Z(n_35212
		));
	notech_ao4 i_2827751(.A(n_59208), .B(n_42704), .C(n_2611), .D(n_60248), 
		.Z(n_2748));
	notech_reg inst_deco2_reg_47(.CP(n_63222), .D(n_35218), .CD(n_62627), .Q
		(inst_deco2[47]));
	notech_mux2 i_37310(.S(n_56504), .A(inst_deco2[47]), .B(n_42162), .Z(n_35218
		));
	notech_reg inst_deco2_reg_48(.CP(n_63222), .D(n_35224), .CD(n_62627), .Q
		(inst_deco2[48]));
	notech_mux2 i_37318(.S(n_56504), .A(inst_deco2[48]), .B(n_42168), .Z(n_35224
		));
	notech_ao4 i_2927752(.A(n_59208), .B(n_42705), .C(n_2619), .D(n_60248), 
		.Z(n_2746));
	notech_reg inst_deco2_reg_49(.CP(n_63222), .D(n_35230), .CD(n_62627), .Q
		(inst_deco2[49]));
	notech_mux2 i_37326(.S(n_56504), .A(inst_deco2[49]), .B(n_42174), .Z(n_35230
		));
	notech_reg inst_deco2_reg_50(.CP(n_63225), .D(n_35236), .CD(n_62627), .Q
		(inst_deco2[50]));
	notech_mux2 i_37334(.S(n_56504), .A(inst_deco2[50]), .B(n_42180), .Z(n_35236
		));
	notech_ao4 i_3027753(.A(n_59213), .B(n_42706), .C(n_2627), .D(n_60248), 
		.Z(n_2744));
	notech_reg inst_deco2_reg_51(.CP(n_63225), .D(n_35242), .CD(n_62627), .Q
		(inst_deco2[51]));
	notech_mux2 i_37342(.S(n_56509), .A(inst_deco2[51]), .B(n_42186), .Z(n_35242
		));
	notech_reg inst_deco2_reg_52(.CP(n_63225), .D(n_35248), .CD(n_62627), .Q
		(inst_deco2[52]));
	notech_mux2 i_37350(.S(n_56509), .A(inst_deco2[52]), .B(n_42192), .Z(n_35248
		));
	notech_ao4 i_3127754(.A(n_59213), .B(n_42707), .C(n_2635), .D(n_60248), 
		.Z(n_2742));
	notech_reg inst_deco2_reg_53(.CP(n_63225), .D(n_35254), .CD(n_62627), .Q
		(inst_deco2[53]));
	notech_mux2 i_37358(.S(n_56509), .A(inst_deco2[53]), .B(n_42198), .Z(n_35254
		));
	notech_reg inst_deco2_reg_54(.CP(n_63225), .D(n_35260), .CD(n_62627), .Q
		(inst_deco2[54]));
	notech_mux2 i_37366(.S(n_56509), .A(inst_deco2[54]), .B(n_42204), .Z(n_35260
		));
	notech_ao4 i_3327756(.A(n_59213), .B(n_42709), .C(n_55701), .D(n_43905),
		 .Z(n_2740));
	notech_reg inst_deco2_reg_55(.CP(n_63192), .D(n_35266), .CD(n_62624), .Q
		(inst_deco2[55]));
	notech_mux2 i_37374(.S(n_56509), .A(inst_deco2[55]), .B(n_42210), .Z(n_35266
		));
	notech_reg inst_deco2_reg_56(.CP(n_63192), .D(n_35272), .CD(n_62624), .Q
		(inst_deco2[56]));
	notech_mux2 i_37382(.S(n_56509), .A(inst_deco2[56]), .B(n_42216), .Z(n_35272
		));
	notech_ao4 i_3427757(.A(n_59208), .B(n_42710), .C(n_55701), .D(n_43903),
		 .Z(n_2738));
	notech_reg inst_deco2_reg_57(.CP(n_63192), .D(n_35278), .CD(n_62627), .Q
		(inst_deco2[57]));
	notech_mux2 i_37390(.S(n_56509), .A(inst_deco2[57]), .B(n_42222), .Z(n_35278
		));
	notech_reg inst_deco2_reg_58(.CP(n_63192), .D(n_35284), .CD(n_62627), .Q
		(inst_deco2[58]));
	notech_mux2 i_37398(.S(n_56522), .A(inst_deco2[58]), .B(n_42228), .Z(n_35284
		));
	notech_ao4 i_3527758(.A(n_59208), .B(n_42711), .C(n_55701), .D(n_43899),
		 .Z(n_2736));
	notech_reg inst_deco2_reg_59(.CP(n_63192), .D(n_35290), .CD(n_62627), .Q
		(inst_deco2[59]));
	notech_mux2 i_37406(.S(n_56538), .A(inst_deco2[59]), .B(n_42234), .Z(n_35290
		));
	notech_reg inst_deco2_reg_60(.CP(n_63194), .D(n_35296), .CD(n_62627), .Q
		(inst_deco2[60]));
	notech_mux2 i_37414(.S(n_56543), .A(inst_deco2[60]), .B(n_42240), .Z(n_35296
		));
	notech_ao4 i_3627759(.A(n_59208), .B(n_42712), .C(n_55701), .D(n_43897),
		 .Z(n_2734));
	notech_reg inst_deco2_reg_61(.CP(n_63194), .D(n_35302), .CD(n_62627), .Q
		(inst_deco2[61]));
	notech_mux2 i_37422(.S(n_56543), .A(inst_deco2[61]), .B(n_42246), .Z(n_35302
		));
	notech_reg inst_deco2_reg_62(.CP(n_63194), .D(n_35308), .CD(n_62610), .Q
		(inst_deco2[62]));
	notech_mux2 i_37430(.S(n_56538), .A(inst_deco2[62]), .B(n_42252), .Z(n_35308
		));
	notech_ao4 i_3727760(.A(n_59208), .B(n_42713), .C(n_55701), .D(n_43893),
		 .Z(n_2732));
	notech_reg inst_deco2_reg_63(.CP(n_63192), .D(n_35314), .CD(n_62594), .Q
		(inst_deco2[63]));
	notech_mux2 i_37438(.S(n_56538), .A(inst_deco2[63]), .B(n_42258), .Z(n_35314
		));
	notech_reg inst_deco2_reg_64(.CP(n_63192), .D(n_35320), .CD(n_62594), .Q
		(inst_deco2[64]));
	notech_mux2 i_37446(.S(n_56538), .A(inst_deco2[64]), .B(n_42264), .Z(n_35320
		));
	notech_ao4 i_3827761(.A(n_59208), .B(n_42714), .C(n_55701), .D(n_43887),
		 .Z(n_2730));
	notech_reg inst_deco2_reg_65(.CP(n_63192), .D(n_35326), .CD(n_62594), .Q
		(inst_deco2[65]));
	notech_mux2 i_37454(.S(n_56543), .A(inst_deco2[65]), .B(n_42270), .Z(n_35326
		));
	notech_reg inst_deco2_reg_66(.CP(n_63192), .D(n_35332), .CD(n_62594), .Q
		(inst_deco2[66]));
	notech_mux2 i_37462(.S(n_56543), .A(inst_deco2[66]), .B(n_42276), .Z(n_35332
		));
	notech_ao4 i_3927762(.A(n_59213), .B(n_42715), .C(n_55701), .D(n_43832),
		 .Z(n_2728));
	notech_reg inst_deco2_reg_67(.CP(n_63192), .D(n_35338), .CD(n_62594), .Q
		(inst_deco2[67]));
	notech_mux2 i_37470(.S(n_56543), .A(inst_deco2[67]), .B(n_42282), .Z(n_35338
		));
	notech_reg inst_deco2_reg_68(.CP(n_63192), .D(n_35344), .CD(n_62596), .Q
		(inst_deco2[68]));
	notech_mux2 i_37478(.S(n_56543), .A(inst_deco2[68]), .B(n_42288), .Z(n_35344
		));
	notech_ao4 i_4027763(.A(n_59213), .B(n_42716), .C(n_55701), .D(n_43879),
		 .Z(n_2726));
	notech_reg inst_deco2_reg_69(.CP(n_63192), .D(n_35350), .CD(n_62596), .Q
		(inst_deco2[69]));
	notech_mux2 i_37486(.S(n_56543), .A(inst_deco2[69]), .B(n_42294), .Z(n_35350
		));
	notech_reg inst_deco2_reg_70(.CP(n_63192), .D(n_35356), .CD(n_62596), .Q
		(inst_deco2[70]));
	notech_mux2 i_37494(.S(n_56543), .A(inst_deco2[70]), .B(n_42300), .Z(n_35356
		));
	notech_ao4 i_4127764(.A(n_59213), .B(n_42717), .C(n_55762), .D(n_43861),
		 .Z(n_2724));
	notech_reg inst_deco2_reg_71(.CP(n_63192), .D(n_35362), .CD(n_62596), .Q
		(inst_deco2[71]));
	notech_mux2 i_37502(.S(n_56543), .A(inst_deco2[71]), .B(n_42306), .Z(n_35362
		));
	notech_reg inst_deco2_reg_72(.CP(n_63192), .D(n_35368), .CD(n_62596), .Q
		(inst_deco2[72]));
	notech_mux2 i_37510(.S(n_56533), .A(inst_deco2[72]), .B(n_42312), .Z(n_35368
		));
	notech_ao4 i_4227765(.A(n_59213), .B(n_42718), .C(n_55762), .D(n_43857),
		 .Z(n_2722));
	notech_reg inst_deco2_reg_73(.CP(n_63192), .D(n_35374), .CD(n_62594), .Q
		(inst_deco2[73]));
	notech_mux2 i_37518(.S(n_56533), .A(inst_deco2[73]), .B(n_42318), .Z(n_35374
		));
	notech_reg inst_deco2_reg_74(.CP(n_63192), .D(n_35380), .CD(n_62594), .Q
		(inst_deco2[74]));
	notech_mux2 i_37526(.S(n_56538), .A(inst_deco2[74]), .B(n_42324), .Z(n_35380
		));
	notech_ao4 i_4327766(.A(n_59213), .B(n_42719), .C(n_55762), .D(n_43855),
		 .Z(n_2720));
	notech_reg inst_deco2_reg_75(.CP(n_63192), .D(n_35386), .CD(n_62594), .Q
		(inst_deco2[75]));
	notech_mux2 i_37534(.S(n_56533), .A(inst_deco2[75]), .B(n_42330), .Z(n_35386
		));
	notech_reg inst_deco2_reg_76(.CP(n_63194), .D(n_35392), .CD(n_62594), .Q
		(inst_deco2[76]));
	notech_mux2 i_37542(.S(n_56533), .A(inst_deco2[76]), .B(n_42336), .Z(n_35392
		));
	notech_ao4 i_4427767(.A(n_59213), .B(n_42720), .C(n_55762), .D(n_43851),
		 .Z(n_2718));
	notech_reg inst_deco2_reg_77(.CP(n_63194), .D(n_35398), .CD(n_62594), .Q
		(inst_deco2[77]));
	notech_mux2 i_37550(.S(n_56533), .A(inst_deco2[77]), .B(n_42342), .Z(n_35398
		));
	notech_reg inst_deco2_reg_78(.CP(n_63194), .D(n_35404), .CD(n_62594), .Q
		(inst_deco2[78]));
	notech_mux2 i_37558(.S(n_56538), .A(inst_deco2[78]), .B(n_42348), .Z(n_35404
		));
	notech_ao4 i_4527768(.A(n_59213), .B(n_42722), .C(n_55762), .D(n_43849),
		 .Z(n_2716));
	notech_reg inst_deco2_reg_79(.CP(n_63194), .D(n_35410), .CD(n_62594), .Q
		(inst_deco2[79]));
	notech_mux2 i_37566(.S(n_56538), .A(inst_deco2[79]), .B(n_42354), .Z(n_35410
		));
	notech_reg inst_deco2_reg_80(.CP(n_63194), .D(n_35416), .CD(n_62594), .Q
		(inst_deco2[80]));
	notech_mux2 i_37574(.S(n_56538), .A(inst_deco2[80]), .B(n_42360), .Z(n_35416
		));
	notech_ao4 i_4627769(.A(n_59213), .B(n_42723), .C(n_55762), .D(n_43845),
		 .Z(n_2714));
	notech_reg inst_deco2_reg_81(.CP(n_63198), .D(n_35422), .CD(n_62594), .Q
		(inst_deco2[81]));
	notech_mux2 i_37582(.S(n_56538), .A(inst_deco2[81]), .B(n_42366), .Z(n_35422
		));
	notech_reg inst_deco2_reg_82(.CP(n_63198), .D(n_35428), .CD(n_62594), .Q
		(inst_deco2[82]));
	notech_mux2 i_37590(.S(n_56538), .A(inst_deco2[82]), .B(n_42372), .Z(n_35428
		));
	notech_ao4 i_4727770(.A(n_59213), .B(n_42725), .C(n_55762), .D(n_43841),
		 .Z(n_2712));
	notech_reg inst_deco2_reg_83(.CP(n_63198), .D(n_35434), .CD(n_62594), .Q
		(inst_deco2[83]));
	notech_mux2 i_37598(.S(n_56538), .A(inst_deco2[83]), .B(n_42378), .Z(n_35434
		));
	notech_reg inst_deco2_reg_84(.CP(n_63194), .D(n_35440), .CD(n_62596), .Q
		(inst_deco2[84]));
	notech_mux2 i_37606(.S(n_56538), .A(inst_deco2[84]), .B(n_42384), .Z(n_35440
		));
	notech_ao4 i_4827771(.A(n_59213), .B(n_42726), .C(n_55762), .D(n_43838),
		 .Z(n_2710));
	notech_reg inst_deco2_reg_85(.CP(n_63198), .D(n_35446), .CD(n_62600), .Q
		(inst_deco2[85]));
	notech_mux2 i_37614(.S(n_56543), .A(inst_deco2[85]), .B(n_42390), .Z(n_35446
		));
	notech_reg inst_deco2_reg_86(.CP(n_63194), .D(n_35452), .CD(n_62596), .Q
		(inst_deco2[86]));
	notech_mux2 i_37622(.S(n_56544), .A(inst_deco2[86]), .B(n_42396), .Z(n_35452
		));
	notech_reg inst_deco2_reg_87(.CP(n_63194), .D(n_35458), .CD(n_62596), .Q
		(inst_deco2[87]));
	notech_mux2 i_37630(.S(n_56544), .A(inst_deco2[87]), .B(n_42402), .Z(n_35458
		));
	notech_reg inst_deco2_reg_88(.CP(n_63194), .D(n_35464), .CD(n_62596), .Q
		(inst_deco2[88]));
	notech_mux2 i_37638(.S(n_56544), .A(inst_deco2[88]), .B(n_42408), .Z(n_35464
		));
	notech_and2 i_942(.A(n_3235), .B(in128[54]), .Z(n_2706));
	notech_reg inst_deco2_reg_89(.CP(n_63194), .D(n_35470), .CD(n_62600), .Q
		(inst_deco2[89]));
	notech_mux2 i_37646(.S(n_56544), .A(inst_deco2[89]), .B(n_42414), .Z(n_35470
		));
	notech_and4 i_58(.A(imm_sz[1]), .B(imm_sz[2]), .C(n_44371), .D(n_3079), 
		.Z(n_2705));
	notech_reg inst_deco2_reg_90(.CP(n_63194), .D(n_35476), .CD(n_62600), .Q
		(inst_deco2[90]));
	notech_mux2 i_37654(.S(n_56544), .A(inst_deco2[90]), .B(n_42420), .Z(n_35476
		));
	notech_or2 i_123154(.A(n_2701), .B(n_2702), .Z(n_2704));
	notech_reg inst_deco2_reg_91(.CP(n_63194), .D(n_35482), .CD(n_62600), .Q
		(inst_deco2[91]));
	notech_mux2 i_37662(.S(n_56544), .A(inst_deco2[91]), .B(n_42426), .Z(n_35482
		));
	notech_ao4 i_936(.A(n_5721), .B(n_2700), .C(db67), .D(n_43465), .Z(n_2703
		));
	notech_reg inst_deco2_reg_92(.CP(n_63194), .D(n_35488), .CD(n_62600), .Q
		(inst_deco2[92]));
	notech_mux2 i_37670(.S(n_56544), .A(inst_deco2[92]), .B(n_42432), .Z(n_35488
		));
	notech_ao3 i_939(.A(\to_acu2_0[4] ), .B(n_42556), .C(n_2703), .Z(n_2702)
		);
	notech_reg inst_deco2_reg_93(.CP(n_63194), .D(n_35494), .CD(n_62600), .Q
		(inst_deco2[93]));
	notech_mux2 i_37678(.S(n_56544), .A(inst_deco2[93]), .B(n_42438), .Z(n_35494
		));
	notech_nor2 i_938(.A(n_2858), .B(n_44729), .Z(n_2701));
	notech_reg inst_deco2_reg_94(.CP(n_63194), .D(n_35500), .CD(n_62596), .Q
		(inst_deco2[94]));
	notech_mux2 i_37686(.S(n_56544), .A(inst_deco2[94]), .B(n_42444), .Z(n_35500
		));
	notech_and2 i_934(.A(n_2867), .B(n_2698), .Z(n_2700));
	notech_reg inst_deco2_reg_95(.CP(n_63194), .D(n_35506), .CD(n_62596), .Q
		(inst_deco2[95]));
	notech_mux2 i_37694(.S(n_56544), .A(inst_deco2[95]), .B(n_42450), .Z(n_35506
		));
	notech_reg inst_deco2_reg_96(.CP(n_63194), .D(n_35512), .CD(n_62596), .Q
		(inst_deco2[96]));
	notech_mux2 i_37702(.S(n_56544), .A(inst_deco2[96]), .B(n_42456), .Z(n_35512
		));
	notech_nand3 i_935(.A(n_44747), .B(n_44748), .C(n_42548), .Z(n_2698));
	notech_reg inst_deco2_reg_97(.CP(n_63192), .D(n_35518), .CD(n_62596), .Q
		(inst_deco2[97]));
	notech_mux2 i_37710(.S(n_56544), .A(inst_deco2[97]), .B(n_42462), .Z(n_35518
		));
	notech_reg inst_deco2_reg_98(.CP(n_63187), .D(n_35524), .CD(n_62596), .Q
		(inst_deco2[98]));
	notech_mux2 i_37718(.S(n_56544), .A(inst_deco2[98]), .B(n_42468), .Z(n_35524
		));
	notech_and4 i_222691(.A(n_60367), .B(n_2975), .C(n_60854), .D(n_44524), 
		.Z(n_2696));
	notech_reg inst_deco2_reg_99(.CP(n_63187), .D(n_35530), .CD(n_62596), .Q
		(inst_deco2[99]));
	notech_mux2 i_37726(.S(n_56543), .A(inst_deco2[99]), .B(n_42474), .Z(n_35530
		));
	notech_nand2 i_211454(.A(n_3029), .B(start), .Z(n_2695));
	notech_reg inst_deco2_reg_100(.CP(n_63187), .D(n_35536), .CD(n_62596), .Q
		(inst_deco2[100]));
	notech_mux2 i_37734(.S(n_56543), .A(inst_deco2[100]), .B(n_42480), .Z(n_35536
		));
	notech_reg inst_deco2_reg_101(.CP(n_63187), .D(n_35542), .CD(n_62596), .Q
		(inst_deco2[101]));
	notech_mux2 i_37742(.S(n_56543), .A(inst_deco2[101]), .B(n_42486), .Z(n_35542
		));
	notech_reg inst_deco2_reg_102(.CP(n_63187), .D(n_35548), .CD(n_62596), .Q
		(inst_deco2[102]));
	notech_mux2 i_37750(.S(n_56543), .A(inst_deco2[102]), .B(n_42492), .Z(n_35548
		));
	notech_and2 i_890(.A(n_3245), .B(in128[63]), .Z(n_2692));
	notech_reg inst_deco2_reg_103(.CP(n_63187), .D(n_35554), .CD(n_62596), .Q
		(inst_deco2[103]));
	notech_mux2 i_37758(.S(n_56543), .A(inst_deco2[103]), .B(n_42498), .Z(n_35554
		));
	notech_reg inst_deco2_reg_104(.CP(n_63187), .D(n_35560), .CD(n_62596), .Q
		(inst_deco2[104]));
	notech_mux2 i_37766(.S(n_56543), .A(inst_deco2[104]), .B(n_42504), .Z(n_35560
		));
	notech_reg inst_deco2_reg_105(.CP(n_63187), .D(n_35566), .CD(n_62589), .Q
		(inst_deco2[105]));
	notech_mux2 i_37774(.S(n_56543), .A(inst_deco2[105]), .B(n_42510), .Z(n_35566
		));
	notech_and2 i_885(.A(n_3245), .B(in128[62]), .Z(n_2689));
	notech_reg inst_deco2_reg_106(.CP(n_63187), .D(n_35572), .CD(n_62589), .Q
		(inst_deco2[106]));
	notech_mux2 i_37782(.S(n_56544), .A(inst_deco2[106]), .B(n_42516), .Z(n_35572
		));
	notech_reg inst_deco2_reg_107(.CP(n_63187), .D(n_35578), .CD(n_62589), .Q
		(inst_deco2[107]));
	notech_mux2 i_37790(.S(n_56544), .A(inst_deco2[107]), .B(n_42522), .Z(n_35578
		));
	notech_reg inst_deco2_reg_108(.CP(n_63187), .D(n_35584), .CD(n_62589), .Q
		(inst_deco2[108]));
	notech_mux2 i_37798(.S(n_56544), .A(inst_deco2[108]), .B(n_42528), .Z(n_35584
		));
	notech_and2 i_880(.A(n_3245), .B(in128[61]), .Z(n_2686));
	notech_reg inst_deco2_reg_109(.CP(n_63187), .D(n_35590), .CD(n_62589), .Q
		(inst_deco2[109]));
	notech_mux2 i_37806(.S(n_56543), .A(inst_deco2[109]), .B(n_42534), .Z(n_35590
		));
	notech_reg inst_deco2_reg_110(.CP(n_63187), .D(n_35596), .CD(n_62589), .Q
		(inst_deco2[110]));
	notech_mux2 i_37814(.S(n_56544), .A(inst_deco2[110]), .B(n_42540), .Z(n_35596
		));
	notech_reg inst_deco2_reg_111(.CP(n_63187), .D(n_35602), .CD(n_62589), .Q
		(inst_deco2[111]));
	notech_mux2 i_37822(.S(n_56544), .A(inst_deco2[111]), .B(n_42546), .Z(n_35602
		));
	notech_and2 i_875(.A(n_3245), .B(in128[60]), .Z(n_2683));
	notech_reg inst_deco2_reg_112(.CP(n_63184), .D(n_35608), .CD(n_62589), .Q
		(inst_deco2[112]));
	notech_mux2 i_37830(.S(n_56527), .A(inst_deco2[112]), .B(n_42552), .Z(n_35608
		));
	notech_reg inst_deco2_reg_113(.CP(n_63184), .D(n_35614), .CD(n_62589), .Q
		(inst_deco2[113]));
	notech_mux2 i_37838(.S(n_56527), .A(inst_deco2[113]), .B(n_42558), .Z(n_35614
		));
	notech_reg inst_deco2_reg_114(.CP(n_63187), .D(n_35620), .CD(n_62589), .Q
		(inst_deco2[114]));
	notech_mux2 i_37846(.S(n_56527), .A(inst_deco2[114]), .B(n_42564), .Z(n_35620
		));
	notech_and2 i_870(.A(n_3245), .B(in128[59]), .Z(n_2680));
	notech_reg inst_deco2_reg_115(.CP(n_63187), .D(n_35626), .CD(n_62589), .Q
		(inst_deco2[115]));
	notech_mux2 i_37854(.S(n_56527), .A(inst_deco2[115]), .B(n_42570), .Z(n_35626
		));
	notech_reg inst_deco2_reg_116(.CP(n_63187), .D(n_35632), .CD(n_62589), .Q
		(inst_deco2[116]));
	notech_mux2 i_37862(.S(n_56527), .A(inst_deco2[116]), .B(n_42576), .Z(n_35632
		));
	notech_reg inst_deco2_reg_117(.CP(n_63187), .D(n_35638), .CD(n_62589), .Q
		(inst_deco2[117]));
	notech_mux2 i_37870(.S(n_56527), .A(inst_deco2[117]), .B(n_42582), .Z(n_35638
		));
	notech_and2 i_865(.A(n_3245), .B(in128[58]), .Z(n_2677));
	notech_reg inst_deco2_reg_118(.CP(n_63187), .D(n_35644), .CD(n_62586), .Q
		(inst_deco2[118]));
	notech_mux2 i_37878(.S(n_56527), .A(inst_deco2[118]), .B(n_42588), .Z(n_35644
		));
	notech_reg inst_deco2_reg_119(.CP(n_63189), .D(n_35650), .CD(n_62586), .Q
		(inst_deco2[119]));
	notech_mux2 i_37886(.S(n_56532), .A(inst_deco2[119]), .B(n_42594), .Z(n_35650
		));
	notech_reg inst_deco2_reg_120(.CP(n_63189), .D(n_35656), .CD(n_62586), .Q
		(inst_deco2[120]));
	notech_mux2 i_37894(.S(n_56532), .A(inst_deco2[120]), .B(n_42600), .Z(n_35656
		));
	notech_and2 i_860(.A(n_3245), .B(in128[57]), .Z(n_2674));
	notech_reg inst_deco2_reg_121(.CP(n_63189), .D(n_35662), .CD(n_62589), .Q
		(inst_deco2[121]));
	notech_mux2 i_37902(.S(n_56532), .A(inst_deco2[121]), .B(n_42606), .Z(n_35662
		));
	notech_reg inst_deco2_reg_122(.CP(n_63189), .D(n_35668), .CD(n_62589), .Q
		(inst_deco2[122]));
	notech_mux2 i_37910(.S(n_56527), .A(inst_deco2[122]), .B(n_42612), .Z(n_35668
		));
	notech_reg inst_deco2_reg_123(.CP(n_63189), .D(n_35674), .CD(n_62589), .Q
		(inst_deco2[123]));
	notech_mux2 i_37918(.S(n_56527), .A(inst_deco2[123]), .B(n_42618), .Z(n_35674
		));
	notech_and2 i_855(.A(n_3245), .B(in128[56]), .Z(n_2671));
	notech_reg inst_deco2_reg_124(.CP(n_63189), .D(n_35680), .CD(n_62589), .Q
		(inst_deco2[124]));
	notech_mux2 i_37926(.S(n_56532), .A(inst_deco2[124]), .B(n_42624), .Z(n_35680
		));
	notech_or2 i_854(.A(n_3245), .B(n_2705), .Z(n_2670));
	notech_reg inst_deco2_reg_125(.CP(n_63192), .D(n_35686), .CD(n_62589), .Q
		(inst_deco2[125]));
	notech_mux2 i_37934(.S(n_56522), .A(inst_deco2[125]), .B(n_42630), .Z(n_35686
		));
	notech_reg inst_deco2_reg_126(.CP(n_63189), .D(n_35692), .CD(n_62591), .Q
		(inst_deco2[126]));
	notech_mux2 i_37942(.S(n_56522), .A(inst_deco2[126]), .B(n_42636), .Z(n_35692
		));
	notech_reg inst_deco2_reg_127(.CP(n_63189), .D(n_35698), .CD(n_62591), .Q
		(inst_deco2[127]));
	notech_mux2 i_37950(.S(n_56522), .A(inst_deco2[127]), .B(n_42642), .Z(n_35698
		));
	notech_and2 i_848(.A(n_3235), .B(in128[55]), .Z(n_2667));
	notech_reg inst_deco1_reg_0(.CP(n_63189), .D(n_35704), .CD(n_62591), .Q(inst_deco1
		[0]));
	notech_mux2 i_37958(.S(n_59377), .A(inst_deco1[0]), .B(n_43077), .Z(n_35704
		));
	notech_reg inst_deco1_reg_1(.CP(n_63189), .D(n_35710), .CD(n_62591), .Q(inst_deco1
		[1]));
	notech_mux2 i_37966(.S(n_59377), .A(inst_deco1[1]), .B(n_43308), .Z(n_35710
		));
	notech_reg inst_deco1_reg_2(.CP(n_63189), .D(n_35716), .CD(n_62591), .Q(inst_deco1
		[2]));
	notech_mux2 i_37974(.S(n_59377), .A(inst_deco1[2]), .B(n_43310), .Z(n_35716
		));
	notech_and2 i_843(.A(n_3235), .B(in128[53]), .Z(n_2664));
	notech_reg inst_deco1_reg_3(.CP(n_63189), .D(n_35722), .CD(n_62594), .Q(inst_deco1
		[3]));
	notech_mux2 i_37982(.S(n_59377), .A(inst_deco1[3]), .B(n_43313), .Z(n_35722
		));
	notech_reg inst_deco1_reg_4(.CP(n_63189), .D(n_35728), .CD(n_62594), .Q(inst_deco1
		[4]));
	notech_mux2 i_37990(.S(n_59377), .A(inst_deco1[4]), .B(n_43315), .Z(n_35728
		));
	notech_reg inst_deco1_reg_5(.CP(n_63189), .D(n_35734), .CD(n_62594), .Q(inst_deco1
		[5]));
	notech_mux2 i_37998(.S(n_59355), .A(inst_deco1[5]), .B(n_43091), .Z(n_35734
		));
	notech_and2 i_838(.A(n_3235), .B(in128[52]), .Z(n_2661));
	notech_reg inst_deco1_reg_6(.CP(n_63189), .D(n_35740), .CD(n_62591), .Q(inst_deco1
		[6]));
	notech_mux2 i_38006(.S(n_59355), .A(inst_deco1[6]), .B(n_43317), .Z(n_35740
		));
	notech_reg inst_deco1_reg_7(.CP(n_63189), .D(n_35746), .CD(n_62591), .Q(inst_deco1
		[7]));
	notech_mux2 i_38014(.S(n_59355), .A(inst_deco1[7]), .B(n_43095), .Z(n_35746
		));
	notech_reg inst_deco1_reg_8(.CP(n_63189), .D(n_35752), .CD(n_62591), .Q(inst_deco1
		[8]));
	notech_mux2 i_38022(.S(n_59355), .A(inst_deco1[8]), .B(n_43099), .Z(n_35752
		));
	notech_and2 i_833(.A(n_3235), .B(in128[51]), .Z(n_2658));
	notech_reg inst_deco1_reg_9(.CP(n_63189), .D(n_35758), .CD(n_62591), .Q(inst_deco1
		[9]));
	notech_mux2 i_38030(.S(n_59355), .A(inst_deco1[9]), .B(n_43320), .Z(n_35758
		));
	notech_reg inst_deco1_reg_10(.CP(n_63189), .D(n_35764), .CD(n_62591), .Q
		(inst_deco1[10]));
	notech_mux2 i_38038(.S(n_59355), .A(inst_deco1[10]), .B(n_43322), .Z(n_35764
		));
	notech_reg inst_deco1_reg_11(.CP(n_63189), .D(n_35770), .CD(n_62591), .Q
		(inst_deco1[11]));
	notech_mux2 i_38046(.S(n_59355), .A(inst_deco1[11]), .B(n_43325), .Z(n_35770
		));
	notech_and2 i_828(.A(n_3235), .B(in128[50]), .Z(n_2655));
	notech_reg inst_deco1_reg_12(.CP(n_63205), .D(n_35776), .CD(n_62591), .Q
		(inst_deco1[12]));
	notech_mux2 i_38054(.S(n_59360), .A(inst_deco1[12]), .B(n_43326), .Z(n_35776
		));
	notech_reg inst_deco1_reg_13(.CP(n_63205), .D(n_35782), .CD(n_62591), .Q
		(inst_deco1[13]));
	notech_mux2 i_38062(.S(n_59360), .A(inst_deco1[13]), .B(n_43328), .Z(n_35782
		));
	notech_reg inst_deco1_reg_14(.CP(n_63205), .D(n_35788), .CD(n_62591), .Q
		(inst_deco1[14]));
	notech_mux2 i_38070(.S(n_59360), .A(inst_deco1[14]), .B(n_43331), .Z(n_35788
		));
	notech_and2 i_823(.A(n_3235), .B(in128[49]), .Z(n_2652));
	notech_reg inst_deco1_reg_15(.CP(n_63203), .D(n_35794), .CD(n_62591), .Q
		(inst_deco1[15]));
	notech_mux2 i_38078(.S(n_59355), .A(inst_deco1[15]), .B(n_43333), .Z(n_35794
		));
	notech_reg inst_deco1_reg_16(.CP(n_63203), .D(n_35800), .CD(n_62591), .Q
		(inst_deco1[16]));
	notech_mux2 i_38086(.S(n_59360), .A(inst_deco1[16]), .B(n_43335), .Z(n_35800
		));
	notech_reg inst_deco1_reg_17(.CP(n_63205), .D(n_35806), .CD(n_62591), .Q
		(inst_deco1[17]));
	notech_mux2 i_38094(.S(n_59360), .A(inst_deco1[17]), .B(n_43338), .Z(n_35806
		));
	notech_and2 i_818(.A(n_3235), .B(in128[48]), .Z(n_2649));
	notech_reg inst_deco1_reg_18(.CP(n_63205), .D(n_35812), .CD(n_62591), .Q
		(inst_deco1[18]));
	notech_mux2 i_38102(.S(n_59355), .A(inst_deco1[18]), .B(n_43340), .Z(n_35812
		));
	notech_or2 i_817(.A(n_3235), .B(n_2705), .Z(n_2648));
	notech_reg inst_deco1_reg_19(.CP(n_63205), .D(n_35818), .CD(n_62600), .Q
		(inst_deco1[19]));
	notech_mux2 i_38110(.S(n_59355), .A(inst_deco1[19]), .B(n_43341), .Z(n_35818
		));
	notech_nor2 i_830119(.A(imm_sz[1]), .B(n_44371), .Z(n_2647));
	notech_reg inst_deco1_reg_20(.CP(n_63205), .D(n_35824), .CD(n_62607), .Q
		(inst_deco1[20]));
	notech_mux2 i_38118(.S(n_59355), .A(inst_deco1[20]), .B(n_43344), .Z(n_35824
		));
	notech_or2 i_810(.A(n_3162), .B(n_44552), .Z(n_2646));
	notech_reg inst_deco1_reg_21(.CP(n_63205), .D(n_35830), .CD(n_62607), .Q
		(inst_deco1[21]));
	notech_mux2 i_38126(.S(n_59354), .A(inst_deco1[21]), .B(n_43346), .Z(n_35830
		));
	notech_reg inst_deco1_reg_22(.CP(n_63203), .D(n_35836), .CD(n_62607), .Q
		(inst_deco1[22]));
	notech_mux2 i_38134(.S(n_59354), .A(inst_deco1[22]), .B(n_43349), .Z(n_35836
		));
	notech_reg inst_deco1_reg_23(.CP(n_63203), .D(n_35842), .CD(n_62607), .Q
		(inst_deco1[23]));
	notech_mux2 i_38142(.S(n_59354), .A(inst_deco1[23]), .B(n_43351), .Z(n_35842
		));
	notech_and4 i_811(.A(n_3232), .B(n_2646), .C(n_2639), .D(n_3230), .Z(n_2643
		));
	notech_reg inst_deco1_reg_24(.CP(n_63203), .D(n_35848), .CD(n_62607), .Q
		(inst_deco1[24]));
	notech_mux2 i_38150(.S(n_59355), .A(inst_deco1[24]), .B(n_43353), .Z(n_35848
		));
	notech_or2 i_804(.A(n_3155), .B(n_44571), .Z(n_2642));
	notech_reg inst_deco1_reg_25(.CP(n_63203), .D(n_35854), .CD(n_62607), .Q
		(inst_deco1[25]));
	notech_mux2 i_38158(.S(n_59355), .A(inst_deco1[25]), .B(n_43356), .Z(n_35854
		));
	notech_reg inst_deco1_reg_26(.CP(n_63203), .D(n_35860), .CD(n_62607), .Q
		(inst_deco1[26]));
	notech_mux2 i_38166(.S(n_59355), .A(inst_deco1[26]), .B(n_43358), .Z(n_35860
		));
	notech_reg inst_deco1_reg_27(.CP(n_63203), .D(n_35866), .CD(n_62607), .Q
		(inst_deco1[27]));
	notech_mux2 i_38174(.S(n_59355), .A(inst_deco1[27]), .B(n_43361), .Z(n_35866
		));
	notech_or2 i_805(.A(n_3198), .B(n_44562), .Z(n_2639));
	notech_reg inst_deco1_reg_28(.CP(n_63203), .D(n_35872), .CD(n_62607), .Q
		(inst_deco1[28]));
	notech_mux2 i_38182(.S(n_59355), .A(inst_deco1[28]), .B(n_43363), .Z(n_35872
		));
	notech_or2 i_797(.A(n_3162), .B(n_44551), .Z(n_2638));
	notech_reg inst_deco1_reg_29(.CP(n_63203), .D(n_35878), .CD(n_62607), .Q
		(inst_deco1[29]));
	notech_mux2 i_38190(.S(n_59355), .A(inst_deco1[29]), .B(n_43365), .Z(n_35878
		));
	notech_reg inst_deco1_reg_30(.CP(n_63203), .D(n_35884), .CD(n_62605), .Q
		(inst_deco1[30]));
	notech_mux2 i_38198(.S(n_59355), .A(inst_deco1[30]), .B(n_43368), .Z(n_35884
		));
	notech_reg inst_deco1_reg_31(.CP(n_63203), .D(n_35890), .CD(n_62605), .Q
		(inst_deco1[31]));
	notech_mux2 i_38206(.S(n_59360), .A(inst_deco1[31]), .B(n_43370), .Z(n_35890
		));
	notech_and4 i_798(.A(n_3227), .B(n_2638), .C(n_2631), .D(n_3225), .Z(n_2635
		));
	notech_reg inst_deco1_reg_32(.CP(n_63203), .D(n_35896), .CD(n_62605), .Q
		(inst_deco1[32]));
	notech_mux2 i_38214(.S(n_59365), .A(inst_deco1[32]), .B(n_43373), .Z(n_35896
		));
	notech_or2 i_791(.A(n_3155), .B(n_44570), .Z(n_2634));
	notech_reg inst_deco1_reg_33(.CP(n_63208), .D(n_35902), .CD(n_62605), .Q
		(inst_deco1[33]));
	notech_mux2 i_38222(.S(n_59365), .A(inst_deco1[33]), .B(n_43375), .Z(n_35902
		));
	notech_reg inst_deco1_reg_34(.CP(n_63208), .D(n_35908), .CD(n_62605), .Q
		(inst_deco1[34]));
	notech_mux2 i_38230(.S(n_59365), .A(inst_deco1[34]), .B(n_43376), .Z(n_35908
		));
	notech_reg inst_deco1_reg_35(.CP(n_63208), .D(n_35914), .CD(n_62605), .Q
		(inst_deco1[35]));
	notech_mux2 i_38238(.S(n_59365), .A(inst_deco1[35]), .B(n_43380), .Z(n_35914
		));
	notech_or2 i_792(.A(n_3198), .B(n_44560), .Z(n_2631));
	notech_reg inst_deco1_reg_36(.CP(n_63205), .D(n_35920), .CD(n_62605), .Q
		(inst_deco1[36]));
	notech_mux2 i_38246(.S(n_59365), .A(inst_deco1[36]), .B(n_43381), .Z(n_35920
		));
	notech_or2 i_784(.A(n_3162), .B(n_44550), .Z(n_2630));
	notech_reg inst_deco1_reg_37(.CP(n_63208), .D(n_35926), .CD(n_62605), .Q
		(inst_deco1[37]));
	notech_mux2 i_38254(.S(n_59365), .A(inst_deco1[37]), .B(n_43382), .Z(n_35926
		));
	notech_reg inst_deco1_reg_38(.CP(n_63208), .D(n_35932), .CD(n_62605), .Q
		(inst_deco1[38]));
	notech_mux2 i_38262(.S(n_59365), .A(inst_deco1[38]), .B(n_43383), .Z(n_35932
		));
	notech_reg inst_deco1_reg_39(.CP(n_63208), .D(n_35938), .CD(n_62605), .Q
		(inst_deco1[39]));
	notech_mux2 i_38270(.S(n_59365), .A(inst_deco1[39]), .B(n_43385), .Z(n_35938
		));
	notech_and4 i_785(.A(n_3222), .B(n_2630), .C(n_2623), .D(n_3220), .Z(n_2627
		));
	notech_reg inst_deco1_reg_40(.CP(n_63208), .D(n_35944), .CD(n_62605), .Q
		(inst_deco1[40]));
	notech_mux2 i_38278(.S(n_59366), .A(inst_deco1[40]), .B(n_43386), .Z(n_35944
		));
	notech_or2 i_778(.A(n_3155), .B(n_44569), .Z(n_2626));
	notech_reg inst_deco1_reg_41(.CP(n_63208), .D(n_35950), .CD(n_62610), .Q
		(inst_deco1[41]));
	notech_mux2 i_38286(.S(n_59366), .A(inst_deco1[41]), .B(n_43176), .Z(n_35950
		));
	notech_reg inst_deco1_reg_42(.CP(n_63208), .D(n_35956), .CD(n_62610), .Q
		(inst_deco1[42]));
	notech_mux2 i_38294(.S(n_59365), .A(inst_deco1[42]), .B(n_43179), .Z(n_35956
		));
	notech_reg inst_deco1_reg_43(.CP(n_63205), .D(n_35962), .CD(n_62610), .Q
		(inst_deco1[43]));
	notech_mux2 i_38302(.S(n_59365), .A(inst_deco1[43]), .B(n_43182), .Z(n_35962
		));
	notech_or2 i_779(.A(n_3198), .B(n_44559), .Z(n_2623));
	notech_reg inst_deco1_reg_44(.CP(n_63205), .D(n_35968), .CD(n_62610), .Q
		(inst_deco1[44]));
	notech_mux2 i_38310(.S(n_59365), .A(inst_deco1[44]), .B(n_43185), .Z(n_35968
		));
	notech_or2 i_771(.A(n_3162), .B(n_44548), .Z(n_2622));
	notech_reg inst_deco1_reg_45(.CP(n_63205), .D(n_35974), .CD(n_62610), .Q
		(inst_deco1[45]));
	notech_mux2 i_38318(.S(n_59360), .A(inst_deco1[45]), .B(n_43188), .Z(n_35974
		));
	notech_reg inst_deco1_reg_46(.CP(n_63205), .D(n_35980), .CD(n_62610), .Q
		(inst_deco1[46]));
	notech_mux2 i_38326(.S(n_59360), .A(inst_deco1[46]), .B(n_43387), .Z(n_35980
		));
	notech_reg inst_deco1_reg_47(.CP(n_63205), .D(n_35986), .CD(n_62610), .Q
		(inst_deco1[47]));
	notech_mux2 i_38334(.S(n_59360), .A(inst_deco1[47]), .B(n_43388), .Z(n_35986
		));
	notech_and4 i_772(.A(n_3217), .B(n_2622), .C(n_2615), .D(n_3215), .Z(n_2619
		));
	notech_reg inst_deco1_reg_48(.CP(n_63205), .D(n_35992), .CD(n_62610), .Q
		(inst_deco1[48]));
	notech_mux2 i_38342(.S(n_59360), .A(inst_deco1[48]), .B(n_43389), .Z(n_35992
		));
	notech_or2 i_765(.A(n_3155), .B(n_44568), .Z(n_2618));
	notech_reg inst_deco1_reg_49(.CP(n_63205), .D(n_35998), .CD(n_62610), .Q
		(inst_deco1[49]));
	notech_mux2 i_38350(.S(n_59360), .A(inst_deco1[49]), .B(n_43391), .Z(n_35998
		));
	notech_reg inst_deco1_reg_50(.CP(n_63205), .D(n_36004), .CD(n_62610), .Q
		(inst_deco1[50]));
	notech_mux2 i_38358(.S(n_59360), .A(inst_deco1[50]), .B(n_43392), .Z(n_36004
		));
	notech_reg inst_deco1_reg_51(.CP(n_63205), .D(n_36010), .CD(n_62610), .Q
		(inst_deco1[51]));
	notech_mux2 i_38366(.S(n_59365), .A(inst_deco1[51]), .B(n_43393), .Z(n_36010
		));
	notech_or2 i_766(.A(n_3198), .B(n_44558), .Z(n_2615));
	notech_reg inst_deco1_reg_52(.CP(n_63205), .D(n_36016), .CD(n_62607), .Q
		(inst_deco1[52]));
	notech_mux2 i_38374(.S(n_59365), .A(inst_deco1[52]), .B(n_43394), .Z(n_36016
		));
	notech_or2 i_758(.A(n_3162), .B(n_44547), .Z(n_2614));
	notech_reg inst_deco1_reg_53(.CP(n_63205), .D(n_36022), .CD(n_62607), .Q
		(inst_deco1[53]));
	notech_mux2 i_38382(.S(n_59365), .A(inst_deco1[53]), .B(n_43395), .Z(n_36022
		));
	notech_reg inst_deco1_reg_54(.CP(n_63203), .D(n_36028), .CD(n_62607), .Q
		(inst_deco1[54]));
	notech_mux2 i_38390(.S(n_59365), .A(inst_deco1[54]), .B(n_43397), .Z(n_36028
		));
	notech_reg inst_deco1_reg_55(.CP(n_63198), .D(n_36034), .CD(n_62607), .Q
		(inst_deco1[55]));
	notech_mux2 i_38398(.S(n_59365), .A(inst_deco1[55]), .B(n_43398), .Z(n_36034
		));
	notech_and4 i_759(.A(n_3212), .B(n_2614), .C(n_2607), .D(n_3210), .Z(n_2611
		));
	notech_reg inst_deco1_reg_56(.CP(n_63198), .D(n_36040), .CD(n_62607), .Q
		(inst_deco1[56]));
	notech_mux2 i_38406(.S(n_59365), .A(inst_deco1[56]), .B(n_43400), .Z(n_36040
		));
	notech_or2 i_752(.A(n_3155), .B(n_44566), .Z(n_2610));
	notech_reg inst_deco1_reg_57(.CP(n_63198), .D(n_36046), .CD(n_62607), .Q
		(inst_deco1[57]));
	notech_mux2 i_38414(.S(n_59365), .A(inst_deco1[57]), .B(n_43404), .Z(n_36046
		));
	notech_reg inst_deco1_reg_58(.CP(n_63198), .D(n_36052), .CD(n_62607), .Q
		(inst_deco1[58]));
	notech_mux2 i_38422(.S(n_59378), .A(inst_deco1[58]), .B(n_43407), .Z(n_36052
		));
	notech_reg inst_deco1_reg_59(.CP(n_63198), .D(n_36058), .CD(n_62607), .Q
		(inst_deco1[59]));
	notech_mux2 i_38430(.S(n_59394), .A(inst_deco1[59]), .B(n_43411), .Z(n_36058
		));
	notech_or2 i_753(.A(n_3198), .B(n_44557), .Z(n_2607));
	notech_reg inst_deco1_reg_60(.CP(n_63200), .D(n_36064), .CD(n_62607), .Q
		(inst_deco1[60]));
	notech_mux2 i_38438(.S(n_59399), .A(inst_deco1[60]), .B(n_43413), .Z(n_36064
		));
	notech_or2 i_745(.A(n_3162), .B(n_44546), .Z(n_2606));
	notech_reg inst_deco1_reg_61(.CP(n_63200), .D(n_36070), .CD(n_62607), .Q
		(inst_deco1[61]));
	notech_mux2 i_38446(.S(n_59399), .A(inst_deco1[61]), .B(n_43415), .Z(n_36070
		));
	notech_reg inst_deco1_reg_62(.CP(n_63200), .D(n_36076), .CD(n_62602), .Q
		(inst_deco1[62]));
	notech_mux2 i_38454(.S(n_59394), .A(inst_deco1[62]), .B(n_43416), .Z(n_36076
		));
	notech_reg inst_deco1_reg_63(.CP(n_63200), .D(n_36082), .CD(n_62602), .Q
		(inst_deco1[63]));
	notech_mux2 i_38462(.S(n_59394), .A(inst_deco1[63]), .B(n_43417), .Z(n_36082
		));
	notech_and4 i_746(.A(n_3207), .B(n_2606), .C(n_2599), .D(n_3205), .Z(n_2603
		));
	notech_reg inst_deco1_reg_64(.CP(n_63200), .D(n_36088), .CD(n_62602), .Q
		(inst_deco1[64]));
	notech_mux2 i_38470(.S(n_59394), .A(inst_deco1[64]), .B(n_43418), .Z(n_36088
		));
	notech_or2 i_739(.A(n_3155), .B(n_44565), .Z(n_2602));
	notech_reg inst_deco1_reg_65(.CP(n_63198), .D(n_36094), .CD(n_62600), .Q
		(inst_deco1[65]));
	notech_mux2 i_38478(.S(n_59399), .A(inst_deco1[65]), .B(n_43419), .Z(n_36094
		));
	notech_reg inst_deco1_reg_66(.CP(n_63198), .D(n_36100), .CD(n_62600), .Q
		(inst_deco1[66]));
	notech_mux2 i_38486(.S(n_59399), .A(inst_deco1[66]), .B(n_43421), .Z(n_36100
		));
	notech_reg inst_deco1_reg_67(.CP(n_63198), .D(n_36106), .CD(n_62602), .Q
		(inst_deco1[67]));
	notech_mux2 i_38494(.S(n_59399), .A(inst_deco1[67]), .B(n_43422), .Z(n_36106
		));
	notech_or2 i_740(.A(n_3198), .B(n_44556), .Z(n_2599));
	notech_reg inst_deco1_reg_68(.CP(n_63198), .D(n_36112), .CD(n_62602), .Q
		(inst_deco1[68]));
	notech_mux2 i_38502(.S(n_59399), .A(inst_deco1[68]), .B(n_43423), .Z(n_36112
		));
	notech_or2 i_732(.A(n_3162), .B(n_44544), .Z(n_2598));
	notech_reg inst_deco1_reg_69(.CP(n_63198), .D(n_36118), .CD(n_62602), .Q
		(inst_deco1[69]));
	notech_mux2 i_38510(.S(n_59399), .A(inst_deco1[69]), .B(n_43424), .Z(n_36118
		));
	notech_reg inst_deco1_reg_70(.CP(n_63198), .D(n_36124), .CD(n_62602), .Q
		(inst_deco1[70]));
	notech_mux2 i_38518(.S(n_59399), .A(inst_deco1[70]), .B(n_43425), .Z(n_36124
		));
	notech_reg inst_deco1_reg_71(.CP(n_63198), .D(n_36130), .CD(n_62602), .Q
		(inst_deco1[71]));
	notech_mux2 i_38526(.S(n_59399), .A(inst_deco1[71]), .B(n_43427), .Z(n_36130
		));
	notech_and4 i_733(.A(n_3202), .B(n_2598), .C(n_2591), .D(n_3200), .Z(n_2595
		));
	notech_reg inst_deco1_reg_72(.CP(n_63198), .D(n_36136), .CD(n_62600), .Q
		(inst_deco1[72]));
	notech_mux2 i_38534(.S(n_59389), .A(inst_deco1[72]), .B(n_43429), .Z(n_36136
		));
	notech_or2 i_726(.A(n_3155), .B(n_44563), .Z(n_2594));
	notech_reg inst_deco1_reg_73(.CP(n_63198), .D(n_36142), .CD(n_62600), .Q
		(inst_deco1[73]));
	notech_mux2 i_38542(.S(n_59389), .A(inst_deco1[73]), .B(n_43430), .Z(n_36142
		));
	notech_reg inst_deco1_reg_74(.CP(n_63198), .D(n_36148), .CD(n_62600), .Q
		(inst_deco1[74]));
	notech_mux2 i_38550(.S(n_59394), .A(inst_deco1[74]), .B(n_43433), .Z(n_36148
		));
	notech_reg inst_deco1_reg_75(.CP(n_63198), .D(n_36154), .CD(n_62600), .Q
		(inst_deco1[75]));
	notech_mux2 i_38558(.S(n_59389), .A(inst_deco1[75]), .B(n_43435), .Z(n_36154
		));
	notech_or2 i_727(.A(n_3198), .B(n_44553), .Z(n_2591));
	notech_reg inst_deco1_reg_76(.CP(n_63200), .D(n_36160), .CD(n_62600), .Q
		(inst_deco1[76]));
	notech_mux2 i_38566(.S(n_59389), .A(inst_deco1[76]), .B(n_43436), .Z(n_36160
		));
	notech_nor2 i_722(.A(n_3197), .B(n_2647), .Z(n_2590));
	notech_reg inst_deco1_reg_77(.CP(n_63203), .D(n_36166), .CD(n_62600), .Q
		(inst_deco1[77]));
	notech_mux2 i_38574(.S(n_59389), .A(inst_deco1[77]), .B(n_43439), .Z(n_36166
		));
	notech_reg inst_deco1_reg_78(.CP(n_63200), .D(n_36172), .CD(n_62600), .Q
		(inst_deco1[78]));
	notech_mux2 i_38582(.S(n_59394), .A(inst_deco1[78]), .B(n_43440), .Z(n_36172
		));
	notech_or2 i_716(.A(n_3162), .B(n_44542), .Z(n_2588));
	notech_reg inst_deco1_reg_79(.CP(n_63200), .D(n_36178), .CD(n_62600), .Q
		(inst_deco1[79]));
	notech_mux2 i_38590(.S(n_59394), .A(inst_deco1[79]), .B(n_43442), .Z(n_36178
		));
	notech_reg inst_deco1_reg_80(.CP(n_63200), .D(n_36184), .CD(n_62600), .Q
		(inst_deco1[80]));
	notech_mux2 i_38598(.S(n_59394), .A(inst_deco1[80]), .B(n_43443), .Z(n_36184
		));
	notech_reg inst_deco1_reg_81(.CP(n_63203), .D(n_36190), .CD(n_62600), .Q
		(inst_deco1[81]));
	notech_mux2 i_38606(.S(n_59394), .A(inst_deco1[81]), .B(n_43447), .Z(n_36190
		));
	notech_and4 i_717(.A(n_3195), .B(n_2581), .C(n_2588), .D(n_3193), .Z(n_2585
		));
	notech_reg inst_deco1_reg_82(.CP(n_63203), .D(n_36196), .CD(n_62600), .Q
		(inst_deco1[82]));
	notech_mux2 i_38614(.S(n_59394), .A(inst_deco1[82]), .B(n_43451), .Z(n_36196
		));
	notech_or2 i_708(.A(n_3156), .B(n_44571), .Z(n_2584));
	notech_reg inst_deco1_reg_83(.CP(n_63203), .D(n_36202), .CD(n_62605), .Q
		(inst_deco1[83]));
	notech_mux2 i_38622(.S(n_59394), .A(inst_deco1[83]), .B(n_43452), .Z(n_36202
		));
	notech_reg inst_deco1_reg_84(.CP(n_63203), .D(n_36208), .CD(n_62605), .Q
		(inst_deco1[84]));
	notech_mux2 i_38630(.S(n_59394), .A(inst_deco1[84]), .B(n_43455), .Z(n_36208
		));
	notech_reg inst_deco1_reg_85(.CP(n_63203), .D(n_36214), .CD(n_62605), .Q
		(inst_deco1[85]));
	notech_mux2 i_38638(.S(n_59399), .A(inst_deco1[85]), .B(n_42586), .Z(n_36214
		));
	notech_or2 i_710(.A(n_3155), .B(n_44562), .Z(n_2581));
	notech_reg inst_deco1_reg_86(.CP(n_63200), .D(n_36220), .CD(n_62602), .Q
		(inst_deco1[86]));
	notech_mux2 i_38646(.S(n_59400), .A(inst_deco1[86]), .B(n_42587), .Z(n_36220
		));
	notech_or2 i_703(.A(n_3162), .B(n_44541), .Z(n_2580));
	notech_reg inst_deco1_reg_87(.CP(n_63200), .D(n_36226), .CD(n_62605), .Q
		(inst_deco1[87]));
	notech_mux2 i_38654(.S(n_59400), .A(inst_deco1[87]), .B(n_42589), .Z(n_36226
		));
	notech_reg inst_deco1_reg_88(.CP(n_63200), .D(n_36232), .CD(n_62605), .Q
		(inst_deco1[88]));
	notech_mux2 i_38662(.S(n_59400), .A(inst_deco1[88]), .B(n_42590), .Z(n_36232
		));
	notech_reg inst_deco1_reg_89(.CP(n_63200), .D(n_36238), .CD(n_62605), .Q
		(inst_deco1[89]));
	notech_mux2 i_38670(.S(n_59400), .A(inst_deco1[89]), .B(n_42591), .Z(n_36238
		));
	notech_and4 i_704(.A(n_3190), .B(n_2573), .C(n_2580), .D(n_3188), .Z(n_2577
		));
	notech_reg inst_deco1_reg_90(.CP(n_63200), .D(n_36244), .CD(n_62605), .Q
		(inst_deco1[90]));
	notech_mux2 i_38678(.S(n_59400), .A(inst_deco1[90]), .B(n_42592), .Z(n_36244
		));
	notech_or2 i_695(.A(n_3156), .B(n_44570), .Z(n_2576));
	notech_reg inst_deco1_reg_91(.CP(n_63200), .D(n_36250), .CD(n_62605), .Q
		(inst_deco1[91]));
	notech_mux2 i_38686(.S(n_59400), .A(inst_deco1[91]), .B(n_42593), .Z(n_36250
		));
	notech_reg inst_deco1_reg_92(.CP(n_63200), .D(n_36256), .CD(n_62605), .Q
		(inst_deco1[92]));
	notech_mux2 i_38694(.S(n_59400), .A(inst_deco1[92]), .B(n_42595), .Z(n_36256
		));
	notech_reg inst_deco1_reg_93(.CP(n_63200), .D(n_36262), .CD(n_62602), .Q
		(inst_deco1[93]));
	notech_mux2 i_38702(.S(n_59400), .A(inst_deco1[93]), .B(n_42596), .Z(n_36262
		));
	notech_or2 i_697(.A(n_3155), .B(n_44560), .Z(n_2573));
	notech_reg inst_deco1_reg_94(.CP(n_63200), .D(n_36268), .CD(n_62602), .Q
		(inst_deco1[94]));
	notech_mux2 i_38710(.S(n_59400), .A(inst_deco1[94]), .B(n_42597), .Z(n_36268
		));
	notech_or2 i_690(.A(n_3162), .B(n_44539), .Z(n_2572));
	notech_reg inst_deco1_reg_95(.CP(n_63200), .D(n_36274), .CD(n_62602), .Q
		(inst_deco1[95]));
	notech_mux2 i_38718(.S(n_59400), .A(inst_deco1[95]), .B(n_42598), .Z(n_36274
		));
	notech_reg inst_deco1_reg_96(.CP(n_63200), .D(n_36280), .CD(n_62602), .Q
		(inst_deco1[96]));
	notech_mux2 i_38726(.S(n_59400), .A(inst_deco1[96]), .B(n_43458), .Z(n_36280
		));
	notech_reg inst_deco1_reg_97(.CP(n_63231), .D(n_36286), .CD(n_62602), .Q
		(inst_deco1[97]));
	notech_mux2 i_38734(.S(n_59400), .A(inst_deco1[97]), .B(n_43460), .Z(n_36286
		));
	notech_and4 i_691(.A(n_3185), .B(n_2565), .C(n_2572), .D(n_3183), .Z(n_2569
		));
	notech_reg inst_deco1_reg_98(.CP(n_63263), .D(n_36292), .CD(n_62602), .Q
		(inst_deco1[98]));
	notech_mux2 i_38742(.S(n_59400), .A(inst_deco1[98]), .B(n_43463), .Z(n_36292
		));
	notech_or2 i_682(.A(n_3156), .B(n_44568), .Z(n_2568));
	notech_reg inst_deco1_reg_99(.CP(n_63263), .D(n_36298), .CD(n_62602), .Q
		(inst_deco1[99]));
	notech_mux2 i_38750(.S(n_59399), .A(inst_deco1[99]), .B(n_43467), .Z(n_36298
		));
	notech_reg inst_deco1_reg_100(.CP(n_63263), .D(n_36304), .CD(n_62602), .Q
		(inst_deco1[100]));
	notech_mux2 i_38758(.S(n_59399), .A(inst_deco1[100]), .B(n_43470), .Z(n_36304
		));
	notech_reg inst_deco1_reg_101(.CP(n_63263), .D(n_36310), .CD(n_62602), .Q
		(inst_deco1[101]));
	notech_mux2 i_38766(.S(n_59399), .A(inst_deco1[101]), .B(n_42599), .Z(n_36310
		));
	notech_or2 i_684(.A(n_3155), .B(n_44558), .Z(n_2565));
	notech_reg inst_deco1_reg_102(.CP(n_63263), .D(n_36316), .CD(n_62602), .Q
		(inst_deco1[102]));
	notech_mux2 i_38774(.S(n_59399), .A(inst_deco1[102]), .B(n_43472), .Z(n_36316
		));
	notech_or2 i_677(.A(n_3162), .B(n_44538), .Z(n_2564));
	notech_reg inst_deco1_reg_103(.CP(n_63263), .D(n_36322), .CD(n_62602), .Q
		(inst_deco1[103]));
	notech_mux2 i_38782(.S(n_59399), .A(inst_deco1[103]), .B(n_42601), .Z(n_36322
		));
	notech_reg inst_deco1_reg_104(.CP(n_63263), .D(n_36328), .CD(n_62665), .Q
		(inst_deco1[104]));
	notech_mux2 i_38790(.S(n_59399), .A(inst_deco1[104]), .B(n_43476), .Z(n_36328
		));
	notech_reg inst_deco1_reg_105(.CP(n_63263), .D(n_36334), .CD(n_62665), .Q
		(inst_deco1[105]));
	notech_mux2 i_38798(.S(n_59399), .A(inst_deco1[105]), .B(n_43479), .Z(n_36334
		));
	notech_and4 i_678(.A(n_3180), .B(n_2557), .C(n_2564), .D(n_3178), .Z(n_2561
		));
	notech_reg inst_deco1_reg_106(.CP(n_63263), .D(n_36340), .CD(n_62665), .Q
		(inst_deco1[106]));
	notech_mux2 i_38806(.S(n_59400), .A(inst_deco1[106]), .B(n_43483), .Z(n_36340
		));
	notech_or2 i_669(.A(n_3156), .B(n_44566), .Z(n_2560));
	notech_reg inst_deco1_reg_107(.CP(n_63263), .D(n_36346), .CD(n_62665), .Q
		(inst_deco1[107]));
	notech_mux2 i_38814(.S(n_59400), .A(inst_deco1[107]), .B(n_42603), .Z(n_36346
		));
	notech_reg inst_deco1_reg_108(.CP(n_63263), .D(n_36352), .CD(n_62665), .Q
		(inst_deco1[108]));
	notech_mux2 i_38822(.S(n_59400), .A(inst_deco1[108]), .B(n_43487), .Z(n_36352
		));
	notech_reg inst_deco1_reg_109(.CP(n_63259), .D(n_36358), .CD(n_62665), .Q
		(inst_deco1[109]));
	notech_mux2 i_38830(.S(n_59399), .A(inst_deco1[109]), .B(n_43490), .Z(n_36358
		));
	notech_or2 i_671(.A(n_3155), .B(n_44557), .Z(n_2557));
	notech_reg inst_deco1_reg_110(.CP(n_63259), .D(n_36364), .CD(n_62665), .Q
		(inst_deco1[110]));
	notech_mux2 i_38838(.S(n_59400), .A(inst_deco1[110]), .B(n_43493), .Z(n_36364
		));
	notech_or2 i_664(.A(n_3162), .B(n_44536), .Z(n_2556));
	notech_reg inst_deco1_reg_111(.CP(n_63259), .D(n_36370), .CD(n_62665), .Q
		(inst_deco1[111]));
	notech_mux2 i_38846(.S(n_59400), .A(inst_deco1[111]), .B(n_43496), .Z(n_36370
		));
	notech_reg inst_deco1_reg_112(.CP(n_63259), .D(n_36376), .CD(n_62665), .Q
		(inst_deco1[112]));
	notech_mux2 i_38854(.S(n_59383), .A(inst_deco1[112]), .B(n_43500), .Z(n_36376
		));
	notech_reg inst_deco1_reg_113(.CP(n_63259), .D(n_36382), .CD(n_62665), .Q
		(inst_deco1[113]));
	notech_mux2 i_38862(.S(n_59383), .A(inst_deco1[113]), .B(n_42605), .Z(n_36382
		));
	notech_and4 i_665(.A(n_3175), .B(n_2549), .C(n_2556), .D(n_3173), .Z(n_2553
		));
	notech_reg inst_deco1_reg_114(.CP(n_63263), .D(n_36388), .CD(n_62665), .Q
		(inst_deco1[114]));
	notech_mux2 i_38870(.S(n_59383), .A(inst_deco1[114]), .B(n_42607), .Z(n_36388
		));
	notech_or2 i_656(.A(n_3156), .B(n_44565), .Z(n_2552));
	notech_reg inst_deco1_reg_115(.CP(n_63263), .D(n_36394), .CD(n_62661), .Q
		(inst_deco1[115]));
	notech_mux2 i_38878(.S(n_59383), .A(inst_deco1[115]), .B(n_42608), .Z(n_36394
		));
	notech_reg inst_deco1_reg_116(.CP(n_63263), .D(n_36400), .CD(n_62661), .Q
		(inst_deco1[116]));
	notech_mux2 i_38886(.S(n_59383), .A(inst_deco1[116]), .B(n_43503), .Z(n_36400
		));
	notech_reg inst_deco1_reg_117(.CP(n_63259), .D(n_36406), .CD(n_62661), .Q
		(inst_deco1[117]));
	notech_mux2 i_38894(.S(n_59383), .A(inst_deco1[117]), .B(n_43507), .Z(n_36406
		));
	notech_or2 i_658(.A(n_3155), .B(n_44556), .Z(n_2549));
	notech_reg inst_deco1_reg_118(.CP(n_63259), .D(n_36412), .CD(n_62661), .Q
		(inst_deco1[118]));
	notech_mux2 i_38902(.S(n_59383), .A(inst_deco1[118]), .B(n_42609), .Z(n_36412
		));
	notech_or2 i_651(.A(n_3162), .B(n_44535), .Z(n_2548));
	notech_reg inst_deco1_reg_119(.CP(n_63265), .D(n_36418), .CD(n_62661), .Q
		(inst_deco1[119]));
	notech_mux2 i_38910(.S(n_59388), .A(inst_deco1[119]), .B(n_43509), .Z(n_36418
		));
	notech_reg inst_deco1_reg_120(.CP(n_63265), .D(n_36424), .CD(n_62665), .Q
		(inst_deco1[120]));
	notech_mux2 i_38918(.S(n_59388), .A(inst_deco1[120]), .B(n_42610), .Z(n_36424
		));
	notech_reg inst_deco1_reg_121(.CP(n_63265), .D(n_36430), .CD(n_62665), .Q
		(inst_deco1[121]));
	notech_mux2 i_38926(.S(n_59388), .A(inst_deco1[121]), .B(n_43512), .Z(n_36430
		));
	notech_and4 i_652(.A(n_3170), .B(n_2541), .C(n_2548), .D(n_3168), .Z(n_2545
		));
	notech_reg inst_deco1_reg_122(.CP(n_63265), .D(n_36436), .CD(n_62665), .Q
		(inst_deco1[122]));
	notech_mux2 i_38934(.S(n_59383), .A(inst_deco1[122]), .B(n_42614), .Z(n_36436
		));
	notech_or2 i_643(.A(n_3156), .B(n_44564), .Z(n_2544));
	notech_reg inst_deco1_reg_123(.CP(n_63265), .D(n_36442), .CD(n_62661), .Q
		(inst_deco1[123]));
	notech_mux2 i_38942(.S(n_59383), .A(inst_deco1[123]), .B(n_43514), .Z(n_36442
		));
	notech_reg inst_deco1_reg_124(.CP(n_63265), .D(n_36448), .CD(n_62661), .Q
		(inst_deco1[124]));
	notech_mux2 i_38950(.S(n_59388), .A(inst_deco1[124]), .B(n_42615), .Z(n_36448
		));
	notech_reg inst_deco1_reg_125(.CP(n_63265), .D(n_36454), .CD(n_62670), .Q
		(inst_deco1[125]));
	notech_mux2 i_38958(.S(n_59378), .A(inst_deco1[125]), .B(n_43517), .Z(n_36454
		));
	notech_or2 i_645(.A(n_3155), .B(n_44554), .Z(n_2541));
	notech_reg inst_deco1_reg_126(.CP(n_63265), .D(n_36460), .CD(n_62670), .Q
		(inst_deco1[126]));
	notech_mux2 i_38966(.S(n_59378), .A(inst_deco1[126]), .B(n_42619), .Z(n_36460
		));
	notech_or2 i_638(.A(n_3162), .B(n_44534), .Z(n_2540));
	notech_reg inst_deco1_reg_127(.CP(n_63265), .D(n_36466), .CD(n_62670), .Q
		(inst_deco1[127]));
	notech_mux2 i_38974(.S(n_59378), .A(inst_deco1[127]), .B(n_42620), .Z(n_36466
		));
	notech_reg trig_it_reg(.CP(n_63265), .D(n_36472), .CD(n_62670), .Q(trig_it
		));
	notech_mux2 i_38982(.S(n_3297), .A(n_42613), .B(trig_it), .Z(n_36472));
	notech_reg trig_itf_reg(.CP(n_63265), .D(trig_it), .CD(n_62670), .Q(trig_itf
		));
	notech_reg intf_reg(.CP(n_63263), .D(int_main), .CD(n_62678), .Q(intf)
		);
	notech_reg_set intff_reg(.CP(n_63263), .D(n_36482), .SD(1'b1), .Q(intff)
		);
	notech_mux2 i_38998(.S(n_62678), .A(intff), .B(intf), .Z(n_36482));
	notech_and4 i_639(.A(n_3165), .B(n_2533), .C(n_2540), .D(n_3160), .Z(n_2537
		));
	notech_reg ififo_rvect4_reg_0(.CP(n_63263), .D(n_36488), .CD(n_62678), .Q
		(ififo_rvect4[0]));
	notech_mux2 i_39006(.S(\nbus_13546[0] ), .A(ififo_rvect4[0]), .B(n_1534100839
		), .Z(n_36488));
	notech_or2 i_630(.A(n_3156), .B(n_44563), .Z(n_2536));
	notech_reg ififo_rvect4_reg_1(.CP(n_63263), .D(n_36494), .CD(n_62678), .Q
		(ififo_rvect4[1]));
	notech_mux2 i_39014(.S(\nbus_13546[0] ), .A(ififo_rvect4[1]), .B(n_1535100840
		), .Z(n_36494));
	notech_reg ififo_rvect4_reg_2(.CP(n_63263), .D(n_36500), .CD(n_62678), .Q
		(ififo_rvect4[2]));
	notech_mux2 i_39022(.S(\nbus_13546[0] ), .A(ififo_rvect4[2]), .B(n_1536100841
		), .Z(n_36500));
	notech_reg ififo_rvect4_reg_3(.CP(n_63265), .D(n_36506), .CD(n_62670), .Q
		(ififo_rvect4[3]));
	notech_mux2 i_39030(.S(\nbus_13546[0] ), .A(ififo_rvect4[3]), .B(n_1537100842
		), .Z(n_36506));
	notech_or2 i_632(.A(n_3155), .B(n_44553), .Z(n_2533));
	notech_reg ififo_rvect4_reg_4(.CP(n_63265), .D(n_36512), .CD(n_62665), .Q
		(ififo_rvect4[4]));
	notech_mux2 i_39038(.S(\nbus_13546[0] ), .A(ififo_rvect4[4]), .B(n_1538100843
		), .Z(n_36512));
	notech_nor2 i_629(.A(n_3117), .B(n_3131), .Z(n_2532));
	notech_reg ififo_rvect4_reg_5(.CP(n_63265), .D(n_36518), .CD(n_62665), .Q
		(ififo_rvect4[5]));
	notech_mux2 i_39046(.S(\nbus_13546[0] ), .A(ififo_rvect4[5]), .B(n_1539100844
		), .Z(n_36518));
	notech_nand2 i_628(.A(n_3121), .B(n_44105), .Z(n_2531));
	notech_reg ififo_rvect4_reg_6(.CP(n_63263), .D(n_36524), .CD(n_62665), .Q
		(ififo_rvect4[6]));
	notech_mux2 i_39054(.S(\nbus_13546[0] ), .A(ififo_rvect4[6]), .B(n_1540100845
		), .Z(n_36524));
	notech_or2 i_623(.A(n_3129), .B(n_44552), .Z(n_2530));
	notech_reg ififo_rvect4_reg_7(.CP(n_63265), .D(n_36530), .CD(n_62665), .Q
		(ififo_rvect4[7]));
	notech_mux2 i_39062(.S(\nbus_13546[0] ), .A(ififo_rvect4[7]), .B(n_1541100846
		), .Z(n_36530));
	notech_reg ififo_rvect3_reg_0(.CP(n_63259), .D(n_36536), .CD(n_62665), .Q
		(ififo_rvect3[0]));
	notech_mux2 i_39070(.S(\nbus_13546[0] ), .A(ififo_rvect3[0]), .B(n_46038
		), .Z(n_36536));
	notech_reg ififo_rvect3_reg_1(.CP(n_63257), .D(n_36542), .CD(n_62670), .Q
		(ififo_rvect3[1]));
	notech_mux2 i_39078(.S(\nbus_13546[0] ), .A(ififo_rvect3[1]), .B(n_46044
		), .Z(n_36542));
	notech_and4 i_624(.A(n_3153), .B(n_2530), .C(n_2523), .D(n_3151), .Z(n_2527
		));
	notech_reg ififo_rvect3_reg_2(.CP(n_63257), .D(n_36548), .CD(n_62670), .Q
		(ififo_rvect3[2]));
	notech_mux2 i_39086(.S(\nbus_13546[0] ), .A(ififo_rvect3[2]), .B(n_46050
		), .Z(n_36548));
	notech_or2 i_618(.A(n_3123), .B(n_44533), .Z(n_2526));
	notech_reg ififo_rvect3_reg_3(.CP(n_63257), .D(n_36554), .CD(n_62670), .Q
		(ififo_rvect3[3]));
	notech_mux2 i_39094(.S(\nbus_13546[0] ), .A(ififo_rvect3[3]), .B(n_46056
		), .Z(n_36554));
	notech_reg ififo_rvect3_reg_4(.CP(n_63257), .D(n_36560), .CD(n_62665), .Q
		(ififo_rvect3[4]));
	notech_mux2 i_39102(.S(\nbus_13546[0] ), .A(ififo_rvect3[4]), .B(n_46062
		), .Z(n_36560));
	notech_reg ififo_rvect3_reg_5(.CP(n_63257), .D(n_36566), .CD(n_62670), .Q
		(ififo_rvect3[5]));
	notech_mux2 i_39110(.S(\nbus_13546[0] ), .A(ififo_rvect3[5]), .B(n_46068
		), .Z(n_36566));
	notech_or2 i_616(.A(n_3119), .B(n_44562), .Z(n_2523));
	notech_reg ififo_rvect3_reg_6(.CP(n_63257), .D(n_36572), .CD(n_62659), .Q
		(ififo_rvect3[6]));
	notech_mux2 i_39118(.S(\nbus_13546[0] ), .A(ififo_rvect3[6]), .B(n_46074
		), .Z(n_36572));
	notech_or2 i_610(.A(n_3129), .B(n_44548), .Z(n_2522));
	notech_reg ififo_rvect3_reg_7(.CP(n_63257), .D(n_36578), .CD(n_62659), .Q
		(ififo_rvect3[7]));
	notech_mux2 i_39126(.S(\nbus_13546[0] ), .A(ififo_rvect3[7]), .B(n_46080
		), .Z(n_36578));
	notech_reg ififo_rvect2_reg_0(.CP(n_63257), .D(n_36584), .CD(n_62659), .Q
		(ififo_rvect2[0]));
	notech_mux2 i_39134(.S(n_56802), .A(ififo_rvect2[0]), .B(n_48361), .Z(n_36584
		));
	notech_reg ififo_rvect2_reg_1(.CP(n_63257), .D(n_36590), .CD(n_62659), .Q
		(ififo_rvect2[1]));
	notech_mux2 i_39142(.S(n_56802), .A(ififo_rvect2[1]), .B(n_48367), .Z(n_36590
		));
	notech_and4 i_611(.A(n_3148), .B(n_2522), .C(n_2515), .D(n_3146), .Z(n_2519
		));
	notech_reg ififo_rvect2_reg_2(.CP(n_63257), .D(n_36596), .CD(n_62659), .Q
		(ififo_rvect2[2]));
	notech_mux2 i_39150(.S(n_56802), .A(ififo_rvect2[2]), .B(n_48373), .Z(n_36596
		));
	notech_or2 i_605(.A(n_3123), .B(n_44529), .Z(n_2518));
	notech_reg ififo_rvect2_reg_3(.CP(n_63257), .D(n_36602), .CD(n_62659), .Q
		(ififo_rvect2[3]));
	notech_mux2 i_39158(.S(n_56802), .A(ififo_rvect2[3]), .B(n_48379), .Z(n_36602
		));
	notech_reg ififo_rvect2_reg_4(.CP(n_63254), .D(n_36608), .CD(n_62659), .Q
		(ififo_rvect2[4]));
	notech_mux2 i_39166(.S(n_56802), .A(ififo_rvect2[4]), .B(n_48385), .Z(n_36608
		));
	notech_reg ififo_rvect2_reg_5(.CP(n_63254), .D(n_36614), .CD(n_62659), .Q
		(ififo_rvect2[5]));
	notech_mux2 i_39174(.S(n_56802), .A(ififo_rvect2[5]), .B(n_48391), .Z(n_36614
		));
	notech_or2 i_603(.A(n_3119), .B(n_44558), .Z(n_2515));
	notech_reg ififo_rvect2_reg_6(.CP(n_63254), .D(n_36620), .CD(n_62659), .Q
		(ififo_rvect2[6]));
	notech_mux2 i_39182(.S(n_56802), .A(ififo_rvect2[6]), .B(n_48397), .Z(n_36620
		));
	notech_or2 i_597(.A(n_3129), .B(n_44547), .Z(n_2514));
	notech_reg ififo_rvect2_reg_7(.CP(n_63254), .D(n_36626), .CD(n_62659), .Q
		(ififo_rvect2[7]));
	notech_mux2 i_39190(.S(n_56802), .A(ififo_rvect2[7]), .B(n_48403), .Z(n_36626
		));
	notech_reg ififo_rvect1_reg_0(.CP(n_63254), .D(n_36632), .CD(n_62659), .Q
		(ififo_rvect1[0]));
	notech_mux2 i_39198(.S(n_56802), .A(ififo_rvect1[0]), .B(n_44292), .Z(n_36632
		));
	notech_reg ififo_rvect1_reg_1(.CP(n_63254), .D(n_36638), .CD(n_62656), .Q
		(ififo_rvect1[1]));
	notech_mux2 i_39206(.S(n_56802), .A(ififo_rvect1[1]), .B(n_44298), .Z(n_36638
		));
	notech_and4 i_598(.A(n_3143), .B(n_2514), .C(n_2507), .D(n_3141), .Z(n_2511
		));
	notech_reg ififo_rvect1_reg_2(.CP(n_63254), .D(n_36644), .CD(n_62656), .Q
		(ififo_rvect1[2]));
	notech_mux2 i_39214(.S(n_56802), .A(ififo_rvect1[2]), .B(n_44304), .Z(n_36644
		));
	notech_or2 i_592(.A(n_3123), .B(n_44528), .Z(n_2510));
	notech_reg ififo_rvect1_reg_3(.CP(n_63254), .D(n_36650), .CD(n_62656), .Q
		(ififo_rvect1[3]));
	notech_mux2 i_39222(.S(n_56802), .A(ififo_rvect1[3]), .B(n_44310), .Z(n_36650
		));
	notech_reg ififo_rvect1_reg_4(.CP(n_63254), .D(n_36656), .CD(n_62656), .Q
		(ififo_rvect1[4]));
	notech_mux2 i_39230(.S(n_56802), .A(ififo_rvect1[4]), .B(n_44316), .Z(n_36656
		));
	notech_reg ififo_rvect1_reg_5(.CP(n_63254), .D(n_36662), .CD(n_62656), .Q
		(ififo_rvect1[5]));
	notech_mux2 i_39238(.S(n_56802), .A(ififo_rvect1[5]), .B(n_44322), .Z(n_36662
		));
	notech_or2 i_590(.A(n_3119), .B(n_44557), .Z(n_2507));
	notech_reg ififo_rvect1_reg_6(.CP(n_63259), .D(n_36668), .CD(n_62656), .Q
		(ififo_rvect1[6]));
	notech_mux2 i_39246(.S(n_56802), .A(ififo_rvect1[6]), .B(n_44328), .Z(n_36668
		));
	notech_or2 i_584(.A(n_3129), .B(n_44546), .Z(n_2506));
	notech_reg ififo_rvect1_reg_7(.CP(n_63259), .D(n_36674), .CD(n_62659), .Q
		(ififo_rvect1[7]));
	notech_mux2 i_39254(.S(n_56802), .A(ififo_rvect1[7]), .B(n_44334), .Z(n_36674
		));
	notech_reg int_excl_reg_0(.CP(n_63259), .D(n_36680), .CD(n_62656), .Q(int_excl
		[0]));
	notech_mux2 i_39262(.S(\nbus_13566[0] ), .A(int_excl[0]), .B(n_1628100933
		), .Z(n_36680));
	notech_reg int_excl_reg_1(.CP(n_63259), .D(n_36686), .CD(n_62656), .Q(int_excl
		[1]));
	notech_mux2 i_39270(.S(\nbus_13566[0] ), .A(int_excl[1]), .B(n_1629100934
		), .Z(n_36686));
	notech_and4 i_585(.A(n_3138), .B(n_2506), .C(n_2499), .D(n_3136), .Z(n_2503
		));
	notech_reg int_excl_reg_2(.CP(n_63259), .D(n_36692), .CD(n_62656), .Q(int_excl
		[2]));
	notech_mux2 i_39278(.S(\nbus_13566[0] ), .A(int_excl[2]), .B(n_49863), .Z
		(n_36692));
	notech_or2 i_579(.A(n_3123), .B(n_44527), .Z(n_2502));
	notech_reg int_excl_reg_3(.CP(n_63259), .D(n_36698), .CD(n_62661), .Q(int_excl
		[3]));
	notech_mux2 i_39286(.S(\nbus_13566[0] ), .A(int_excl[3]), .B(n_1630100935
		), .Z(n_36698));
	notech_reg int_excl_reg_4(.CP(n_63259), .D(n_36704), .CD(n_62661), .Q(int_excl
		[4]));
	notech_mux2 i_39294(.S(\nbus_13566[0] ), .A(int_excl[4]), .B(n_2844), .Z
		(n_36704));
	notech_reg int_excl_reg_5(.CP(n_63259), .D(n_36710), .CD(n_62661), .Q(int_excl
		[5]));
	notech_mux2 i_39302(.S(\nbus_13566[0] ), .A(int_excl[5]), .B(n_1631100936
		), .Z(n_36710));
	notech_or2 i_577(.A(n_3119), .B(n_44556), .Z(n_2499));
	notech_reg fpu_reg(.CP(n_63259), .D(n_36716), .CD(n_62661), .Q(fpu));
	notech_mux2 i_39310(.S(n_3298), .A(n_1627100932), .B(fpu), .Z(n_36716)
		);
	notech_or2 i_571(.A(n_3129), .B(n_44544), .Z(n_2498));
	notech_reg imm_sz_reg_0(.CP(n_63259), .D(n_36722), .CD(n_62661), .Q(imm_sz
		[0]));
	notech_mux2 i_39318(.S(n_2351), .A(n_41801), .B(imm_sz[0]), .Z(n_36722)
		);
	notech_reg imm_sz_reg_1(.CP(n_63259), .D(n_36728), .CD(n_62661), .Q(imm_sz
		[1]));
	notech_mux2 i_39326(.S(n_2351), .A(n_41807), .B(imm_sz[1]), .Z(n_36728)
		);
	notech_reg imm_sz_reg_2(.CP(n_63257), .D(n_36734), .CD(n_62661), .Q(imm_sz
		[2]));
	notech_mux2 i_39334(.S(n_2351), .A(n_41813), .B(imm_sz[2]), .Z(n_36734)
		);
	notech_and4 i_572(.A(n_3133), .B(n_2498), .C(n_2491), .D(n_3127), .Z(n_2495
		));
	notech_reg i_ptr_reg_0(.CP(n_63257), .D(n_36740), .CD(n_62661), .Q(i_ptr
		[0]));
	notech_mux2 i_39342(.S(n_2388), .A(n_42585), .B(i_ptr[0]), .Z(n_36740)
		);
	notech_or2 i_566(.A(n_3123), .B(n_44525), .Z(n_2494));
	notech_reg i_ptr_reg_1(.CP(n_63257), .D(n_36746), .CD(n_62661), .Q(i_ptr
		[1]));
	notech_mux2 i_39350(.S(n_2388), .A(n_2861), .B(i_ptr[1]), .Z(n_36746));
	notech_reg i_ptr_reg_2(.CP(n_63257), .D(n_36752), .CD(n_62661), .Q(i_ptr
		[2]));
	notech_mux2 i_39358(.S(n_2388), .A(n_2855), .B(i_ptr[2]), .Z(n_36752));
	notech_reg i_ptr_reg_3(.CP(n_63257), .D(n_36761), .CD(n_62661), .Q(i_ptr
		[3]));
	notech_and2 i_39368(.A(n_2388), .B(i_ptr[3]), .Z(n_36761));
	notech_or2 i_564(.A(n_3119), .B(n_44553), .Z(n_2491));
	notech_reg idx_deco_reg_0(.CP(n_63257), .D(n_36764), .CD(n_62659), .Q(idx_deco
		[0]));
	notech_mux2 i_39374(.S(n_3468), .A(n_3574), .B(idx_deco[0]), .Z(n_36764)
		);
	notech_nand2 i_630113(.A(n_44371), .B(n_44372), .Z(n_2490));
	notech_reg idx_deco_reg_1(.CP(n_63259), .D(n_36770), .CD(n_62659), .Q(idx_deco
		[1]));
	notech_mux2 i_39382(.S(n_3468), .A(n_2875), .B(idx_deco[1]), .Z(n_36770)
		);
	notech_nao3 i_561(.A(n_2490), .B(n_3121), .C(n_3117), .Z(n_2489));
	notech_reg fsm_reg_0(.CP(n_63257), .D(n_36776), .CD(n_62659), .Q(fsm[0])
		);
	notech_mux2 i_39390(.S(n_3299), .A(n_42581), .B(fsm[0]), .Z(n_36776));
	notech_nao3 i_559(.A(n_3118), .B(n_44372), .C(imm_sz[1]), .Z(n_2488));
	notech_reg fsm_reg_1(.CP(n_63257), .D(n_36782), .CD(n_62659), .Q(fsm[1])
		);
	notech_mux2 i_39398(.S(n_3299), .A(n_42583), .B(fsm[1]), .Z(n_36782));
	notech_nao3 i_552(.A(n_3060), .B(in128[23]), .C(n_3068), .Z(n_2487));
	notech_reg fsm_reg_2(.CP(n_63257), .D(n_36788), .CD(n_62659), .Q(fsm[2])
		);
	notech_mux2 i_39406(.S(n_3299), .A(n_42584), .B(fsm[2]), .Z(n_36788));
	notech_reg fsm_reg_3(.CP(n_63273), .D(n_36797), .CD(n_62661), .Q(fsm[3])
		);
	notech_and2 i_39416(.A(n_3299), .B(fsm[3]), .Z(n_36797));
	notech_reg fsm_reg_4(.CP(n_63273), .D(n_36803), .CD(n_62661), .Q(fsm[4])
		);
	notech_and2 i_39424(.A(n_3299), .B(fsm[4]), .Z(n_36803));
	notech_and4 i_553(.A(n_3115), .B(n_2487), .C(n_2480), .D(n_3113), .Z(n_2484
		));
	notech_reg repz_reg(.CP(n_63273), .D(n_36806), .CD(n_62659), .Q(repz));
	notech_mux2 i_39430(.S(n_42755), .A(repz), .B(n_1626100931), .Z(n_36806)
		);
	notech_or4 i_544(.A(n_2420), .B(n_2419), .C(n_3064), .D(n_44542), .Z(n_2483
		));
	notech_reg rep_reg(.CP(n_63273), .D(n_36812), .CD(n_62659), .Q(rep));
	notech_mux2 i_39438(.S(n_42755), .A(rep), .B(n_41609), .Z(n_36812));
	notech_reg opz2_reg_0(.CP(n_63273), .D(n_36818), .CD(n_62659), .Q(opz2[0
		]));
	notech_mux2 i_39446(.S(n_56522), .A(opz2[0]), .B(n_1907), .Z(n_36818));
	notech_reg opz2_reg_1(.CP(n_63273), .D(n_36824), .CD(n_62678), .Q(opz2[1
		]));
	notech_mux2 i_39454(.S(n_56522), .A(opz2[1]), .B(n_1902), .Z(n_36824));
	notech_nao3 i_545(.A(n_3057), .B(in128[39]), .C(n_3064), .Z(n_2480));
	notech_reg_set opz2_reg_2(.CP(n_63273), .D(n_36830), .SD(n_62676), .Q(opz2
		[2]));
	notech_mux2 i_39462(.S(n_56522), .A(opz2[2]), .B(n_2892), .Z(n_36830));
	notech_nao3 i_539(.A(n_3060), .B(in128[22]), .C(n_3068), .Z(n_2479));
	notech_reg reps2_reg_0(.CP(n_63273), .D(n_36836), .CD(n_62676), .Q(reps2
		[0]));
	notech_mux2 i_39470(.S(n_56522), .A(reps2[0]), .B(n_1905), .Z(n_36836)
		);
	notech_reg reps2_reg_1(.CP(n_63273), .D(n_36842), .CD(n_62676), .Q(reps2
		[1]));
	notech_mux2 i_39478(.S(n_56527), .A(reps2[1]), .B(n_1909), .Z(n_36842)
		);
	notech_reg reps2_reg_2(.CP(n_63273), .D(n_36848), .CD(n_62676), .Q(reps2
		[2]));
	notech_mux2 i_39486(.S(n_56527), .A(reps2[2]), .B(n_49797), .Z(n_36848)
		);
	notech_and4 i_540(.A(n_3110), .B(n_2479), .C(n_2472), .D(n_3108), .Z(n_2476
		));
	notech_reg reps1_reg_0(.CP(n_63273), .D(n_36854), .CD(n_62676), .Q(reps1
		[0]));
	notech_mux2 i_39494(.S(n_59378), .A(reps1[0]), .B(n_43303), .Z(n_36854)
		);
	notech_or4 i_531(.A(n_2420), .B(n_2419), .C(n_3064), .D(n_44541), .Z(n_2475
		));
	notech_reg reps1_reg_1(.CP(n_63273), .D(n_36860), .CD(n_62676), .Q(reps1
		[1]));
	notech_mux2 i_39502(.S(n_59378), .A(reps1[1]), .B(n_43305), .Z(n_36860)
		);
	notech_reg reps1_reg_2(.CP(n_63273), .D(n_36866), .CD(n_62676), .Q(reps1
		[2]));
	notech_mux2 i_39510(.S(n_59378), .A(reps1[2]), .B(n_42580), .Z(n_36866)
		);
	notech_reg overgs_reg(.CP(n_63273), .D(n_36872), .CD(n_62676), .Q(overgs
		));
	notech_mux2 i_39518(.S(n_3300), .A(n_41609), .B(overgs), .Z(n_36872));
	notech_nao3 i_532(.A(n_3057), .B(in128[38]), .C(n_3064), .Z(n_2472));
	notech_reg over_seg2_reg_5(.CP(n_63270), .D(n_36878), .CD(n_62676), .Q(\over_seg2[5] 
		));
	notech_mux2 i_39526(.S(n_56527), .A(\over_seg2[5] ), .B(n_45639), .Z(n_36878
		));
	notech_nao3 i_526(.A(n_3060), .B(in128[21]), .C(n_3068), .Z(n_2471));
	notech_reg over_seg1_reg_5(.CP(n_63270), .D(n_36884), .CD(n_62676), .Q(\over_seg1[5] 
		));
	notech_mux2 i_39534(.S(n_59378), .A(\over_seg1[5] ), .B(n_42579), .Z(n_36884
		));
	notech_reg to_acu2_reg_0(.CP(n_63273), .D(n_36890), .CD(n_62675), .Q(to_acu2
		[0]));
	notech_mux2 i_39542(.S(n_56522), .A(to_acu2[0]), .B(n_1904), .Z(n_36890)
		);
	notech_reg to_acu2_reg_1(.CP(n_63273), .D(n_36896), .CD(n_62675), .Q(to_acu2
		[1]));
	notech_mux2 i_39550(.S(n_56522), .A(to_acu2[1]), .B(n_1901), .Z(n_36896)
		);
	notech_and4 i_527(.A(n_3105), .B(n_2471), .C(n_2464), .D(n_3103), .Z(n_2468
		));
	notech_reg to_acu2_reg_2(.CP(n_63273), .D(n_36902), .CD(n_62675), .Q(to_acu2
		[2]));
	notech_mux2 i_39558(.S(n_56522), .A(to_acu2[2]), .B(n_1903), .Z(n_36902)
		);
	notech_or4 i_518(.A(n_2420), .B(n_2419), .C(n_3064), .D(n_44540), .Z(n_2467
		));
	notech_reg to_acu2_reg_3(.CP(n_63273), .D(n_36908), .CD(n_62675), .Q(to_acu2
		[3]));
	notech_mux2 i_39566(.S(n_56532), .A(to_acu2[3]), .B(n_1908), .Z(n_36908)
		);
	notech_reg to_acu2_reg_4(.CP(n_63273), .D(n_36914), .CD(n_62675), .Q(to_acu2
		[4]));
	notech_mux2 i_39574(.S(n_56533), .A(to_acu2[4]), .B(n_1906), .Z(n_36914)
		);
	notech_reg to_acu2_reg_5(.CP(n_63275), .D(n_36920), .CD(n_62675), .Q(to_acu2
		[5]));
	notech_mux2 i_39582(.S(n_56533), .A(to_acu2[5]), .B(n_1900), .Z(n_36920)
		);
	notech_nao3 i_519(.A(n_3057), .B(in128[37]), .C(n_3064), .Z(n_2464));
	notech_reg to_acu2_reg_6(.CP(n_63275), .D(n_36926), .CD(n_62675), .Q(to_acu2
		[6]));
	notech_mux2 i_39590(.S(n_56533), .A(to_acu2[6]), .B(n_1910), .Z(n_36926)
		);
	notech_nao3 i_513(.A(n_3060), .B(in128[20]), .C(n_3068), .Z(n_2463));
	notech_reg to_acu2_reg_7(.CP(n_63275), .D(n_36932), .CD(n_62675), .Q(to_acu2
		[7]));
	notech_mux2 i_39598(.S(n_56533), .A(to_acu2[7]), .B(n_3337), .Z(n_36932)
		);
	notech_reg to_acu2_reg_8(.CP(n_63275), .D(n_36938), .CD(n_62675), .Q(to_acu2
		[8]));
	notech_mux2 i_39606(.S(n_56533), .A(to_acu2[8]), .B(n_3335), .Z(n_36938)
		);
	notech_reg to_acu2_reg_9(.CP(n_63275), .D(n_36944), .CD(n_62675), .Q(to_acu2
		[9]));
	notech_mux2 i_39614(.S(n_56533), .A(to_acu2[9]), .B(n_3333), .Z(n_36944)
		);
	notech_and4 i_514(.A(n_3100), .B(n_2463), .C(n_2456), .D(n_3098), .Z(n_2460
		));
	notech_reg to_acu2_reg_10(.CP(n_63275), .D(n_36950), .CD(n_62675), .Q(to_acu2
		[10]));
	notech_mux2 i_39622(.S(n_56533), .A(to_acu2[10]), .B(n_11899519), .Z(n_36950
		));
	notech_or4 i_505(.A(n_2420), .B(n_2419), .C(n_3064), .D(n_44539), .Z(n_2459
		));
	notech_reg to_acu2_reg_11(.CP(n_63275), .D(n_36956), .CD(n_62678), .Q(to_acu2
		[11]));
	notech_mux2 i_39630(.S(n_56533), .A(to_acu2[11]), .B(n_3331), .Z(n_36956
		));
	notech_reg to_acu2_reg_12(.CP(n_63275), .D(n_36962), .CD(n_62678), .Q(to_acu2
		[12]));
	notech_mux2 i_39638(.S(n_56533), .A(to_acu2[12]), .B(n_3329), .Z(n_36962
		));
	notech_reg to_acu2_reg_13(.CP(n_63275), .D(n_36968), .CD(n_62678), .Q(to_acu2
		[13]));
	notech_mux2 i_39646(.S(n_56533), .A(to_acu2[13]), .B(n_3327), .Z(n_36968
		));
	notech_nao3 i_506(.A(n_3057), .B(in128[36]), .C(n_3064), .Z(n_2456));
	notech_reg to_acu2_reg_14(.CP(n_63275), .D(n_36974), .CD(n_62678), .Q(to_acu2
		[14]));
	notech_mux2 i_39654(.S(n_56533), .A(to_acu2[14]), .B(n_3325), .Z(n_36974
		));
	notech_nao3 i_500(.A(n_3060), .B(in128[19]), .C(n_3068), .Z(n_2455));
	notech_reg to_acu2_reg_15(.CP(n_63275), .D(n_36980), .CD(n_62678), .Q(to_acu2
		[15]));
	notech_mux2 i_39662(.S(n_56533), .A(to_acu2[15]), .B(n_3323), .Z(n_36980
		));
	notech_reg to_acu2_reg_16(.CP(n_63275), .D(n_36986), .CD(n_62678), .Q(to_acu2
		[16]));
	notech_mux2 i_39670(.S(n_56533), .A(to_acu2[16]), .B(n_3321), .Z(n_36986
		));
	notech_reg to_acu2_reg_17(.CP(n_63275), .D(n_36992), .CD(n_62678), .Q(to_acu2
		[17]));
	notech_mux2 i_39678(.S(n_56532), .A(to_acu2[17]), .B(n_3319), .Z(n_36992
		));
	notech_and4 i_501(.A(n_3095), .B(n_2455), .C(n_2448), .D(n_3093), .Z(n_2452
		));
	notech_reg to_acu2_reg_18(.CP(n_63275), .D(n_36998), .CD(n_62678), .Q(to_acu2
		[18]));
	notech_mux2 i_39686(.S(n_56532), .A(to_acu2[18]), .B(n_3317), .Z(n_36998
		));
	notech_or4 i_492(.A(n_2420), .B(n_2419), .C(n_3064), .D(n_44538), .Z(n_2451
		));
	notech_reg to_acu2_reg_19(.CP(n_63273), .D(n_37004), .CD(n_62678), .Q(to_acu2
		[19]));
	notech_mux2 i_39694(.S(n_56532), .A(to_acu2[19]), .B(n_73954424), .Z(n_37004
		));
	notech_reg to_acu2_reg_20(.CP(n_63275), .D(n_37010), .CD(n_62678), .Q(to_acu2
		[20]));
	notech_mux2 i_39702(.S(n_56532), .A(to_acu2[20]), .B(n_1521100826), .Z(n_37010
		));
	notech_reg to_acu2_reg_21(.CP(n_63275), .D(n_37016), .CD(n_62678), .Q(to_acu2
		[21]));
	notech_mux2 i_39710(.S(n_56532), .A(to_acu2[21]), .B(n_72154406), .Z(n_37016
		));
	notech_nao3 i_493(.A(n_3057), .B(in128[35]), .C(n_3064), .Z(n_2448));
	notech_reg to_acu2_reg_22(.CP(n_63275), .D(n_37022), .CD(n_62676), .Q(to_acu2
		[22]));
	notech_mux2 i_39718(.S(n_56532), .A(to_acu2[22]), .B(n_72054405), .Z(n_37022
		));
	notech_nao3 i_487(.A(n_3060), .B(in128[18]), .C(n_3068), .Z(n_2447));
	notech_reg to_acu2_reg_23(.CP(n_63275), .D(n_37028), .CD(n_62676), .Q(to_acu2
		[23]));
	notech_mux2 i_39726(.S(n_56532), .A(to_acu2[23]), .B(n_71954404), .Z(n_37028
		));
	notech_reg to_acu2_reg_24(.CP(n_63275), .D(n_37034), .CD(n_62676), .Q(to_acu2
		[24]));
	notech_mux2 i_39734(.S(n_56532), .A(to_acu2[24]), .B(n_73754422), .Z(n_37034
		));
	notech_reg to_acu2_reg_25(.CP(n_63275), .D(n_37040), .CD(n_62676), .Q(to_acu2
		[25]));
	notech_mux2 i_39742(.S(n_56532), .A(to_acu2[25]), .B(n_73654421), .Z(n_37040
		));
	notech_and4 i_488(.A(n_3090), .B(n_2447), .C(n_2440), .D(n_3088), .Z(n_2444
		));
	notech_reg to_acu2_reg_26(.CP(n_63270), .D(n_37046), .CD(n_62676), .Q(to_acu2
		[26]));
	notech_mux2 i_39750(.S(n_56532), .A(to_acu2[26]), .B(n_80654491), .Z(n_37046
		));
	notech_or4 i_479(.A(n_2420), .B(n_2419), .C(n_3064), .D(n_44536), .Z(n_2443
		));
	notech_reg to_acu2_reg_27(.CP(n_63268), .D(n_37052), .CD(n_62676), .Q(to_acu2
		[27]));
	notech_mux2 i_39758(.S(n_56532), .A(to_acu2[27]), .B(n_73554420), .Z(n_37052
		));
	notech_reg to_acu2_reg_28(.CP(n_63268), .D(n_37058), .CD(n_62676), .Q(to_acu2
		[28]));
	notech_mux2 i_39766(.S(n_56532), .A(to_acu2[28]), .B(n_73454419), .Z(n_37058
		));
	notech_reg to_acu2_reg_29(.CP(n_63268), .D(n_37064), .CD(n_62676), .Q(to_acu2
		[29]));
	notech_mux2 i_39774(.S(n_56532), .A(to_acu2[29]), .B(n_1522100827), .Z(n_37064
		));
	notech_nao3 i_480(.A(n_3057), .B(in128[34]), .C(n_3064), .Z(n_2440));
	notech_reg to_acu2_reg_30(.CP(n_63268), .D(n_37070), .CD(n_62676), .Q(to_acu2
		[30]));
	notech_mux2 i_39782(.S(n_56464), .A(to_acu2[30]), .B(n_1523100828), .Z(n_37070
		));
	notech_nao3 i_474(.A(n_3060), .B(in128[17]), .C(n_3068), .Z(n_2439));
	notech_reg to_acu2_reg_31(.CP(n_63268), .D(n_37076), .CD(n_62676), .Q(to_acu2
		[31]));
	notech_mux2 i_39790(.S(n_56464), .A(to_acu2[31]), .B(n_3795), .Z(n_37076
		));
	notech_reg to_acu2_reg_32(.CP(n_63268), .D(n_37082), .CD(n_62671), .Q(to_acu2
		[32]));
	notech_mux2 i_39798(.S(n_56464), .A(to_acu2[32]), .B(n_3793), .Z(n_37082
		));
	notech_reg to_acu2_reg_33(.CP(n_63268), .D(n_37088), .CD(n_62671), .Q(to_acu2
		[33]));
	notech_mux2 i_39806(.S(n_56464), .A(to_acu2[33]), .B(n_3791), .Z(n_37088
		));
	notech_and4 i_475(.A(n_3085), .B(n_2439), .C(n_2432), .D(n_3083), .Z(n_2436
		));
	notech_reg to_acu2_reg_34(.CP(n_63268), .D(n_37094), .CD(n_62671), .Q(to_acu2
		[34]));
	notech_mux2 i_39814(.S(n_56464), .A(to_acu2[34]), .B(n_3789), .Z(n_37094
		));
	notech_or4 i_466(.A(n_2420), .B(n_2419), .C(n_3064), .D(n_44535), .Z(n_2435
		));
	notech_reg to_acu2_reg_35(.CP(n_63268), .D(n_37100), .CD(n_62670), .Q(to_acu2
		[35]));
	notech_mux2 i_39822(.S(n_56464), .A(to_acu2[35]), .B(n_3787), .Z(n_37100
		));
	notech_reg to_acu2_reg_36(.CP(n_63268), .D(n_37106), .CD(n_62670), .Q(to_acu2
		[36]));
	notech_mux2 i_39830(.S(n_56465), .A(to_acu2[36]), .B(n_3785), .Z(n_37106
		));
	notech_reg to_acu2_reg_37(.CP(n_63268), .D(n_37112), .CD(n_62671), .Q(to_acu2
		[37]));
	notech_mux2 i_39838(.S(n_56465), .A(to_acu2[37]), .B(n_3783), .Z(n_37112
		));
	notech_nao3 i_467(.A(n_3057), .B(in128[33]), .C(n_3064), .Z(n_2432));
	notech_reg to_acu2_reg_38(.CP(n_63265), .D(n_37118), .CD(n_62671), .Q(to_acu2
		[38]));
	notech_mux2 i_39846(.S(n_56465), .A(to_acu2[38]), .B(n_3781), .Z(n_37118
		));
	notech_nao3 i_461(.A(n_3060), .B(in128[16]), .C(n_3068), .Z(n_2431));
	notech_reg to_acu2_reg_39(.CP(n_63265), .D(n_37128), .CD(n_62671), .Q(to_acu2
		[39]));
	notech_ao3 i_39858(.A(to_acu2[39]), .B(1'b1), .C(n_56465), .Z(n_37128)
		);
	notech_reg to_acu2_reg_40(.CP(n_63265), .D(n_37130), .CD(n_62671), .Q(to_acu2
		[40]));
	notech_mux2 i_39862(.S(n_56465), .A(to_acu2[40]), .B(n_3779), .Z(n_37130
		));
	notech_reg to_acu2_reg_41(.CP(n_63265), .D(n_37136), .CD(n_62671), .Q(to_acu2
		[41]));
	notech_mux2 i_39870(.S(n_56465), .A(to_acu2[41]), .B(n_65554341), .Z(n_37136
		));
	notech_and4 i_462(.A(n_3080), .B(n_2431), .C(n_2424), .D(n_3074), .Z(n_2428
		));
	notech_reg to_acu2_reg_42(.CP(n_63265), .D(n_37142), .CD(n_62670), .Q(to_acu2
		[42]));
	notech_mux2 i_39878(.S(n_56465), .A(to_acu2[42]), .B(n_3777), .Z(n_37142
		));
	notech_or4 i_453(.A(n_3064), .B(n_2420), .C(n_2419), .D(n_44534), .Z(n_2427
		));
	notech_reg to_acu2_reg_43(.CP(n_63268), .D(n_37148), .CD(n_62670), .Q(to_acu2
		[43]));
	notech_mux2 i_39886(.S(n_56464), .A(to_acu2[43]), .B(n_3775), .Z(n_37148
		));
	notech_reg to_acu2_reg_44(.CP(n_63268), .D(n_37155), .CD(n_62670), .Q(to_acu2
		[44]));
	notech_mux2 i_39894(.S(n_56464), .A(to_acu2[44]), .B(n_3773), .Z(n_37155
		));
	notech_reg to_acu2_reg_45(.CP(n_63268), .D(n_37161), .CD(n_62678), .Q(to_acu2
		[45]));
	notech_mux2 i_39902(.S(n_56464), .A(to_acu2[45]), .B(n_1524100829), .Z(n_37161
		));
	notech_nao3 i_454(.A(n_3057), .B(in128[32]), .C(n_3064), .Z(n_2424));
	notech_reg to_acu2_reg_46(.CP(n_63268), .D(n_37167), .CD(n_62678), .Q(to_acu2
		[46]));
	notech_mux2 i_39910(.S(n_56459), .A(to_acu2[46]), .B(n_3771), .Z(n_37167
		));
	notech_ao3 i_630080(.A(n_44372), .B(n_44371), .C(imm_sz[1]), .Z(n_2423)
		);
	notech_reg to_acu2_reg_47(.CP(n_63268), .D(n_37173), .CD(n_62678), .Q(to_acu2
		[47]));
	notech_mux2 i_39918(.S(n_56464), .A(to_acu2[47]), .B(n_3769), .Z(n_37173
		));
	notech_reg to_acu2_reg_48(.CP(n_63270), .D(n_37179), .CD(n_62670), .Q(to_acu2
		[48]));
	notech_mux2 i_39926(.S(n_56464), .A(to_acu2[48]), .B(n_3767), .Z(n_37179
		));
	notech_reg to_acu2_reg_49(.CP(n_63270), .D(n_37185), .CD(n_62670), .Q(to_acu2
		[49]));
	notech_mux2 i_39934(.S(n_56464), .A(to_acu2[49]), .B(n_3765), .Z(n_37185
		));
	notech_nor2 i_441(.A(displc[0]), .B(n_3056), .Z(n_2420));
	notech_reg to_acu2_reg_50(.CP(n_63270), .D(n_37191), .CD(n_62670), .Q(to_acu2
		[50]));
	notech_mux2 i_39942(.S(n_56464), .A(to_acu2[50]), .B(n_3763), .Z(n_37191
		));
	notech_and2 i_440(.A(displc[0]), .B(n_3056), .Z(n_2419));
	notech_reg to_acu2_reg_51(.CP(n_63270), .D(n_37197), .CD(n_62670), .Q(to_acu2
		[51]));
	notech_mux2 i_39950(.S(n_56464), .A(to_acu2[51]), .B(n_3761), .Z(n_37197
		));
	notech_ao3 i_437(.A(displc[1]), .B(n_44163), .C(displc[2]), .Z(n_2418)
		);
	notech_reg to_acu2_reg_52(.CP(n_63270), .D(n_37203), .CD(n_62670), .Q(to_acu2
		[52]));
	notech_mux2 i_39958(.S(n_56464), .A(to_acu2[52]), .B(n_3759), .Z(n_37203
		));
	notech_and2 i_436(.A(displc[2]), .B(n_3059), .Z(n_2417));
	notech_reg to_acu2_reg_53(.CP(n_63270), .D(n_37209), .CD(n_62675), .Q(to_acu2
		[53]));
	notech_mux2 i_39966(.S(n_56464), .A(to_acu2[53]), .B(n_3757), .Z(n_37209
		));
	notech_and2 i_432(.A(n_44731), .B(n_44730), .Z(n_2416));
	notech_reg to_acu2_reg_54(.CP(n_63270), .D(n_37215), .CD(n_62675), .Q(to_acu2
		[54]));
	notech_mux2 i_39974(.S(n_56464), .A(to_acu2[54]), .B(n_1899), .Z(n_37215
		));
	notech_reg to_acu2_reg_55(.CP(n_63270), .D(n_37221), .CD(n_62675), .Q(to_acu2
		[55]));
	notech_mux2 i_39982(.S(n_56464), .A(to_acu2[55]), .B(n_3755), .Z(n_37221
		));
	notech_reg to_acu2_reg_56(.CP(n_63270), .D(n_37227), .CD(n_62671), .Q(to_acu2
		[56]));
	notech_mux2 i_39990(.S(n_56465), .A(to_acu2[56]), .B(n_3753), .Z(n_37227
		));
	notech_and4 i_320(.A(n_44526), .B(\to_acu2_0[7] ), .C(in128[16]), .D(in128
		[18]), .Z(n_2413));
	notech_reg to_acu2_reg_57(.CP(n_63270), .D(n_37233), .CD(n_62675), .Q(to_acu2
		[57]));
	notech_mux2 i_39998(.S(n_56448), .A(to_acu2[57]), .B(n_3751), .Z(n_37233
		));
	notech_ao3 i_313(.A(\fpu_modrm[0] ), .B(n_3052), .C(\fpu_modrm[1] ), .Z(n_2412
		));
	notech_reg to_acu2_reg_58(.CP(n_63270), .D(n_37239), .CD(n_62675), .Q(to_acu2
		[58]));
	notech_mux2 i_40006(.S(n_56448), .A(to_acu2[58]), .B(n_3749), .Z(n_37239
		));
	notech_and4 i_311(.A(n_2408), .B(n_3046), .C(n_2407), .D(twobyte), .Z(n_2411
		));
	notech_reg to_acu2_reg_59(.CP(n_63268), .D(n_37245), .CD(n_62675), .Q(to_acu2
		[59]));
	notech_mux2 i_40014(.S(n_56448), .A(to_acu2[59]), .B(n_3747), .Z(n_37245
		));
	notech_nand3 i_65795(.A(n_2405), .B(n_3041), .C(n_2403), .Z(n_2410));
	notech_reg to_acu2_reg_60(.CP(n_63270), .D(n_37251), .CD(n_62675), .Q(to_acu2
		[60]));
	notech_mux2 i_40022(.S(n_56448), .A(to_acu2[60]), .B(n_3745), .Z(n_37251
		));
	notech_and2 i_310(.A(n_44745), .B(n_2410), .Z(n_2409));
	notech_reg to_acu2_reg_61(.CP(n_63268), .D(n_37257), .CD(n_62675), .Q(to_acu2
		[61]));
	notech_mux2 i_40030(.S(n_56448), .A(to_acu2[61]), .B(n_3743), .Z(n_37257
		));
	notech_nand2 i_303(.A(n_2406), .B(\to_acu2_0[26] ), .Z(n_2408));
	notech_reg to_acu2_reg_62(.CP(n_63268), .D(n_37263), .CD(n_62675), .Q(to_acu2
		[62]));
	notech_mux2 i_40038(.S(n_56448), .A(to_acu2[62]), .B(n_3741), .Z(n_37263
		));
	notech_nand3 i_305(.A(\to_acu2_0[21] ), .B(\to_acu2_0[23] ), .C(\to_acu2_0[22] 
		), .Z(n_2407));
	notech_reg to_acu2_reg_63(.CP(n_63268), .D(n_37269), .CD(n_62671), .Q(to_acu2
		[63]));
	notech_mux2 i_40046(.S(n_56448), .A(to_acu2[63]), .B(n_3739), .Z(n_37269
		));
	notech_nand2 i_304(.A(n_44746), .B(n_44717), .Z(n_2406));
	notech_reg to_acu2_reg_64(.CP(n_63270), .D(n_37275), .CD(n_62671), .Q(to_acu2
		[64]));
	notech_mux2 i_40054(.S(n_56475), .A(to_acu2[64]), .B(n_3737), .Z(n_37275
		));
	notech_nand2 i_294(.A(\to_acu2_0[17] ), .B(\to_acu2_0[18] ), .Z(n_2405)
		);
	notech_reg to_acu2_reg_65(.CP(n_63270), .D(n_37281), .CD(n_62671), .Q(to_acu2
		[65]));
	notech_mux2 i_40062(.S(n_56475), .A(to_acu2[65]), .B(n_3735), .Z(n_37281
		));
	notech_nand2 i_296(.A(n_44712), .B(n_44711), .Z(n_2404));
	notech_reg to_acu2_reg_66(.CP(n_63270), .D(n_37287), .CD(n_62671), .Q(to_acu2
		[66]));
	notech_mux2 i_40070(.S(n_56475), .A(to_acu2[66]), .B(n_3733), .Z(n_37287
		));
	notech_nand2 i_295(.A(n_2404), .B(\to_acu2_0[13] ), .Z(n_2403));
	notech_reg to_acu2_reg_67(.CP(n_63270), .D(n_37293), .CD(n_62671), .Q(to_acu2
		[67]));
	notech_mux2 i_40078(.S(n_56448), .A(to_acu2[67]), .B(n_3731), .Z(n_37293
		));
	notech_nao3 i_44(.A(n_60854), .B(n_44744), .C(n_2975), .Z(n_2402));
	notech_reg to_acu2_reg_68(.CP(n_63270), .D(n_37299), .CD(n_62671), .Q(to_acu2
		[68]));
	notech_mux2 i_40086(.S(n_56448), .A(to_acu2[68]), .B(n_3729), .Z(n_37299
		));
	notech_ao3 i_6258(.A(n_2399), .B(n_3037), .C(n_3029), .Z(n_2401));
	notech_reg to_acu2_reg_69(.CP(n_63238), .D(n_37305), .CD(n_62671), .Q(to_acu2
		[69]));
	notech_mux2 i_40094(.S(n_56475), .A(to_acu2[69]), .B(n_3727), .Z(n_37305
		));
	notech_reg to_acu2_reg_70(.CP(n_63238), .D(n_37311), .CD(n_62671), .Q(to_acu2
		[70]));
	notech_mux2 i_40102(.S(n_56465), .A(to_acu2[70]), .B(n_3725), .Z(n_37311
		));
	notech_or4 i_269(.A(ififo_rvect1[1]), .B(ififo_rvect1[0]), .C(n_3033), .D
		(n_3032), .Z(n_2399));
	notech_reg to_acu2_reg_71(.CP(n_63238), .D(n_37317), .CD(n_62671), .Q(to_acu2
		[71]));
	notech_mux2 i_40110(.S(n_56465), .A(to_acu2[71]), .B(n_3723), .Z(n_37317
		));
	notech_ao4 i_254(.A(n_60248), .B(n_3027), .C(pc_req), .D(n_2393), .Z(n_2398
		));
	notech_reg to_acu2_reg_72(.CP(n_63238), .D(n_37323), .CD(n_62671), .Q(to_acu2
		[72]));
	notech_mux2 i_40118(.S(n_56465), .A(to_acu2[72]), .B(n_3721), .Z(n_37323
		));
	notech_reg to_acu2_reg_73(.CP(n_63238), .D(n_37329), .CD(n_62671), .Q(to_acu2
		[73]));
	notech_mux2 i_40126(.S(n_56465), .A(to_acu2[73]), .B(n_3719), .Z(n_37329
		));
	notech_reg to_acu2_reg_74(.CP(n_63241), .D(n_37335), .CD(n_62656), .Q(to_acu2
		[74]));
	notech_mux2 i_40134(.S(n_56465), .A(to_acu2[74]), .B(n_3717), .Z(n_37335
		));
	notech_nao3 i_3230218(.A(n_2376), .B(n_2335), .C(valid_len[5]), .Z(n_2395
		));
	notech_reg to_acu2_reg_75(.CP(n_63241), .D(n_37341), .CD(n_62640), .Q(to_acu2
		[75]));
	notech_mux2 i_40142(.S(n_56465), .A(to_acu2[75]), .B(n_3715), .Z(n_37341
		));
	notech_reg to_acu2_reg_76(.CP(n_63241), .D(n_37347), .CD(n_62640), .Q(to_acu2
		[76]));
	notech_mux2 i_40150(.S(n_56465), .A(to_acu2[76]), .B(n_3713), .Z(n_37347
		));
	notech_mux2 i_251(.S(n_5405), .A(n_230099379), .B(n_2391), .Z(n_2393));
	notech_reg to_acu2_reg_77(.CP(n_63238), .D(n_37353), .CD(n_62640), .Q(to_acu2
		[77]));
	notech_mux2 i_40158(.S(n_56448), .A(to_acu2[77]), .B(n_3711), .Z(n_37353
		));
	notech_reg to_acu2_reg_78(.CP(n_63241), .D(n_37359), .CD(n_62640), .Q(to_acu2
		[78]));
	notech_mux2 i_40166(.S(n_56448), .A(to_acu2[78]), .B(n_3709), .Z(n_37359
		));
	notech_ao3 i_65854(.A(fsm[0]), .B(fsm[1]), .C(n_2970), .Z(n_2391));
	notech_reg to_acu2_reg_79(.CP(n_63238), .D(n_37365), .CD(n_62640), .Q(to_acu2
		[79]));
	notech_mux2 i_40174(.S(n_56448), .A(to_acu2[79]), .B(n_3707), .Z(n_37365
		));
	notech_reg to_acu2_reg_80(.CP(n_63238), .D(n_37371), .CD(n_62643), .Q(to_acu2
		[80]));
	notech_mux2 i_40182(.S(n_56465), .A(to_acu2[80]), .B(n_3705), .Z(n_37371
		));
	notech_reg to_acu2_reg_81(.CP(n_63238), .D(n_37377), .CD(n_62643), .Q(to_acu2
		[81]));
	notech_mux2 i_40190(.S(n_56465), .A(to_acu2[81]), .B(n_3703), .Z(n_37377
		));
	notech_and4 i_70795(.A(n_60127), .B(n_2386), .C(n_3022), .D(n_2387), .Z(n_2388
		));
	notech_reg to_acu2_reg_82(.CP(n_63238), .D(n_37383), .CD(n_62643), .Q(to_acu2
		[82]));
	notech_mux2 i_40198(.S(n_56465), .A(to_acu2[82]), .B(n_3701), .Z(n_37383
		));
	notech_nao3 i_2289(.A(n_60921), .B(n_60854), .C(pg_fault), .Z(n_2387));
	notech_reg to_acu2_reg_83(.CP(n_63238), .D(n_37389), .CD(n_62640), .Q(to_acu2
		[83]));
	notech_mux2 i_40206(.S(n_56453), .A(to_acu2[83]), .B(n_3699), .Z(n_37389
		));
	notech_nand3 i_2744(.A(n_2379), .B(fpu), .C(n_2337), .Z(n_2386));
	notech_reg to_acu2_reg_84(.CP(n_63238), .D(n_37395), .CD(n_62643), .Q(to_acu2
		[84]));
	notech_mux2 i_40214(.S(n_56453), .A(to_acu2[84]), .B(n_47596), .Z(n_37395
		));
	notech_nand2 i_245(.A(n_3020), .B(n_2379), .Z(n_2385));
	notech_reg to_acu2_reg_85(.CP(n_63238), .D(n_37401), .CD(n_62640), .Q(to_acu2
		[85]));
	notech_mux2 i_40222(.S(n_56453), .A(to_acu2[85]), .B(n_3697), .Z(n_37401
		));
	notech_nao3 i_244(.A(n_60859), .B(n_44744), .C(n_3017), .Z(n_2384));
	notech_reg to_acu2_reg_86(.CP(n_63238), .D(n_37407), .CD(n_62640), .Q(to_acu2
		[86]));
	notech_mux2 i_40230(.S(n_56453), .A(to_acu2[86]), .B(n_3695), .Z(n_37407
		));
	notech_nand2 i_68(.A(n_1676), .B(n_44165), .Z(n_2383));
	notech_reg to_acu2_reg_87(.CP(n_63238), .D(n_37413), .CD(n_62640), .Q(to_acu2
		[87]));
	notech_mux2 i_40238(.S(n_56453), .A(to_acu2[87]), .B(n_3693), .Z(n_37413
		));
	notech_nand2 i_188(.A(n_42724), .B(n_2975), .Z(n_2382));
	notech_reg to_acu2_reg_88(.CP(n_63238), .D(n_37419), .CD(n_62640), .Q(to_acu2
		[88]));
	notech_mux2 i_40246(.S(n_56453), .A(to_acu2[88]), .B(n_3691), .Z(n_37419
		));
	notech_nand2 i_117(.A(n_2379), .B(fpu), .Z(n_2381));
	notech_reg to_acu2_reg_89(.CP(n_63238), .D(n_37425), .CD(n_62640), .Q(to_acu2
		[89]));
	notech_mux2 i_40254(.S(n_56453), .A(to_acu2[89]), .B(n_3689), .Z(n_37425
		));
	notech_or4 i_175(.A(\to_acu2_0[9] ), .B(\to_acu2_0[10] ), .C(\to_acu2_0[11] 
		), .D(\to_acu2_0[8] ), .Z(n_2380));
	notech_reg to_acu2_reg_90(.CP(n_63241), .D(n_37431), .CD(n_62640), .Q(to_acu2
		[90]));
	notech_mux2 i_40262(.S(n_56453), .A(to_acu2[90]), .B(n_3687), .Z(n_37431
		));
	notech_and4 i_28(.A(n_2378), .B(n_2999), .C(n_2395), .D(n_2996), .Z(n_2379
		));
	notech_reg to_acu2_reg_91(.CP(n_63241), .D(n_37437), .CD(n_62640), .Q(to_acu2
		[91]));
	notech_mux2 i_40270(.S(n_56453), .A(to_acu2[91]), .B(n_3685), .Z(n_37437
		));
	notech_or4 i_16(.A(valid_len[5]), .B(valid_len[4]), .C(n_2989), .D(n_2377
		), .Z(n_2378));
	notech_reg to_acu2_reg_92(.CP(n_63241), .D(n_37443), .CD(n_62640), .Q(to_acu2
		[92]));
	notech_mux2 i_40278(.S(n_56454), .A(to_acu2[92]), .B(n_3683), .Z(n_37443
		));
	notech_and2 i_167(.A(valid_len[1]), .B(valid_len[0]), .Z(n_2377));
	notech_reg to_acu2_reg_93(.CP(n_63241), .D(n_37449), .CD(n_62640), .Q(to_acu2
		[93]));
	notech_mux2 i_40286(.S(n_56453), .A(to_acu2[93]), .B(n_3681), .Z(n_37449
		));
	notech_nand2 i_162(.A(n_2980), .B(valid_len[4]), .Z(n_2376));
	notech_reg to_acu2_reg_94(.CP(n_63241), .D(n_37455), .CD(n_62640), .Q(to_acu2
		[94]));
	notech_mux2 i_40294(.S(n_56453), .A(to_acu2[94]), .B(n_3679), .Z(n_37455
		));
	notech_or2 i_156(.A(n_2981), .B(n_2367), .Z(n_2375));
	notech_reg to_acu2_reg_95(.CP(n_63243), .D(n_37461), .CD(n_62640), .Q(to_acu2
		[95]));
	notech_mux2 i_40302(.S(n_56453), .A(to_acu2[95]), .B(n_3677), .Z(n_37461
		));
	notech_reg to_acu2_reg_96(.CP(n_63243), .D(n_37467), .CD(n_62643), .Q(to_acu2
		[96]));
	notech_mux2 i_40310(.S(n_56448), .A(to_acu2[96]), .B(n_3675), .Z(n_37467
		));
	notech_reg to_acu2_reg_97(.CP(n_63243), .D(n_37473), .CD(n_62643), .Q(to_acu2
		[97]));
	notech_mux2 i_40318(.S(n_56448), .A(to_acu2[97]), .B(n_3673), .Z(n_37473
		));
	notech_and2 i_151(.A(valid_len[2]), .B(n_44186), .Z(n_2372));
	notech_reg to_acu2_reg_98(.CP(n_63243), .D(n_37479), .CD(n_62643), .Q(to_acu2
		[98]));
	notech_mux2 i_40326(.S(n_56453), .A(to_acu2[98]), .B(n_3671), .Z(n_37479
		));
	notech_and2 i_9(.A(valid_len[1]), .B(n_44185), .Z(n_2371));
	notech_reg to_acu2_reg_99(.CP(n_63243), .D(n_37485), .CD(n_62643), .Q(to_acu2
		[99]));
	notech_mux2 i_40334(.S(n_56448), .A(to_acu2[99]), .B(n_1525100830), .Z(n_37485
		));
	notech_ao3 i_2775(.A(valid_len[0]), .B(n_2357), .C(n_2358), .Z(n_2370)
		);
	notech_reg to_acu2_reg_100(.CP(n_63241), .D(n_37491), .CD(n_62643), .Q(to_acu2
		[100]));
	notech_mux2 i_40342(.S(n_56448), .A(to_acu2[100]), .B(n_81454499), .Z(n_37491
		));
	notech_and2 i_26(.A(n_2981), .B(valid_len[3]), .Z(n_2369));
	notech_reg to_acu2_reg_101(.CP(n_63241), .D(n_37497), .CD(n_62645), .Q(to_acu2
		[101]));
	notech_mux2 i_40350(.S(n_56448), .A(to_acu2[101]), .B(n_77554460), .Z(n_37497
		));
	notech_or4 i_157(.A(n_2371), .B(n_2370), .C(n_2372), .D(n_2369), .Z(n_2368
		));
	notech_reg to_acu2_reg_102(.CP(n_63241), .D(n_37503), .CD(n_62645), .Q(to_acu2
		[102]));
	notech_mux2 i_40358(.S(n_56453), .A(to_acu2[102]), .B(n_79554480), .Z(n_37503
		));
	notech_and2 i_152(.A(valid_len[3]), .B(n_2366), .Z(n_2367));
	notech_reg to_acu2_reg_103(.CP(n_63241), .D(n_37509), .CD(n_62645), .Q(to_acu2
		[103]));
	notech_mux2 i_40366(.S(n_56453), .A(to_acu2[103]), .B(n_76854453), .Z(n_37509
		));
	notech_or2 i_153(.A(valid_len[2]), .B(n_44186), .Z(n_2366));
	notech_reg to_acu2_reg_104(.CP(n_63241), .D(n_37515), .CD(n_62645), .Q(to_acu2
		[104]));
	notech_mux2 i_40374(.S(n_56453), .A(to_acu2[104]), .B(n_81654501), .Z(n_37515
		));
	notech_reg to_acu2_reg_105(.CP(n_63241), .D(n_37521), .CD(n_62645), .Q(to_acu2
		[105]));
	notech_mux2 i_40382(.S(n_56453), .A(to_acu2[105]), .B(n_81754502), .Z(n_37521
		));
	notech_reg to_acu2_reg_106(.CP(n_63241), .D(n_37527), .CD(n_62643), .Q(to_acu2
		[106]));
	notech_mux2 i_40390(.S(n_56453), .A(to_acu2[106]), .B(n_80554490), .Z(n_37527
		));
	notech_reg to_acu2_reg_107(.CP(n_63241), .D(n_37533), .CD(n_62643), .Q(to_acu2
		[107]));
	notech_mux2 i_40398(.S(n_56453), .A(to_acu2[107]), .B(n_79154476), .Z(n_37533
		));
	notech_and2 i_143(.A(n_44372), .B(n_43428), .Z(n_2362));
	notech_reg to_acu2_reg_108(.CP(n_63241), .D(n_37539), .CD(n_62643), .Q(to_acu2
		[108]));
	notech_mux2 i_40406(.S(n_56453), .A(to_acu2[108]), .B(n_1526100831), .Z(n_37539
		));
	notech_reg to_acu2_reg_109(.CP(n_63241), .D(n_37545), .CD(n_62643), .Q(to_acu2
		[109]));
	notech_mux2 i_40414(.S(n_56454), .A(to_acu2[109]), .B(n_77454459), .Z(n_37545
		));
	notech_reg to_acu2_reg_110(.CP(n_63241), .D(n_37551), .CD(n_62643), .Q(to_acu2
		[110]));
	notech_mux2 i_40422(.S(n_56459), .A(to_acu2[110]), .B(n_1527100832), .Z(n_37551
		));
	notech_reg to_acu2_reg_111(.CP(n_63238), .D(n_37557), .CD(n_62643), .Q(to_acu2
		[111]));
	notech_mux2 i_40430(.S(n_56459), .A(to_acu2[111]), .B(n_74154426), .Z(n_37557
		));
	notech_xor2 i_6240(.A(imm_sz[0]), .B(i_ptr[0]), .Z(n_2358));
	notech_reg to_acu2_reg_112(.CP(n_63233), .D(n_37563), .CD(n_62643), .Q(to_acu2
		[112]));
	notech_mux2 i_40438(.S(n_56459), .A(to_acu2[112]), .B(n_82654511), .Z(n_37563
		));
	notech_or2 i_138(.A(valid_len[1]), .B(n_44185), .Z(n_2357));
	notech_reg to_acu2_reg_113(.CP(n_63233), .D(n_37569), .CD(n_62643), .Q(to_acu2
		[113]));
	notech_mux2 i_40446(.S(n_56454), .A(to_acu2[113]), .B(n_82354508), .Z(n_37569
		));
	notech_reg to_acu2_reg_114(.CP(n_63233), .D(n_37575), .CD(n_62643), .Q(to_acu2
		[114]));
	notech_mux2 i_40454(.S(n_56454), .A(to_acu2[114]), .B(n_76354448), .Z(n_37575
		));
	notech_reg to_acu2_reg_115(.CP(n_63233), .D(n_37581), .CD(n_62643), .Q(to_acu2
		[115]));
	notech_mux2 i_40462(.S(n_56459), .A(to_acu2[115]), .B(n_74954434), .Z(n_37581
		));
	notech_reg to_acu2_reg_116(.CP(n_63233), .D(n_37587), .CD(n_62643), .Q(to_acu2
		[116]));
	notech_mux2 i_40470(.S(n_56459), .A(to_acu2[116]), .B(n_82954514), .Z(n_37587
		));
	notech_reg to_acu2_reg_117(.CP(n_63233), .D(n_37593), .CD(n_62635), .Q(to_acu2
		[117]));
	notech_mux2 i_40478(.S(n_56459), .A(to_acu2[117]), .B(n_74854433), .Z(n_37593
		));
	notech_and2 i_133(.A(imm_sz[1]), .B(i_ptr[1]), .Z(n_2352));
	notech_reg to_acu2_reg_118(.CP(n_63236), .D(n_37599), .CD(n_62635), .Q(to_acu2
		[118]));
	notech_mux2 i_40486(.S(n_56459), .A(to_acu2[118]), .B(n_75854443), .Z(n_37599
		));
	notech_and2 i_70886(.A(n_5765), .B(n_2349), .Z(n_2351));
	notech_reg to_acu2_reg_119(.CP(n_63233), .D(n_37605), .CD(n_62635), .Q(to_acu2
		[119]));
	notech_mux2 i_40494(.S(n_56459), .A(to_acu2[119]), .B(n_75354438), .Z(n_37605
		));
	notech_and4 i_126(.A(n_2960), .B(n_2342), .C(n_2341), .D(n_2348), .Z(n_2350
		));
	notech_reg to_acu2_reg_120(.CP(n_63233), .D(n_37611), .CD(n_62635), .Q(to_acu2
		[120]));
	notech_mux2 i_40502(.S(n_56459), .A(to_acu2[120]), .B(n_83054515), .Z(n_37611
		));
	notech_or2 i_127(.A(n_44164), .B(n_2350), .Z(n_2349));
	notech_reg to_acu2_reg_121(.CP(n_63233), .D(n_37617), .CD(n_62635), .Q(to_acu2
		[121]));
	notech_mux2 i_40510(.S(n_56459), .A(to_acu2[121]), .B(n_82254507), .Z(n_37617
		));
	notech_nand2 i_125(.A(n_1744), .B(n_2957), .Z(n_2348));
	notech_reg to_acu2_reg_122(.CP(n_63233), .D(n_37623), .CD(n_62638), .Q(to_acu2
		[122]));
	notech_mux2 i_40518(.S(n_56459), .A(to_acu2[122]), .B(n_76554450), .Z(n_37623
		));
	notech_and4 i_115(.A(n_44685), .B(n_44680), .C(n_44681), .D(n_1878), .Z(n_2347
		));
	notech_reg to_acu2_reg_123(.CP(n_63233), .D(n_37629), .CD(n_62638), .Q(to_acu2
		[123]));
	notech_mux2 i_40526(.S(n_56454), .A(to_acu2[123]), .B(n_74454429), .Z(n_37629
		));
	notech_reg to_acu2_reg_124(.CP(n_63233), .D(n_37635), .CD(n_62635), .Q(to_acu2
		[124]));
	notech_mux2 i_40534(.S(n_56454), .A(to_acu2[124]), .B(n_1528100833), .Z(n_37635
		));
	notech_and2 i_107(.A(n_44718), .B(n_44679), .Z(n_2345));
	notech_reg to_acu2_reg_125(.CP(n_63233), .D(n_37641), .CD(n_62635), .Q(to_acu2
		[125]));
	notech_mux2 i_40542(.S(n_56454), .A(to_acu2[125]), .B(n_75654441), .Z(n_37641
		));
	notech_reg to_acu2_reg_126(.CP(n_63233), .D(n_37647), .CD(n_62635), .Q(to_acu2
		[126]));
	notech_mux2 i_40550(.S(n_56454), .A(to_acu2[126]), .B(n_75254437), .Z(n_37647
		));
	notech_nand2 i_100(.A(n_44707), .B(n_44706), .Z(n_2343));
	notech_reg to_acu2_reg_127(.CP(n_63233), .D(n_37653), .CD(n_62635), .Q(to_acu2
		[127]));
	notech_mux2 i_40558(.S(n_56454), .A(to_acu2[127]), .B(n_76454449), .Z(n_37653
		));
	notech_nand3 i_103(.A(n_44718), .B(twobyte), .C(n_2343), .Z(n_2342));
	notech_reg to_acu2_reg_128(.CP(n_63233), .D(n_37659), .CD(n_62635), .Q(to_acu2
		[128]));
	notech_mux2 i_40566(.S(n_56454), .A(to_acu2[128]), .B(n_65354339), .Z(n_37659
		));
	notech_nand2 i_102(.A(n_44745), .B(n_2956), .Z(n_2341));
	notech_reg to_acu2_reg_129(.CP(n_63233), .D(n_37665), .CD(n_62635), .Q(to_acu2
		[129]));
	notech_mux2 i_40574(.S(n_56454), .A(to_acu2[129]), .B(n_81954504), .Z(n_37665
		));
	notech_nand2 i_57(.A(\to_acu2_0[5] ), .B(\to_acu2_0[48] ), .Z(n_2340));
	notech_reg to_acu2_reg_130(.CP(n_63233), .D(n_37671), .CD(n_62635), .Q(to_acu2
		[130]));
	notech_mux2 i_40582(.S(n_56454), .A(to_acu2[130]), .B(n_77354458), .Z(n_37671
		));
	notech_nand2 i_49(.A(n_1879), .B(n_44685), .Z(n_2339));
	notech_reg to_acu2_reg_131(.CP(n_63233), .D(n_37677), .CD(n_62635), .Q(to_acu2
		[131]));
	notech_mux2 i_40590(.S(n_56454), .A(to_acu2[131]), .B(n_74554430), .Z(n_37677
		));
	notech_nand2 i_38(.A(\to_acu2_0[5] ), .B(\to_acu2_0[59] ), .Z(n_2338));
	notech_reg to_acu2_reg_132(.CP(n_63233), .D(n_37683), .CD(n_62635), .Q(to_acu2
		[132]));
	notech_mux2 i_40598(.S(n_56454), .A(to_acu2[132]), .B(n_64954335), .Z(n_37683
		));
	notech_nao3 i_71370(.A(n_1733), .B(n_44751), .C(db67), .Z(n_2337));
	notech_reg to_acu2_reg_133(.CP(n_63236), .D(n_37689), .CD(n_62635), .Q(to_acu2
		[133]));
	notech_mux2 i_40606(.S(n_56454), .A(to_acu2[133]), .B(n_75454439), .Z(n_37689
		));
	notech_nand2 i_6229(.A(idx_deco[1]), .B(idx_deco[0]), .Z(n_2336));
	notech_reg to_acu2_reg_134(.CP(n_63236), .D(n_37695), .CD(n_62635), .Q(to_acu2
		[134]));
	notech_mux2 i_40614(.S(n_56454), .A(to_acu2[134]), .B(n_75754442), .Z(n_37695
		));
	notech_nand3 i_2769(.A(n_2990), .B(n_2375), .C(n_2368), .Z(n_2335));
	notech_reg to_acu2_reg_135(.CP(n_63236), .D(n_37701), .CD(n_62635), .Q(to_acu2
		[135]));
	notech_mux2 i_40622(.S(n_56454), .A(to_acu2[135]), .B(n_78354468), .Z(n_37701
		));
	notech_reg to_acu2_reg_136(.CP(n_63236), .D(n_37707), .CD(n_62635), .Q(to_acu2
		[136]));
	notech_mux2 i_40630(.S(n_56475), .A(to_acu2[136]), .B(n_65154337), .Z(n_37707
		));
	notech_reg to_acu2_reg_137(.CP(n_63236), .D(n_37713), .CD(n_62635), .Q(to_acu2
		[137]));
	notech_mux2 i_40638(.S(n_56488), .A(to_acu2[137]), .B(n_81854503), .Z(n_37713
		));
	notech_reg to_acu2_reg_138(.CP(n_63238), .D(n_37719), .CD(n_62638), .Q(to_acu2
		[138]));
	notech_mux2 i_40646(.S(n_56488), .A(to_acu2[138]), .B(n_77154456), .Z(n_37719
		));
	notech_reg to_acu2_reg_139(.CP(n_63238), .D(n_37725), .CD(n_62638), .Q(to_acu2
		[139]));
	notech_mux2 i_40654(.S(n_56488), .A(to_acu2[139]), .B(n_76254447), .Z(n_37725
		));
	notech_reg to_acu2_reg_140(.CP(n_63236), .D(n_37731), .CD(n_62638), .Q(to_acu2
		[140]));
	notech_mux2 i_40662(.S(n_56488), .A(to_acu2[140]), .B(n_65454340), .Z(n_37731
		));
	notech_ao4 i_104078014(.A(n_44545), .B(n_3162), .C(n_3163), .D(n_44602),
		 .Z(n_2329));
	notech_reg to_acu2_reg_141(.CP(n_63236), .D(n_37737), .CD(n_62638), .Q(to_acu2
		[141]));
	notech_mux2 i_40670(.S(n_56488), .A(to_acu2[141]), .B(n_78454469), .Z(n_37737
		));
	notech_reg to_acu2_reg_142(.CP(n_63236), .D(n_37743), .CD(n_62638), .Q(to_acu2
		[142]));
	notech_mux2 i_40678(.S(n_56488), .A(to_acu2[142]), .B(n_76154446), .Z(n_37743
		));
	notech_reg to_acu2_reg_143(.CP(n_63236), .D(n_37749), .CD(n_62640), .Q(to_acu2
		[143]));
	notech_mux2 i_40686(.S(n_56488), .A(to_acu2[143]), .B(n_76054445), .Z(n_37749
		));
	notech_ao4 i_104278012(.A(n_3198), .B(n_44554), .C(n_3155), .D(n_44564),
		 .Z(n_2326));
	notech_reg to_acu2_reg_144(.CP(n_63236), .D(n_37755), .CD(n_62640), .Q(to_acu2
		[144]));
	notech_mux2 i_40694(.S(n_56488), .A(to_acu2[144]), .B(n_82454509), .Z(n_37755
		));
	notech_ao4 i_104378011(.A(n_3157), .B(n_44593), .C(n_3156), .D(n_44574),
		 .Z(n_2325));
	notech_reg to_acu2_reg_145(.CP(n_63236), .D(n_37761), .CD(n_62640), .Q(to_acu2
		[145]));
	notech_mux2 i_40702(.S(n_56488), .A(to_acu2[145]), .B(n_82154506), .Z(n_37761
		));
	notech_ao4 i_104478010(.A(n_3162), .B(n_44540), .C(n_3163), .D(n_44598),
		 .Z(n_2324));
	notech_reg to_acu2_reg_146(.CP(n_63236), .D(n_37767), .CD(n_62638), .Q(to_acu2
		[146]));
	notech_mux2 i_40710(.S(n_56488), .A(to_acu2[146]), .B(n_75954444), .Z(n_37767
		));
	notech_reg to_acu2_reg_147(.CP(n_63236), .D(n_37773), .CD(n_62638), .Q(to_acu2
		[147]));
	notech_mux2 i_40718(.S(n_56488), .A(to_acu2[147]), .B(n_77254457), .Z(n_37773
		));
	notech_reg to_acu2_reg_148(.CP(n_63236), .D(n_37779), .CD(n_62638), .Q(to_acu2
		[148]));
	notech_mux2 i_40726(.S(n_56488), .A(to_acu2[148]), .B(n_82754512), .Z(n_37779
		));
	notech_ao4 i_104678008(.A(n_3158), .B(n_44550), .C(n_3155), .D(n_44559),
		 .Z(n_232199400));
	notech_reg to_acu2_reg_149(.CP(n_63236), .D(n_37785), .CD(n_62638), .Q(to_acu2
		[149]));
	notech_mux2 i_40734(.S(n_56488), .A(to_acu2[149]), .B(n_79354478), .Z(n_37785
		));
	notech_ao4 i_104778007(.A(n_3157), .B(n_44588), .C(n_3156), .D(n_44569),
		 .Z(n_232099399));
	notech_reg to_acu2_reg_150(.CP(n_63236), .D(n_37791), .CD(n_62638), .Q(to_acu2
		[150]));
	notech_mux2 i_40742(.S(n_56487), .A(to_acu2[150]), .B(n_79254477), .Z(n_37791
		));
	notech_reg to_acu2_reg_151(.CP(n_63236), .D(n_37797), .CD(n_62638), .Q(to_acu2
		[151]));
	notech_mux2 i_40750(.S(n_56487), .A(to_acu2[151]), .B(n_74354428), .Z(n_37797
		));
	notech_ao4 i_104878006(.A(n_44551), .B(n_3129), .C(n_44580), .D(n_3130),
		 .Z(n_231899397));
	notech_reg to_acu2_reg_152(.CP(n_63236), .D(n_37803), .CD(n_62638), .Q(to_acu2
		[152]));
	notech_mux2 i_40758(.S(n_56487), .A(to_acu2[152]), .B(n_65254338), .Z(n_37803
		));
	notech_reg to_acu2_reg_153(.CP(n_63236), .D(n_37809), .CD(n_62638), .Q(to_acu2
		[153]));
	notech_mux2 i_40766(.S(n_56487), .A(to_acu2[153]), .B(n_82054505), .Z(n_37809
		));
	notech_ao4 i_105078004(.A(n_3124), .B(n_44589), .C(n_44560), .D(n_3119),
		 .Z(n_231699395));
	notech_reg to_acu2_reg_154(.CP(n_63252), .D(n_37815), .CD(n_62638), .Q(to_acu2
		[154]));
	notech_mux2 i_40774(.S(n_56487), .A(to_acu2[154]), .B(n_77754462), .Z(n_37815
		));
	notech_ao4 i_105178003(.A(n_3125), .B(n_44570), .C(n_3123), .D(n_44532),
		 .Z(n_231599394));
	notech_reg to_acu2_reg_155(.CP(n_63252), .D(n_37821), .CD(n_62638), .Q(to_acu2
		[155]));
	notech_mux2 i_40782(.S(n_56487), .A(to_acu2[155]), .B(n_78054465), .Z(n_37821
		));
	notech_reg to_acu2_reg_156(.CP(n_63252), .D(n_37827), .CD(n_62638), .Q(to_acu2
		[156]));
	notech_mux2 i_40790(.S(n_56487), .A(to_acu2[156]), .B(n_64854334), .Z(n_37827
		));
	notech_ao4 i_105378001(.A(n_3130), .B(n_44578), .C(n_3125), .D(n_44569),
		 .Z(n_231399392));
	notech_reg to_acu2_reg_157(.CP(n_63249), .D(n_37833), .CD(n_62638), .Q(to_acu2
		[157]));
	notech_mux2 i_40798(.S(n_56488), .A(to_acu2[157]), .B(n_75154436), .Z(n_37833
		));
	notech_reg to_acu2_reg_158(.CP(n_63252), .D(n_37839), .CD(n_62638), .Q(to_acu2
		[158]));
	notech_mux2 i_40806(.S(n_56488), .A(to_acu2[158]), .B(n_79954484), .Z(n_37839
		));
	notech_ao4 i_105577999(.A(n_3124), .B(n_44588), .C(n_3119), .D(n_44559),
		 .Z(n_231199390));
	notech_reg to_acu2_reg_159(.CP(n_63252), .D(n_37845), .CD(n_62645), .Q(to_acu2
		[159]));
	notech_mux2 i_40814(.S(n_56488), .A(to_acu2[159]), .B(n_75554440), .Z(n_37845
		));
	notech_ao4 i_105677998(.A(n_3129), .B(n_44550), .C(n_44530), .D(n_3123),
		 .Z(n_231099389));
	notech_reg to_acu2_reg_160(.CP(n_63252), .D(n_37851), .CD(n_62654), .Q(to_acu2
		[160]));
	notech_mux2 i_40822(.S(n_56487), .A(to_acu2[160]), .B(n_82554510), .Z(n_37851
		));
	notech_reg to_acu2_reg_161(.CP(n_63252), .D(n_37857), .CD(n_62654), .Q(to_acu2
		[161]));
	notech_mux2 i_40830(.S(n_56488), .A(to_acu2[161]), .B(n_76754452), .Z(n_37857
		));
	notech_ao4 i_105877996(.A(n_3124), .B(n_44583), .C(n_3130), .D(n_44574),
		 .Z(n_230899387));
	notech_reg to_acu2_reg_162(.CP(n_63252), .D(n_37863), .CD(n_62654), .Q(to_acu2
		[162]));
	notech_mux2 i_40838(.S(n_56488), .A(to_acu2[162]), .B(n_80054485), .Z(n_37863
		));
	notech_reg to_acu2_reg_163(.CP(n_63252), .D(n_37869), .CD(n_62651), .Q(to_acu2
		[163]));
	notech_mux2 i_40846(.S(n_56493), .A(to_acu2[163]), .B(n_80154486), .Z(n_37869
		));
	notech_ao4 i_106077994(.A(n_44564), .B(n_3125), .C(n_3119), .D(n_44554),
		 .Z(n_230699385));
	notech_reg to_acu2_reg_164(.CP(n_63249), .D(n_37875), .CD(n_62654), .Q(to_acu2
		[164]));
	notech_mux2 i_40854(.S(n_56498), .A(to_acu2[164]), .B(n_82854513), .Z(n_37875
		));
	notech_ao4 i_106177993(.A(n_3132), .B(n_44535), .C(n_3123), .D(n_44526),
		 .Z(n_230599384));
	notech_reg to_acu2_reg_165(.CP(n_63249), .D(n_37881), .CD(n_62654), .Q(to_acu2
		[165]));
	notech_mux2 i_40862(.S(n_56498), .A(to_acu2[165]), .B(n_81254497), .Z(n_37881
		));
	notech_reg to_acu2_reg_166(.CP(n_63249), .D(n_37887), .CD(n_62654), .Q(to_acu2
		[166]));
	notech_mux2 i_40870(.S(n_56498), .A(to_acu2[166]), .B(n_80954494), .Z(n_37887
		));
	notech_ao4 i_106777987(.A(n_225799336), .B(n_5767), .C(n_194199020), .D(n_225699335
		), .Z(n_230399382));
	notech_reg to_acu2_reg_167(.CP(n_63249), .D(n_37893), .CD(n_62654), .Q(to_acu2
		[167]));
	notech_mux2 i_40878(.S(n_56498), .A(to_acu2[167]), .B(n_80254487), .Z(n_37893
		));
	notech_and2 i_2779014(.A(n_1669), .B(n_3026), .Z(n_230299381));
	notech_reg to_acu2_reg_168(.CP(n_63249), .D(n_37899), .CD(n_62654), .Q(to_acu2
		[168]));
	notech_mux2 i_40886(.S(n_56498), .A(to_acu2[168]), .B(n_78654471), .Z(n_37899
		));
	notech_reg to_acu2_reg_169(.CP(n_63249), .D(n_37905), .CD(n_62654), .Q(to_acu2
		[169]));
	notech_mux2 i_40894(.S(n_56498), .A(to_acu2[169]), .B(n_80354488), .Z(n_37905
		));
	notech_and2 i_3379008(.A(n_1669), .B(n_2336), .Z(n_230099379));
	notech_reg to_acu2_reg_170(.CP(n_63249), .D(n_37911), .CD(n_62651), .Q(to_acu2
		[170]));
	notech_mux2 i_40902(.S(n_56498), .A(to_acu2[170]), .B(n_78754472), .Z(n_37911
		));
	notech_and2 i_1879023(.A(n_42724), .B(n_194099019), .Z(n_229999378));
	notech_reg to_acu2_reg_171(.CP(n_63249), .D(n_37917), .CD(n_62651), .Q(to_acu2
		[171]));
	notech_mux2 i_40910(.S(n_56498), .A(to_acu2[171]), .B(n_67454360), .Z(n_37917
		));
	notech_reg to_acu2_reg_172(.CP(n_63249), .D(n_37923), .CD(n_62651), .Q(to_acu2
		[172]));
	notech_mux2 i_40918(.S(n_56498), .A(to_acu2[172]), .B(n_67554361), .Z(n_37923
		));
	notech_reg to_acu2_reg_173(.CP(n_63249), .D(n_37929), .CD(n_62651), .Q(to_acu2
		[173]));
	notech_mux2 i_40926(.S(n_56498), .A(to_acu2[173]), .B(n_67654362), .Z(n_37929
		));
	notech_or2 i_79478255(.A(n_42549), .B(n_1912), .Z(n_229699375));
	notech_reg to_acu2_reg_174(.CP(n_63249), .D(n_37935), .CD(n_62651), .Q(to_acu2
		[174]));
	notech_mux2 i_40934(.S(n_56498), .A(to_acu2[174]), .B(n_67854363), .Z(n_37935
		));
	notech_reg to_acu2_reg_175(.CP(n_63254), .D(n_37941), .CD(n_62651), .Q(to_acu2
		[175]));
	notech_mux2 i_40942(.S(n_56498), .A(to_acu2[175]), .B(n_67954364), .Z(n_37941
		));
	notech_reg to_acu2_reg_176(.CP(n_63254), .D(n_37947), .CD(n_62651), .Q(to_acu2
		[176]));
	notech_mux2 i_40950(.S(n_56498), .A(to_acu2[176]), .B(n_3469), .Z(n_37947
		));
	notech_reg to_acu2_reg_177(.CP(n_63254), .D(n_37953), .CD(n_62651), .Q(to_acu2
		[177]));
	notech_mux2 i_40958(.S(n_56493), .A(to_acu2[177]), .B(n_68054365), .Z(n_37953
		));
	notech_reg to_acu2_reg_178(.CP(n_63254), .D(n_37959), .CD(n_62651), .Q(to_acu2
		[178]));
	notech_mux2 i_40966(.S(n_56493), .A(to_acu2[178]), .B(n_3313), .Z(n_37959
		));
	notech_reg to_acu2_reg_179(.CP(n_63254), .D(n_37965), .CD(n_62651), .Q(to_acu2
		[179]));
	notech_mux2 i_40974(.S(n_56493), .A(to_acu2[179]), .B(n_3311), .Z(n_37965
		));
	notech_or2 i_2479017(.A(n_3129), .B(n_44545), .Z(n_229199370));
	notech_reg to_acu2_reg_180(.CP(n_63254), .D(n_37971), .CD(n_62651), .Q(to_acu2
		[180]));
	notech_mux2 i_40982(.S(n_56493), .A(to_acu2[180]), .B(n_3309), .Z(n_37971
		));
	notech_reg to_acu2_reg_181(.CP(n_63254), .D(n_37977), .CD(n_62656), .Q(to_acu2
		[181]));
	notech_mux2 i_40990(.S(n_56493), .A(to_acu2[181]), .B(n_3307), .Z(n_37977
		));
	notech_reg to_acu2_reg_182(.CP(n_63254), .D(n_37983), .CD(n_62656), .Q(to_acu2
		[182]));
	notech_mux2 i_40998(.S(n_56493), .A(to_acu2[182]), .B(n_3305), .Z(n_37983
		));
	notech_reg to_acu2_reg_183(.CP(n_63254), .D(n_37989), .CD(n_62656), .Q(to_acu2
		[183]));
	notech_mux2 i_41006(.S(n_56493), .A(to_acu2[183]), .B(n_68154366), .Z(n_37989
		));
	notech_reg to_acu2_reg_184(.CP(n_63254), .D(n_37995), .CD(n_62656), .Q(to_acu2
		[184]));
	notech_mux2 i_41014(.S(n_56493), .A(to_acu2[184]), .B(n_68254367), .Z(n_37995
		));
	notech_reg to_acu2_reg_185(.CP(n_63252), .D(n_38001), .CD(n_62656), .Q(to_acu2
		[185]));
	notech_mux2 i_41022(.S(n_56498), .A(to_acu2[185]), .B(n_68354368), .Z(n_38001
		));
	notech_reg to_acu2_reg_186(.CP(n_63252), .D(n_38007), .CD(n_62656), .Q(to_acu2
		[186]));
	notech_mux2 i_41030(.S(n_56498), .A(to_acu2[186]), .B(n_68454369), .Z(n_38007
		));
	notech_or2 i_2579016(.A(n_3132), .B(n_44540), .Z(n_228499363));
	notech_reg to_acu2_reg_187(.CP(n_63252), .D(n_38013), .CD(n_62656), .Q(to_acu2
		[187]));
	notech_mux2 i_41038(.S(n_56493), .A(to_acu2[187]), .B(n_68554370), .Z(n_38013
		));
	notech_reg to_acu2_reg_188(.CP(n_63252), .D(n_38019), .CD(n_62656), .Q(to_acu2
		[188]));
	notech_mux2 i_41046(.S(n_56493), .A(to_acu2[188]), .B(n_68654371), .Z(n_38019
		));
	notech_reg to_acu2_reg_189(.CP(n_63252), .D(n_38025), .CD(n_62656), .Q(to_acu2
		[189]));
	notech_mux2 i_41054(.S(n_56493), .A(to_acu2[189]), .B(n_68754372), .Z(n_38025
		));
	notech_reg to_acu2_reg_190(.CP(n_63252), .D(n_38031), .CD(n_62656), .Q(to_acu2
		[190]));
	notech_mux2 i_41062(.S(n_56476), .A(to_acu2[190]), .B(n_1529100834), .Z(n_38031
		));
	notech_reg to_acu2_reg_191(.CP(n_63252), .D(n_38037), .CD(n_62654), .Q(to_acu2
		[191]));
	notech_mux2 i_41070(.S(n_56476), .A(to_acu2[191]), .B(n_1530100835), .Z(n_38037
		));
	notech_reg to_acu2_reg_192(.CP(n_63252), .D(n_38043), .CD(n_62654), .Q(to_acu2
		[192]));
	notech_mux2 i_41078(.S(n_56476), .A(to_acu2[192]), .B(n_1531100836), .Z(n_38043
		));
	notech_reg to_acu2_reg_193(.CP(n_63252), .D(n_38049), .CD(n_62654), .Q(to_acu2
		[193]));
	notech_mux2 i_41086(.S(n_56476), .A(to_acu2[193]), .B(n_69154376), .Z(n_38049
		));
	notech_or2 i_2679015(.A(n_3132), .B(n_44541), .Z(n_227799356));
	notech_reg to_acu2_reg_194(.CP(n_63252), .D(n_38055), .CD(n_62654), .Q(to_acu2
		[194]));
	notech_mux2 i_41094(.S(n_56476), .A(to_acu2[194]), .B(n_3604), .Z(n_38055
		));
	notech_reg to_acu2_reg_195(.CP(n_63252), .D(n_38061), .CD(n_62654), .Q(to_acu2
		[195]));
	notech_mux2 i_41102(.S(n_56476), .A(to_acu2[195]), .B(n_3602), .Z(n_38061
		));
	notech_reg to_acu2_reg_196(.CP(n_63249), .D(n_38067), .CD(n_62654), .Q(to_acu2
		[196]));
	notech_mux2 i_41110(.S(n_56476), .A(to_acu2[196]), .B(n_3600), .Z(n_38067
		));
	notech_reg to_acu2_reg_197(.CP(n_63243), .D(n_38073), .CD(n_62654), .Q(to_acu2
		[197]));
	notech_mux2 i_41118(.S(n_56476), .A(to_acu2[197]), .B(n_3598), .Z(n_38073
		));
	notech_reg to_acu2_reg_198(.CP(n_63247), .D(n_38079), .CD(n_62654), .Q(to_acu2
		[198]));
	notech_mux2 i_41126(.S(n_56476), .A(to_acu2[198]), .B(n_3596), .Z(n_38079
		));
	notech_reg to_acu2_reg_199(.CP(n_63243), .D(n_38085), .CD(n_62654), .Q(to_acu2
		[199]));
	notech_mux2 i_41134(.S(n_56476), .A(to_acu2[199]), .B(n_3594), .Z(n_38085
		));
	notech_reg to_acu2_reg_200(.CP(n_63243), .D(n_38091), .CD(n_62654), .Q(to_acu2
		[200]));
	notech_mux2 i_41142(.S(n_56476), .A(to_acu2[200]), .B(n_3592), .Z(n_38091
		));
	notech_or2 i_1679025(.A(n_3164), .B(n_44578), .Z(n_227099349));
	notech_reg to_acu2_reg_201(.CP(n_63243), .D(n_38097), .CD(n_62654), .Q(to_acu2
		[201]));
	notech_mux2 i_41150(.S(n_56476), .A(to_acu2[201]), .B(n_3590), .Z(n_38097
		));
	notech_reg to_acu2_reg_202(.CP(n_63247), .D(n_38103), .CD(n_62649), .Q(to_acu2
		[202]));
	notech_mux2 i_41158(.S(n_56476), .A(to_acu2[202]), .B(n_3588), .Z(n_38103
		));
	notech_reg to_acu2_reg_203(.CP(n_63247), .D(n_38109), .CD(n_62649), .Q(to_acu2
		[203]));
	notech_mux2 i_41166(.S(n_56475), .A(to_acu2[203]), .B(n_3586), .Z(n_38109
		));
	notech_reg to_acu2_reg_204(.CP(n_63247), .D(n_38115), .CD(n_62645), .Q(to_acu2
		[204]));
	notech_mux2 i_41174(.S(n_56475), .A(to_acu2[204]), .B(n_3584), .Z(n_38115
		));
	notech_reg to_acu2_reg_205(.CP(n_63247), .D(n_38121), .CD(n_62645), .Q(to_acu2
		[205]));
	notech_mux2 i_41182(.S(n_56475), .A(to_acu2[205]), .B(n_3582), .Z(n_38121
		));
	notech_reg to_acu2_reg_206(.CP(n_63247), .D(n_38127), .CD(n_62645), .Q(to_acu2
		[206]));
	notech_mux2 i_41190(.S(n_56475), .A(to_acu2[206]), .B(n_3580), .Z(n_38127
		));
	notech_reg to_acu2_reg_207(.CP(n_63243), .D(n_38133), .CD(n_62649), .Q(to_acu2
		[207]));
	notech_mux2 i_41198(.S(n_56475), .A(to_acu2[207]), .B(n_1532100837), .Z(n_38133
		));
	notech_or2 i_1779024(.A(n_3164), .B(n_44583), .Z(n_226399342));
	notech_reg to_acu2_reg_208(.CP(n_63243), .D(n_38139), .CD(n_62649), .Q(to_acu2
		[208]));
	notech_mux2 i_41206(.S(n_56475), .A(to_acu2[208]), .B(n_3578), .Z(n_38139
		));
	notech_reg to_acu2_reg_209(.CP(n_63243), .D(n_38145), .CD(n_62649), .Q(to_acu2
		[209]));
	notech_mux2 i_41214(.S(n_56475), .A(to_acu2[209]), .B(n_1533100838), .Z(n_38145
		));
	notech_reg to_acu2_reg_210(.CP(n_63243), .D(n_38151), .CD(n_62649), .Q(to_acu2
		[210]));
	notech_mux2 i_41222(.S(n_56475), .A(to_acu2[210]), .B(n_48352), .Z(n_38151
		));
	notech_or4 i_61678433(.A(n_60367), .B(pc_req), .C(pg_fault), .D(n_230299381
		), .Z(n_226099339));
	notech_reg to_acu1_reg_0(.CP(n_63243), .D(n_38157), .CD(n_62649), .Q(to_acu1
		[0]));
	notech_mux2 i_41230(.S(n_59383), .A(to_acu1[0]), .B(n_43709), .Z(n_38157
		));
	notech_nao3 i_61578434(.A(idx_deco[1]), .B(n_43431), .C(n_59153), .Z(n_225999338
		));
	notech_reg to_acu1_reg_1(.CP(n_63243), .D(n_38163), .CD(n_62645), .Q(to_acu1
		[1]));
	notech_mux2 i_41238(.S(n_59383), .A(to_acu1[1]), .B(n_43711), .Z(n_38163
		));
	notech_and3 i_2962(.A(n_60921), .B(lenpc2[10]), .C(n_60859), .Z(n_44118)
		);
	notech_reg to_acu1_reg_2(.CP(n_63243), .D(n_38169), .CD(n_62645), .Q(to_acu1
		[2]));
	notech_mux2 i_41246(.S(n_59383), .A(to_acu1[2]), .B(n_43713), .Z(n_38169
		));
	notech_and3 i_2959(.A(n_60921), .B(lenpc2[7]), .C(n_60859), .Z(n_44100)
		);
	notech_reg to_acu1_reg_3(.CP(n_63243), .D(n_38175), .CD(n_62645), .Q(to_acu1
		[3]));
	notech_mux2 i_41254(.S(n_59378), .A(to_acu1[3]), .B(n_43716), .Z(n_38175
		));
	notech_reg to_acu1_reg_4(.CP(n_63243), .D(n_38181), .CD(n_62645), .Q(to_acu1
		[4]));
	notech_mux2 i_41262(.S(n_59378), .A(to_acu1[4]), .B(n_43718), .Z(n_38181
		));
	notech_ao3 i_22578824(.A(n_1669), .B(n_3026), .C(n_5405), .Z(n_225799336
		));
	notech_reg to_acu1_reg_5(.CP(n_63243), .D(n_38187), .CD(n_62645), .Q(to_acu1
		[5]));
	notech_mux2 i_41270(.S(n_59378), .A(to_acu1[5]), .B(n_43721), .Z(n_38187
		));
	notech_ao3 i_3479007(.A(n_2336), .B(n_1669), .C(n_5405), .Z(n_225699335)
		);
	notech_reg to_acu1_reg_6(.CP(n_63243), .D(n_38193), .CD(n_62645), .Q(to_acu1
		[6]));
	notech_mux2 i_41278(.S(n_59388), .A(to_acu1[6]), .B(n_43723), .Z(n_38193
		));
	notech_and4 i_79078259(.A(n_230899387), .B(n_230699385), .C(n_230599384)
		, .D(n_229199370), .Z(n_225599334));
	notech_reg to_acu1_reg_7(.CP(n_63249), .D(n_38199), .CD(n_62645), .Q(to_acu1
		[7]));
	notech_mux2 i_41286(.S(n_59389), .A(to_acu1[7]), .B(n_43725), .Z(n_38199
		));
	notech_and4 i_78978260(.A(n_231399392), .B(n_231199390), .C(n_231099389)
		, .D(n_228499363), .Z(n_225499333));
	notech_reg to_acu1_reg_8(.CP(n_63249), .D(n_38205), .CD(n_62645), .Q(to_acu1
		[8]));
	notech_mux2 i_41294(.S(n_59389), .A(to_acu1[8]), .B(n_43728), .Z(n_38205
		));
	notech_and4 i_78878261(.A(n_231899397), .B(n_231699395), .C(n_231599394)
		, .D(n_227799356), .Z(n_225399332));
	notech_reg to_acu1_reg_9(.CP(n_63247), .D(n_38211), .CD(n_62645), .Q(to_acu1
		[9]));
	notech_mux2 i_41302(.S(n_59389), .A(to_acu1[9]), .B(n_43730), .Z(n_38211
		));
	notech_and4 i_78378266(.A(n_232199400), .B(n_232099399), .C(n_2324), .D(n_227099349
		), .Z(n_225299331));
	notech_reg to_acu1_reg_10(.CP(n_63247), .D(n_38217), .CD(n_62645), .Q(to_acu1
		[10]));
	notech_mux2 i_41310(.S(n_59389), .A(to_acu1[10]), .B(n_43843), .Z(n_38217
		));
	notech_and4 i_77878271(.A(n_2326), .B(n_2325), .C(n_2329), .D(n_226399342
		), .Z(n_225199330));
	notech_reg to_acu1_reg_11(.CP(n_63247), .D(n_38223), .CD(n_62645), .Q(to_acu1
		[11]));
	notech_mux2 i_41318(.S(n_59389), .A(to_acu1[11]), .B(n_43733), .Z(n_38223
		));
	notech_reg to_acu1_reg_12(.CP(n_63249), .D(n_38229), .CD(n_62651), .Q(to_acu1
		[12]));
	notech_mux2 i_41326(.S(n_59389), .A(to_acu1[12]), .B(n_43735), .Z(n_38229
		));
	notech_reg to_acu1_reg_13(.CP(n_63249), .D(n_38235), .CD(n_62651), .Q(to_acu1
		[13]));
	notech_mux2 i_41334(.S(n_59389), .A(to_acu1[13]), .B(n_43737), .Z(n_38235
		));
	notech_reg to_acu1_reg_14(.CP(n_63249), .D(n_38241), .CD(n_62651), .Q(to_acu1
		[14]));
	notech_mux2 i_41342(.S(n_59389), .A(to_acu1[14]), .B(n_43740), .Z(n_38241
		));
	notech_reg to_acu1_reg_15(.CP(n_63249), .D(n_38247), .CD(n_62649), .Q(to_acu1
		[15]));
	notech_mux2 i_41350(.S(n_59389), .A(to_acu1[15]), .B(n_43742), .Z(n_38247
		));
	notech_reg to_acu1_reg_16(.CP(n_63249), .D(n_38253), .CD(n_62649), .Q(to_acu1
		[16]));
	notech_mux2 i_41358(.S(n_59389), .A(to_acu1[16]), .B(n_43745), .Z(n_38253
		));
	notech_reg to_acu1_reg_17(.CP(n_63247), .D(n_38259), .CD(n_62651), .Q(to_acu1
		[17]));
	notech_mux2 i_41366(.S(n_59389), .A(to_acu1[17]), .B(n_43747), .Z(n_38259
		));
	notech_reg to_acu1_reg_18(.CP(n_63247), .D(n_38265), .CD(n_62651), .Q(to_acu1
		[18]));
	notech_mux2 i_41374(.S(n_59389), .A(to_acu1[18]), .B(n_43749), .Z(n_38265
		));
	notech_reg to_acu1_reg_19(.CP(n_63247), .D(n_38271), .CD(n_62651), .Q(to_acu1
		[19]));
	notech_mux2 i_41382(.S(n_59389), .A(to_acu1[19]), .B(n_43862), .Z(n_38271
		));
	notech_reg to_acu1_reg_20(.CP(n_63247), .D(n_38277), .CD(n_62651), .Q(to_acu1
		[20]));
	notech_mux2 i_41390(.S(n_59388), .A(to_acu1[20]), .B(n_43865), .Z(n_38277
		));
	notech_reg to_acu1_reg_21(.CP(n_63247), .D(n_38283), .CD(n_62651), .Q(to_acu1
		[21]));
	notech_mux2 i_41398(.S(n_59388), .A(to_acu1[21]), .B(n_43867), .Z(n_38283
		));
	notech_reg to_acu1_reg_22(.CP(n_63247), .D(n_38289), .CD(n_62649), .Q(to_acu1
		[22]));
	notech_mux2 i_41406(.S(n_59388), .A(to_acu1[22]), .B(n_43869), .Z(n_38289
		));
	notech_reg to_acu1_reg_23(.CP(n_63247), .D(n_38295), .CD(n_62649), .Q(to_acu1
		[23]));
	notech_mux2 i_41414(.S(n_59388), .A(to_acu1[23]), .B(n_43872), .Z(n_38295
		));
	notech_reg to_acu1_reg_24(.CP(n_63247), .D(n_38301), .CD(n_62649), .Q(to_acu1
		[24]));
	notech_mux2 i_41422(.S(n_59388), .A(to_acu1[24]), .B(n_43874), .Z(n_38301
		));
	notech_reg to_acu1_reg_25(.CP(n_63247), .D(n_38307), .CD(n_62649), .Q(to_acu1
		[25]));
	notech_mux2 i_41430(.S(n_59388), .A(to_acu1[25]), .B(n_43877), .Z(n_38307
		));
	notech_reg to_acu1_reg_26(.CP(n_63247), .D(n_38313), .CD(n_62649), .Q(to_acu1
		[26]));
	notech_mux2 i_41438(.S(n_59388), .A(to_acu1[26]), .B(n_43880), .Z(n_38313
		));
	notech_reg to_acu1_reg_27(.CP(n_63247), .D(n_38319), .CD(n_62649), .Q(to_acu1
		[27]));
	notech_mux2 i_41446(.S(n_59388), .A(to_acu1[27]), .B(n_43883), .Z(n_38319
		));
	notech_reg to_acu1_reg_28(.CP(n_63184), .D(n_38325), .CD(n_62649), .Q(to_acu1
		[28]));
	notech_mux2 i_41454(.S(n_59388), .A(to_acu1[28]), .B(n_43885), .Z(n_38325
		));
	notech_reg to_acu1_reg_29(.CP(n_63117), .D(n_38331), .CD(n_62649), .Q(to_acu1
		[29]));
	notech_mux2 i_41462(.S(n_59388), .A(to_acu1[29]), .B(n_43889), .Z(n_38331
		));
	notech_reg to_acu1_reg_30(.CP(n_63117), .D(n_38337), .CD(n_62649), .Q(to_acu1
		[30]));
	notech_mux2 i_41470(.S(n_59388), .A(to_acu1[30]), .B(n_43891), .Z(n_38337
		));
	notech_reg to_acu1_reg_31(.CP(n_63117), .D(n_38343), .CD(n_62649), .Q(to_acu1
		[31]));
	notech_mux2 i_41478(.S(n_59388), .A(to_acu1[31]), .B(n_42903), .Z(n_38343
		));
	notech_reg to_acu1_reg_32(.CP(n_63117), .D(n_38349), .CD(n_62649), .Q(to_acu1
		[32]));
	notech_mux2 i_41486(.S(n_59388), .A(to_acu1[32]), .B(n_42907), .Z(n_38349
		));
	notech_reg to_acu1_reg_33(.CP(n_63117), .D(n_38355), .CD(n_62586), .Q(to_acu1
		[33]));
	notech_mux2 i_41494(.S(n_59320), .A(to_acu1[33]), .B(n_42911), .Z(n_38355
		));
	notech_reg to_acu1_reg_34(.CP(n_63117), .D(n_38361), .CD(n_62519), .Q(to_acu1
		[34]));
	notech_mux2 i_41502(.S(n_59320), .A(to_acu1[34]), .B(n_42914), .Z(n_38361
		));
	notech_reg to_acu1_reg_35(.CP(n_63117), .D(n_38367), .CD(n_62519), .Q(to_acu1
		[35]));
	notech_mux2 i_41510(.S(n_59320), .A(to_acu1[35]), .B(n_42917), .Z(n_38367
		));
	notech_reg to_acu1_reg_36(.CP(n_63117), .D(n_38373), .CD(n_62519), .Q(to_acu1
		[36]));
	notech_mux2 i_41518(.S(n_59320), .A(to_acu1[36]), .B(n_42919), .Z(n_38373
		));
	notech_reg to_acu1_reg_37(.CP(n_63117), .D(n_38379), .CD(n_62519), .Q(to_acu1
		[37]));
	notech_mux2 i_41526(.S(n_59320), .A(to_acu1[37]), .B(n_42921), .Z(n_38379
		));
	notech_reg to_acu1_reg_38(.CP(n_63117), .D(n_38385), .CD(n_62519), .Q(to_acu1
		[38]));
	notech_mux2 i_41534(.S(n_59320), .A(to_acu1[38]), .B(n_42924), .Z(n_38385
		));
	notech_reg to_acu1_reg_39(.CP(n_63117), .D(n_38391), .CD(n_62519), .Q(to_acu1
		[39]));
	notech_mux2 i_41542(.S(n_59321), .A(to_acu1[39]), .B(n_1196100504), .Z(n_38391
		));
	notech_reg to_acu1_reg_40(.CP(n_63117), .D(n_38397), .CD(n_62519), .Q(to_acu1
		[40]));
	notech_mux2 i_41550(.S(n_59321), .A(to_acu1[40]), .B(n_42926), .Z(n_38397
		));
	notech_reg to_acu1_reg_41(.CP(n_63117), .D(n_38403), .CD(n_62519), .Q(to_acu1
		[41]));
	notech_mux2 i_41558(.S(n_59321), .A(to_acu1[41]), .B(n_43911), .Z(n_38403
		));
	notech_reg to_acu1_reg_42(.CP(n_63113), .D(n_38409), .CD(n_62519), .Q(to_acu1
		[42]));
	notech_mux2 i_41566(.S(n_59321), .A(to_acu1[42]), .B(n_42930), .Z(n_38409
		));
	notech_reg to_acu1_reg_43(.CP(n_63113), .D(n_38415), .CD(n_62519), .Q(to_acu1
		[43]));
	notech_mux2 i_41574(.S(n_59321), .A(to_acu1[43]), .B(n_42933), .Z(n_38415
		));
	notech_reg to_acu1_reg_44(.CP(n_63113), .D(n_38421), .CD(n_62519), .Q(to_acu1
		[44]));
	notech_mux2 i_41582(.S(n_59321), .A(to_acu1[44]), .B(n_42937), .Z(n_38421
		));
	notech_reg to_acu1_reg_45(.CP(n_63117), .D(n_38427), .CD(n_62515), .Q(to_acu1
		[45]));
	notech_mux2 i_41590(.S(n_59321), .A(to_acu1[45]), .B(n_43917), .Z(n_38427
		));
	notech_reg to_acu1_reg_46(.CP(n_63117), .D(n_38433), .CD(n_62519), .Q(to_acu1
		[46]));
	notech_mux2 i_41598(.S(n_59320), .A(to_acu1[46]), .B(n_42941), .Z(n_38433
		));
	notech_reg to_acu1_reg_47(.CP(n_63117), .D(n_38439), .CD(n_62515), .Q(to_acu1
		[47]));
	notech_mux2 i_41606(.S(n_59320), .A(to_acu1[47]), .B(n_42944), .Z(n_38439
		));
	notech_reg to_acu1_reg_48(.CP(n_63117), .D(n_38445), .CD(n_62515), .Q(to_acu1
		[48]));
	notech_mux2 i_41614(.S(n_59320), .A(to_acu1[48]), .B(n_42948), .Z(n_38445
		));
	notech_reg to_acu1_reg_49(.CP(n_63117), .D(n_38451), .CD(n_62515), .Q(to_acu1
		[49]));
	notech_mux2 i_41622(.S(n_59315), .A(to_acu1[49]), .B(n_42951), .Z(n_38451
		));
	notech_reg to_acu1_reg_50(.CP(n_63119), .D(n_38457), .CD(n_62519), .Q(to_acu1
		[50]));
	notech_mux2 i_41630(.S(n_59320), .A(to_acu1[50]), .B(n_42955), .Z(n_38457
		));
	notech_reg to_acu1_reg_51(.CP(n_63119), .D(n_38463), .CD(n_62519), .Q(to_acu1
		[51]));
	notech_mux2 i_41638(.S(n_59320), .A(to_acu1[51]), .B(n_42959), .Z(n_38463
		));
	notech_reg to_acu1_reg_52(.CP(n_63119), .D(n_38469), .CD(n_62519), .Q(to_acu1
		[52]));
	notech_mux2 i_41646(.S(n_59320), .A(to_acu1[52]), .B(n_42962), .Z(n_38469
		));
	notech_reg to_acu1_reg_53(.CP(n_63119), .D(n_38475), .CD(n_62519), .Q(to_acu1
		[53]));
	notech_mux2 i_41654(.S(n_59320), .A(to_acu1[53]), .B(n_42966), .Z(n_38475
		));
	notech_reg to_acu1_reg_54(.CP(n_63119), .D(n_38481), .CD(n_62519), .Q(to_acu1
		[54]));
	notech_mux2 i_41662(.S(n_59320), .A(to_acu1[54]), .B(n_43752), .Z(n_38481
		));
	notech_reg to_acu1_reg_55(.CP(n_63122), .D(n_38487), .CD(n_62521), .Q(to_acu1
		[55]));
	notech_mux2 i_41670(.S(n_59320), .A(to_acu1[55]), .B(n_42969), .Z(n_38487
		));
	notech_reg to_acu1_reg_56(.CP(n_63122), .D(n_38493), .CD(n_62521), .Q(to_acu1
		[56]));
	notech_mux2 i_41678(.S(n_59320), .A(to_acu1[56]), .B(n_42973), .Z(n_38493
		));
	notech_reg to_acu1_reg_57(.CP(n_63122), .D(n_38499), .CD(n_62521), .Q(to_acu1
		[57]));
	notech_mux2 i_41686(.S(n_59320), .A(to_acu1[57]), .B(n_42977), .Z(n_38499
		));
	notech_reg to_acu1_reg_58(.CP(n_63119), .D(n_38505), .CD(n_62521), .Q(to_acu1
		[58]));
	notech_mux2 i_41694(.S(n_59320), .A(to_acu1[58]), .B(n_42980), .Z(n_38505
		));
	notech_reg to_acu1_reg_59(.CP(n_63119), .D(n_38511), .CD(n_62521), .Q(to_acu1
		[59]));
	notech_mux2 i_41702(.S(n_59321), .A(to_acu1[59]), .B(n_42984), .Z(n_38511
		));
	notech_reg to_acu1_reg_60(.CP(n_63119), .D(n_38517), .CD(n_62524), .Q(to_acu1
		[60]));
	notech_mux2 i_41710(.S(n_59304), .A(to_acu1[60]), .B(n_42987), .Z(n_38517
		));
	notech_reg to_acu1_reg_61(.CP(n_63119), .D(n_38523), .CD(n_62524), .Q(to_acu1
		[61]));
	notech_mux2 i_41718(.S(n_59304), .A(to_acu1[61]), .B(n_42991), .Z(n_38523
		));
	notech_reg to_acu1_reg_62(.CP(n_63119), .D(n_38529), .CD(n_62521), .Q(to_acu1
		[62]));
	notech_mux2 i_41726(.S(n_59304), .A(to_acu1[62]), .B(n_42995), .Z(n_38529
		));
	notech_reg to_acu1_reg_63(.CP(n_63119), .D(n_38535), .CD(n_62521), .Q(to_acu1
		[63]));
	notech_mux2 i_41734(.S(n_59304), .A(to_acu1[63]), .B(n_42998), .Z(n_38535
		));
	notech_reg to_acu1_reg_64(.CP(n_63119), .D(n_38541), .CD(n_62521), .Q(to_acu1
		[64]));
	notech_mux2 i_41742(.S(n_59304), .A(to_acu1[64]), .B(n_43002), .Z(n_38541
		));
	notech_reg to_acu1_reg_65(.CP(n_63119), .D(n_38547), .CD(n_62521), .Q(to_acu1
		[65]));
	notech_mux2 i_41750(.S(n_59304), .A(to_acu1[65]), .B(n_43005), .Z(n_38547
		));
	notech_reg to_acu1_reg_66(.CP(n_63119), .D(n_38553), .CD(n_62521), .Q(to_acu1
		[66]));
	notech_mux2 i_41758(.S(n_59304), .A(to_acu1[66]), .B(n_43009), .Z(n_38553
		));
	notech_reg to_acu1_reg_67(.CP(n_63119), .D(n_38559), .CD(n_62521), .Q(to_acu1
		[67]));
	notech_mux2 i_41766(.S(n_59331), .A(to_acu1[67]), .B(n_43013), .Z(n_38559
		));
	notech_reg to_acu1_reg_68(.CP(n_63119), .D(n_38565), .CD(n_62521), .Q(to_acu1
		[68]));
	notech_mux2 i_41774(.S(n_59331), .A(to_acu1[68]), .B(n_43016), .Z(n_38565
		));
	notech_reg to_acu1_reg_69(.CP(n_63119), .D(n_38571), .CD(n_62519), .Q(to_acu1
		[69]));
	notech_mux2 i_41782(.S(n_59331), .A(to_acu1[69]), .B(n_43020), .Z(n_38571
		));
	notech_reg to_acu1_reg_70(.CP(n_63119), .D(n_38577), .CD(n_62521), .Q(to_acu1
		[70]));
	notech_mux2 i_41790(.S(n_59304), .A(to_acu1[70]), .B(n_43023), .Z(n_38577
		));
	notech_reg to_acu1_reg_71(.CP(n_63113), .D(n_38583), .CD(n_62521), .Q(to_acu1
		[71]));
	notech_mux2 i_41798(.S(n_59304), .A(to_acu1[71]), .B(n_43027), .Z(n_38583
		));
	notech_reg to_acu1_reg_72(.CP(n_63111), .D(n_38589), .CD(n_62521), .Q(to_acu1
		[72]));
	notech_mux2 i_41806(.S(n_59331), .A(to_acu1[72]), .B(n_43031), .Z(n_38589
		));
	notech_reg to_acu1_reg_73(.CP(n_63111), .D(n_38595), .CD(n_62521), .Q(to_acu1
		[73]));
	notech_mux2 i_41814(.S(n_59321), .A(to_acu1[73]), .B(n_43035), .Z(n_38595
		));
	notech_reg to_acu1_reg_74(.CP(n_63111), .D(n_38601), .CD(n_62521), .Q(to_acu1
		[74]));
	notech_mux2 i_41822(.S(n_59321), .A(to_acu1[74]), .B(n_43039), .Z(n_38601
		));
	notech_reg to_acu1_reg_75(.CP(n_63111), .D(n_38607), .CD(n_62521), .Q(to_acu1
		[75]));
	notech_mux2 i_41830(.S(n_59321), .A(to_acu1[75]), .B(n_43043), .Z(n_38607
		));
	notech_reg to_acu1_reg_76(.CP(n_63111), .D(n_38613), .CD(n_62513), .Q(to_acu1
		[76]));
	notech_mux2 i_41838(.S(n_59321), .A(to_acu1[76]), .B(n_43046), .Z(n_38613
		));
	notech_reg to_acu1_reg_77(.CP(n_63111), .D(n_38619), .CD(n_62513), .Q(to_acu1
		[77]));
	notech_mux2 i_41846(.S(n_59321), .A(to_acu1[77]), .B(n_43050), .Z(n_38619
		));
	notech_reg to_acu1_reg_78(.CP(n_63111), .D(n_38625), .CD(n_62513), .Q(to_acu1
		[78]));
	notech_mux2 i_41854(.S(n_59321), .A(to_acu1[78]), .B(n_43053), .Z(n_38625
		));
	notech_reg to_acu1_reg_79(.CP(n_63111), .D(n_38631), .CD(n_62513), .Q(to_acu1
		[79]));
	notech_mux2 i_41862(.S(n_59321), .A(to_acu1[79]), .B(n_43057), .Z(n_38631
		));
	notech_reg to_acu1_reg_80(.CP(n_63111), .D(n_38637), .CD(n_62513), .Q(to_acu1
		[80]));
	notech_mux2 i_41870(.S(n_59304), .A(to_acu1[80]), .B(n_43061), .Z(n_38637
		));
	notech_reg to_acu1_reg_81(.CP(n_63111), .D(n_38643), .CD(n_62513), .Q(to_acu1
		[81]));
	notech_mux2 i_41878(.S(n_59304), .A(to_acu1[81]), .B(n_43064), .Z(n_38643
		));
	notech_reg to_acu1_reg_82(.CP(n_63111), .D(n_38649), .CD(n_62513), .Q(to_acu1
		[82]));
	notech_mux2 i_41886(.S(n_59304), .A(to_acu1[82]), .B(n_43068), .Z(n_38649
		));
	notech_reg to_acu1_reg_83(.CP(n_63108), .D(n_38655), .CD(n_62513), .Q(to_acu1
		[83]));
	notech_mux2 i_41894(.S(n_59321), .A(to_acu1[83]), .B(n_43071), .Z(n_38655
		));
	notech_reg to_acu1_reg_84(.CP(n_63108), .D(n_38661), .CD(n_62513), .Q(to_acu1
		[84]));
	notech_mux2 i_41902(.S(n_59321), .A(to_acu1[84]), .B(n_43754), .Z(n_38661
		));
	notech_reg to_acu1_reg_85(.CP(n_63108), .D(n_38667), .CD(n_62513), .Q(to_acu1
		[85]));
	notech_mux2 i_41910(.S(n_59321), .A(to_acu1[85]), .B(n_43075), .Z(n_38667
		));
	notech_reg to_acu1_reg_86(.CP(n_63108), .D(n_38673), .CD(n_62513), .Q(to_acu1
		[86]));
	notech_mux2 i_41918(.S(n_59309), .A(to_acu1[86]), .B(n_43080), .Z(n_38673
		));
	notech_reg to_acu1_reg_87(.CP(n_63108), .D(n_38679), .CD(n_62510), .Q(to_acu1
		[87]));
	notech_mux2 i_41926(.S(n_59309), .A(to_acu1[87]), .B(n_43082), .Z(n_38679
		));
	notech_reg to_acu1_reg_88(.CP(n_63108), .D(n_38685), .CD(n_62510), .Q(to_acu1
		[88]));
	notech_mux2 i_41934(.S(n_59309), .A(to_acu1[88]), .B(n_43085), .Z(n_38685
		));
	notech_reg to_acu1_reg_89(.CP(n_63108), .D(n_38691), .CD(n_62510), .Q(to_acu1
		[89]));
	notech_mux2 i_41942(.S(n_59309), .A(to_acu1[89]), .B(n_43087), .Z(n_38691
		));
	notech_reg to_acu1_reg_90(.CP(n_63108), .D(n_38697), .CD(n_62510), .Q(to_acu1
		[90]));
	notech_mux2 i_41950(.S(n_59309), .A(to_acu1[90]), .B(n_43089), .Z(n_38697
		));
	notech_reg to_acu1_reg_91(.CP(n_63108), .D(n_38703), .CD(n_62510), .Q(to_acu1
		[91]));
	notech_mux2 i_41958(.S(n_59309), .A(to_acu1[91]), .B(n_43093), .Z(n_38703
		));
	notech_reg to_acu1_reg_92(.CP(n_63108), .D(n_38709), .CD(n_62510), .Q(to_acu1
		[92]));
	notech_mux2 i_41966(.S(n_59309), .A(to_acu1[92]), .B(n_43098), .Z(n_38709
		));
	notech_reg to_acu1_reg_93(.CP(n_63113), .D(n_38715), .CD(n_62510), .Q(to_acu1
		[93]));
	notech_mux2 i_41974(.S(n_59309), .A(to_acu1[93]), .B(n_43101), .Z(n_38715
		));
	notech_reg to_acu1_reg_94(.CP(n_63113), .D(n_38721), .CD(n_62510), .Q(to_acu1
		[94]));
	notech_mux2 i_41982(.S(n_59309), .A(to_acu1[94]), .B(n_43104), .Z(n_38721
		));
	notech_reg to_acu1_reg_95(.CP(n_63113), .D(n_38727), .CD(n_62510), .Q(to_acu1
		[95]));
	notech_mux2 i_41990(.S(n_59310), .A(to_acu1[95]), .B(n_43106), .Z(n_38727
		));
	notech_reg to_acu1_reg_96(.CP(n_63113), .D(n_38733), .CD(n_62510), .Q(to_acu1
		[96]));
	notech_mux2 i_41998(.S(n_59309), .A(to_acu1[96]), .B(n_43109), .Z(n_38733
		));
	notech_reg to_acu1_reg_97(.CP(n_63113), .D(n_38739), .CD(n_62515), .Q(to_acu1
		[97]));
	notech_mux2 i_42006(.S(n_59309), .A(to_acu1[97]), .B(n_43111), .Z(n_38739
		));
	notech_reg to_acu1_reg_98(.CP(n_63113), .D(n_38745), .CD(n_62515), .Q(to_acu1
		[98]));
	notech_mux2 i_42014(.S(n_59309), .A(to_acu1[98]), .B(n_43113), .Z(n_38745
		));
	notech_reg to_acu1_reg_99(.CP(n_63113), .D(n_38751), .CD(n_62515), .Q(to_acu1
		[99]));
	notech_mux2 i_42022(.S(n_59304), .A(to_acu1[99]), .B(n_43983), .Z(n_38751
		));
	notech_reg to_acu1_reg_100(.CP(n_63113), .D(n_38757), .CD(n_62515), .Q(to_acu1
		[100]));
	notech_mux2 i_42030(.S(n_59304), .A(to_acu1[100]), .B(n_43986), .Z(n_38757
		));
	notech_reg to_acu1_reg_101(.CP(n_63113), .D(n_38763), .CD(n_62515), .Q(to_acu1
		[101]));
	notech_mux2 i_42038(.S(n_59309), .A(to_acu1[101]), .B(n_43116), .Z(n_38763
		));
	notech_reg to_acu1_reg_102(.CP(n_63113), .D(n_38769), .CD(n_62515), .Q(to_acu1
		[102]));
	notech_mux2 i_42046(.S(n_59304), .A(to_acu1[102]), .B(n_43989), .Z(n_38769
		));
	notech_reg to_acu1_reg_103(.CP(n_63113), .D(n_38775), .CD(n_62515), .Q(to_acu1
		[103]));
	notech_mux2 i_42054(.S(n_59304), .A(to_acu1[103]), .B(n_43992), .Z(n_38775
		));
	notech_reg to_acu1_reg_104(.CP(n_63111), .D(n_38781), .CD(n_62515), .Q(to_acu1
		[104]));
	notech_mux2 i_42062(.S(n_59304), .A(to_acu1[104]), .B(n_43118), .Z(n_38781
		));
	notech_reg to_acu1_reg_105(.CP(n_63111), .D(n_38787), .CD(n_62515), .Q(to_acu1
		[105]));
	notech_mux2 i_42070(.S(n_59309), .A(to_acu1[105]), .B(n_43995), .Z(n_38787
		));
	notech_reg to_acu1_reg_106(.CP(n_63111), .D(n_38793), .CD(n_62515), .Q(to_acu1
		[106]));
	notech_mux2 i_42078(.S(n_59309), .A(to_acu1[106]), .B(n_43121), .Z(n_38793
		));
	notech_reg to_acu1_reg_107(.CP(n_63111), .D(n_38799), .CD(n_62515), .Q(to_acu1
		[107]));
	notech_mux2 i_42086(.S(n_59309), .A(to_acu1[107]), .B(n_43999), .Z(n_38799
		));
	notech_reg to_acu1_reg_108(.CP(n_63111), .D(n_38805), .CD(n_62513), .Q(to_acu1
		[108]));
	notech_mux2 i_42094(.S(n_59309), .A(to_acu1[108]), .B(n_44001), .Z(n_38805
		));
	notech_reg to_acu1_reg_109(.CP(n_63113), .D(n_38811), .CD(n_62513), .Q(to_acu1
		[109]));
	notech_mux2 i_42102(.S(n_59309), .A(to_acu1[109]), .B(n_44004), .Z(n_38811
		));
	notech_reg to_acu1_reg_110(.CP(n_63113), .D(n_38817), .CD(n_62513), .Q(to_acu1
		[110]));
	notech_mux2 i_42110(.S(n_59309), .A(to_acu1[110]), .B(n_44006), .Z(n_38817
		));
	notech_reg to_acu1_reg_111(.CP(n_63113), .D(n_38823), .CD(n_62513), .Q(to_acu1
		[111]));
	notech_mux2 i_42118(.S(n_59309), .A(to_acu1[111]), .B(n_44009), .Z(n_38823
		));
	notech_reg to_acu1_reg_112(.CP(n_63111), .D(n_38829), .CD(n_62513), .Q(to_acu1
		[112]));
	notech_mux2 i_42126(.S(n_59310), .A(to_acu1[112]), .B(n_44011), .Z(n_38829
		));
	notech_reg to_acu1_reg_113(.CP(n_63111), .D(n_38835), .CD(n_62515), .Q(to_acu1
		[113]));
	notech_mux2 i_42134(.S(n_59315), .A(to_acu1[113]), .B(n_43122), .Z(n_38835
		));
	notech_reg to_acu1_reg_114(.CP(n_63129), .D(n_38841), .CD(n_62515), .Q(to_acu1
		[114]));
	notech_mux2 i_42142(.S(n_59315), .A(to_acu1[114]), .B(n_44015), .Z(n_38841
		));
	notech_reg to_acu1_reg_115(.CP(n_63129), .D(n_38847), .CD(n_62515), .Q(to_acu1
		[115]));
	notech_mux2 i_42150(.S(n_59315), .A(to_acu1[115]), .B(n_44017), .Z(n_38847
		));
	notech_reg to_acu1_reg_116(.CP(n_63129), .D(n_38853), .CD(n_62513), .Q(to_acu1
		[116]));
	notech_mux2 i_42158(.S(n_59310), .A(to_acu1[116]), .B(n_44019), .Z(n_38853
		));
	notech_reg to_acu1_reg_117(.CP(n_63129), .D(n_38859), .CD(n_62513), .Q(to_acu1
		[117]));
	notech_mux2 i_42166(.S(n_59310), .A(to_acu1[117]), .B(n_44022), .Z(n_38859
		));
	notech_reg to_acu1_reg_118(.CP(n_63129), .D(n_38865), .CD(n_62524), .Q(to_acu1
		[118]));
	notech_mux2 i_42174(.S(n_59315), .A(to_acu1[118]), .B(n_44024), .Z(n_38865
		));
	notech_reg to_acu1_reg_119(.CP(n_63129), .D(n_38871), .CD(n_62531), .Q(to_acu1
		[119]));
	notech_mux2 i_42182(.S(n_59315), .A(to_acu1[119]), .B(n_44027), .Z(n_38871
		));
	notech_reg to_acu1_reg_120(.CP(n_63129), .D(n_38877), .CD(n_62531), .Q(to_acu1
		[120]));
	notech_mux2 i_42190(.S(n_59315), .A(to_acu1[120]), .B(n_44029), .Z(n_38877
		));
	notech_reg to_acu1_reg_121(.CP(n_63129), .D(n_38883), .CD(n_62531), .Q(to_acu1
		[121]));
	notech_mux2 i_42198(.S(n_59315), .A(to_acu1[121]), .B(n_44031), .Z(n_38883
		));
	notech_reg to_acu1_reg_122(.CP(n_63129), .D(n_38889), .CD(n_62531), .Q(to_acu1
		[122]));
	notech_mux2 i_42206(.S(n_59315), .A(to_acu1[122]), .B(n_44034), .Z(n_38889
		));
	notech_reg to_acu1_reg_123(.CP(n_63129), .D(n_38895), .CD(n_62531), .Q(to_acu1
		[123]));
	notech_mux2 i_42214(.S(n_59315), .A(to_acu1[123]), .B(n_43124), .Z(n_38895
		));
	notech_reg to_acu1_reg_124(.CP(n_63129), .D(n_38901), .CD(n_62531), .Q(to_acu1
		[124]));
	notech_mux2 i_42222(.S(n_59315), .A(to_acu1[124]), .B(n_44037), .Z(n_38901
		));
	notech_reg to_acu1_reg_125(.CP(n_63127), .D(n_38907), .CD(n_62531), .Q(to_acu1
		[125]));
	notech_mux2 i_42230(.S(n_59315), .A(to_acu1[125]), .B(n_43127), .Z(n_38907
		));
	notech_reg to_acu1_reg_126(.CP(n_63127), .D(n_38913), .CD(n_62531), .Q(to_acu1
		[126]));
	notech_mux2 i_42238(.S(n_59310), .A(to_acu1[126]), .B(n_43129), .Z(n_38913
		));
	notech_reg to_acu1_reg_127(.CP(n_63127), .D(n_38919), .CD(n_62531), .Q(to_acu1
		[127]));
	notech_mux2 i_42246(.S(n_59310), .A(to_acu1[127]), .B(n_43130), .Z(n_38919
		));
	notech_reg to_acu1_reg_128(.CP(n_63127), .D(n_38925), .CD(n_62531), .Q(to_acu1
		[128]));
	notech_mux2 i_42254(.S(n_59310), .A(to_acu1[128]), .B(n_43133), .Z(n_38925
		));
	notech_reg to_acu1_reg_129(.CP(n_63127), .D(n_38931), .CD(n_62531), .Q(to_acu1
		[129]));
	notech_mux2 i_42262(.S(n_59310), .A(to_acu1[129]), .B(n_43135), .Z(n_38931
		));
	notech_reg to_acu1_reg_130(.CP(n_63129), .D(n_38937), .CD(n_62529), .Q(to_acu1
		[130]));
	notech_mux2 i_42270(.S(n_59310), .A(to_acu1[130]), .B(n_43137), .Z(n_38937
		));
	notech_reg to_acu1_reg_131(.CP(n_63129), .D(n_38943), .CD(n_62529), .Q(to_acu1
		[131]));
	notech_mux2 i_42278(.S(n_59310), .A(to_acu1[131]), .B(n_43140), .Z(n_38943
		));
	notech_reg to_acu1_reg_132(.CP(n_63127), .D(n_38949), .CD(n_62529), .Q(to_acu1
		[132]));
	notech_mux2 i_42286(.S(n_59310), .A(to_acu1[132]), .B(n_43142), .Z(n_38949
		));
	notech_reg to_acu1_reg_133(.CP(n_63127), .D(n_38955), .CD(n_62529), .Q(to_acu1
		[133]));
	notech_mux2 i_42294(.S(n_59310), .A(to_acu1[133]), .B(n_43145), .Z(n_38955
		));
	notech_reg to_acu1_reg_134(.CP(n_63127), .D(n_38961), .CD(n_62529), .Q(to_acu1
		[134]));
	notech_mux2 i_42302(.S(n_59310), .A(to_acu1[134]), .B(n_43147), .Z(n_38961
		));
	notech_reg to_acu1_reg_135(.CP(n_63133), .D(n_38967), .CD(n_62529), .Q(to_acu1
		[135]));
	notech_mux2 i_42310(.S(n_59310), .A(to_acu1[135]), .B(n_43149), .Z(n_38967
		));
	notech_reg to_acu1_reg_136(.CP(n_63133), .D(n_38973), .CD(n_62531), .Q(to_acu1
		[136]));
	notech_mux2 i_42318(.S(n_59310), .A(to_acu1[136]), .B(n_43152), .Z(n_38973
		));
	notech_reg to_acu1_reg_137(.CP(n_63133), .D(n_38979), .CD(n_62529), .Q(to_acu1
		[137]));
	notech_mux2 i_42326(.S(n_59310), .A(to_acu1[137]), .B(n_43154), .Z(n_38979
		));
	notech_reg to_acu1_reg_138(.CP(n_63133), .D(n_38985), .CD(n_62529), .Q(to_acu1
		[138]));
	notech_mux2 i_42334(.S(n_59310), .A(to_acu1[138]), .B(n_43157), .Z(n_38985
		));
	notech_reg to_acu1_reg_139(.CP(n_63133), .D(n_38991), .CD(n_62529), .Q(to_acu1
		[139]));
	notech_mux2 i_42342(.S(n_59331), .A(to_acu1[139]), .B(n_43159), .Z(n_38991
		));
	notech_reg to_acu1_reg_140(.CP(n_63133), .D(n_38997), .CD(n_62535), .Q(to_acu1
		[140]));
	notech_mux2 i_42350(.S(n_59344), .A(to_acu1[140]), .B(n_43161), .Z(n_38997
		));
	notech_reg to_acu1_reg_141(.CP(n_63133), .D(n_39003), .CD(n_62535), .Q(to_acu1
		[141]));
	notech_mux2 i_42358(.S(n_59344), .A(to_acu1[141]), .B(n_43164), .Z(n_39003
		));
	notech_reg to_acu1_reg_142(.CP(n_63133), .D(n_39009), .CD(n_62535), .Q(to_acu1
		[142]));
	notech_mux2 i_42366(.S(n_59344), .A(to_acu1[142]), .B(n_43166), .Z(n_39009
		));
	notech_reg to_acu1_reg_143(.CP(n_63133), .D(n_39015), .CD(n_62535), .Q(to_acu1
		[143]));
	notech_mux2 i_42374(.S(n_59344), .A(to_acu1[143]), .B(n_43169), .Z(n_39015
		));
	notech_reg to_acu1_reg_144(.CP(n_63133), .D(n_39021), .CD(n_62535), .Q(to_acu1
		[144]));
	notech_mux2 i_42382(.S(n_59344), .A(to_acu1[144]), .B(n_43171), .Z(n_39021
		));
	notech_reg to_acu1_reg_145(.CP(n_63133), .D(n_39027), .CD(n_62535), .Q(to_acu1
		[145]));
	notech_mux2 i_42390(.S(n_59344), .A(to_acu1[145]), .B(n_43173), .Z(n_39027
		));
	notech_reg to_acu1_reg_146(.CP(n_63129), .D(n_39033), .CD(n_62535), .Q(to_acu1
		[146]));
	notech_mux2 i_42398(.S(n_59344), .A(to_acu1[146]), .B(n_43178), .Z(n_39033
		));
	notech_reg to_acu1_reg_147(.CP(n_63129), .D(n_39039), .CD(n_62535), .Q(to_acu1
		[147]));
	notech_mux2 i_42406(.S(n_59344), .A(to_acu1[147]), .B(n_43184), .Z(n_39039
		));
	notech_reg to_acu1_reg_148(.CP(n_63129), .D(n_39045), .CD(n_62535), .Q(to_acu1
		[148]));
	notech_mux2 i_42414(.S(n_59344), .A(to_acu1[148]), .B(n_43190), .Z(n_39045
		));
	notech_reg to_acu1_reg_149(.CP(n_63129), .D(n_39051), .CD(n_62535), .Q(to_acu1
		[149]));
	notech_mux2 i_42422(.S(n_59344), .A(to_acu1[149]), .B(n_43193), .Z(n_39051
		));
	notech_reg to_acu1_reg_150(.CP(n_63129), .D(n_39057), .CD(n_62535), .Q(to_acu1
		[150]));
	notech_mux2 i_42430(.S(n_59344), .A(to_acu1[150]), .B(n_43195), .Z(n_39057
		));
	notech_reg to_acu1_reg_151(.CP(n_63133), .D(n_39063), .CD(n_62531), .Q(to_acu1
		[151]));
	notech_mux2 i_42438(.S(n_59344), .A(to_acu1[151]), .B(n_43197), .Z(n_39063
		));
	notech_reg to_acu1_reg_152(.CP(n_63133), .D(n_39069), .CD(n_62531), .Q(to_acu1
		[152]));
	notech_mux2 i_42446(.S(n_59344), .A(to_acu1[152]), .B(n_43200), .Z(n_39069
		));
	notech_reg to_acu1_reg_153(.CP(n_63133), .D(n_39075), .CD(n_62531), .Q(to_acu1
		[153]));
	notech_mux2 i_42454(.S(n_59343), .A(to_acu1[153]), .B(n_43202), .Z(n_39075
		));
	notech_reg to_acu1_reg_154(.CP(n_63133), .D(n_39081), .CD(n_62531), .Q(to_acu1
		[154]));
	notech_mux2 i_42462(.S(n_59343), .A(to_acu1[154]), .B(n_43205), .Z(n_39081
		));
	notech_reg to_acu1_reg_155(.CP(n_63133), .D(n_39087), .CD(n_62531), .Q(to_acu1
		[155]));
	notech_mux2 i_42470(.S(n_59343), .A(to_acu1[155]), .B(n_43207), .Z(n_39087
		));
	notech_reg to_acu1_reg_156(.CP(n_63127), .D(n_39093), .CD(n_62535), .Q(to_acu1
		[156]));
	notech_mux2 i_42478(.S(n_59343), .A(to_acu1[156]), .B(n_43209), .Z(n_39093
		));
	notech_reg to_acu1_reg_157(.CP(n_63122), .D(n_39099), .CD(n_62535), .Q(to_acu1
		[157]));
	notech_mux2 i_42486(.S(n_59343), .A(to_acu1[157]), .B(n_43212), .Z(n_39099
		));
	notech_reg to_acu1_reg_158(.CP(n_63124), .D(n_39105), .CD(n_62535), .Q(to_acu1
		[158]));
	notech_mux2 i_42494(.S(n_59343), .A(to_acu1[158]), .B(n_43214), .Z(n_39105
		));
	notech_reg to_acu1_reg_159(.CP(n_63122), .D(n_39111), .CD(n_62531), .Q(to_acu1
		[159]));
	notech_mux2 i_42502(.S(n_59343), .A(to_acu1[159]), .B(n_43217), .Z(n_39111
		));
	notech_reg to_acu1_reg_160(.CP(n_63122), .D(n_39117), .CD(n_62535), .Q(to_acu1
		[160]));
	notech_mux2 i_42510(.S(n_59344), .A(to_acu1[160]), .B(n_43219), .Z(n_39117
		));
	notech_reg to_acu1_reg_161(.CP(n_63122), .D(n_39123), .CD(n_62524), .Q(to_acu1
		[161]));
	notech_mux2 i_42518(.S(n_59344), .A(to_acu1[161]), .B(n_43221), .Z(n_39123
		));
	notech_reg to_acu1_reg_162(.CP(n_63124), .D(n_39129), .CD(n_62526), .Q(to_acu1
		[162]));
	notech_mux2 i_42526(.S(n_59344), .A(to_acu1[162]), .B(n_43224), .Z(n_39129
		));
	notech_reg to_acu1_reg_163(.CP(n_63124), .D(n_39135), .CD(n_62524), .Q(to_acu1
		[163]));
	notech_mux2 i_42534(.S(n_59343), .A(to_acu1[163]), .B(n_43226), .Z(n_39135
		));
	notech_reg to_acu1_reg_164(.CP(n_63124), .D(n_39141), .CD(n_62524), .Q(to_acu1
		[164]));
	notech_mux2 i_42542(.S(n_59344), .A(to_acu1[164]), .B(n_43229), .Z(n_39141
		));
	notech_reg to_acu1_reg_165(.CP(n_63124), .D(n_39147), .CD(n_62524), .Q(to_acu1
		[165]));
	notech_mux2 i_42550(.S(n_59344), .A(to_acu1[165]), .B(n_43231), .Z(n_39147
		));
	notech_reg to_acu1_reg_166(.CP(n_63124), .D(n_39153), .CD(n_62526), .Q(to_acu1
		[166]));
	notech_mux2 i_42558(.S(n_59349), .A(to_acu1[166]), .B(n_43233), .Z(n_39153
		));
	notech_reg to_acu1_reg_167(.CP(n_63122), .D(n_39159), .CD(n_62526), .Q(to_acu1
		[167]));
	notech_mux2 i_42566(.S(n_59354), .A(to_acu1[167]), .B(n_43236), .Z(n_39159
		));
	notech_reg to_acu1_reg_168(.CP(n_63122), .D(n_39165), .CD(n_62526), .Q(to_acu1
		[168]));
	notech_mux2 i_42574(.S(n_59354), .A(to_acu1[168]), .B(n_43238), .Z(n_39165
		));
	notech_reg to_acu1_reg_169(.CP(n_63122), .D(n_39171), .CD(n_62526), .Q(to_acu1
		[169]));
	notech_mux2 i_42582(.S(n_59354), .A(to_acu1[169]), .B(n_43241), .Z(n_39171
		));
	notech_reg to_acu1_reg_170(.CP(n_63122), .D(n_39177), .CD(n_62526), .Q(to_acu1
		[170]));
	notech_mux2 i_42590(.S(n_59354), .A(to_acu1[170]), .B(n_43243), .Z(n_39177
		));
	notech_reg to_acu1_reg_171(.CP(n_63122), .D(n_39183), .CD(n_62524), .Q(to_acu1
		[171]));
	notech_mux2 i_42598(.S(n_59354), .A(to_acu1[171]), .B(n_43245), .Z(n_39183
		));
	notech_reg to_acu1_reg_172(.CP(n_63122), .D(n_39189), .CD(n_62524), .Q(to_acu1
		[172]));
	notech_mux2 i_42606(.S(n_59354), .A(to_acu1[172]), .B(n_43248), .Z(n_39189
		));
	notech_reg to_acu1_reg_173(.CP(n_63122), .D(n_39195), .CD(n_62524), .Q(to_acu1
		[173]));
	notech_mux2 i_42614(.S(n_59354), .A(to_acu1[173]), .B(n_43250), .Z(n_39195
		));
	notech_reg to_acu1_reg_174(.CP(n_63122), .D(n_39201), .CD(n_62524), .Q(to_acu1
		[174]));
	notech_mux2 i_42622(.S(n_59354), .A(to_acu1[174]), .B(n_43253), .Z(n_39201
		));
	notech_reg to_acu1_reg_175(.CP(n_63122), .D(n_39207), .CD(n_62524), .Q(to_acu1
		[175]));
	notech_mux2 i_42630(.S(n_59354), .A(to_acu1[175]), .B(n_43255), .Z(n_39207
		));
	notech_reg to_acu1_reg_176(.CP(n_63122), .D(n_39213), .CD(n_62524), .Q(to_acu1
		[176]));
	notech_mux2 i_42638(.S(n_59354), .A(to_acu1[176]), .B(n_42578), .Z(n_39213
		));
	notech_reg to_acu1_reg_177(.CP(n_63122), .D(n_39219), .CD(n_62524), .Q(to_acu1
		[177]));
	notech_mux2 i_42646(.S(n_59354), .A(to_acu1[177]), .B(n_43257), .Z(n_39219
		));
	notech_reg to_acu1_reg_178(.CP(n_63127), .D(n_39225), .CD(n_62524), .Q(to_acu1
		[178]));
	notech_mux2 i_42654(.S(n_59354), .A(to_acu1[178]), .B(n_43757), .Z(n_39225
		));
	notech_reg to_acu1_reg_179(.CP(n_63127), .D(n_39231), .CD(n_62524), .Q(to_acu1
		[179]));
	notech_mux2 i_42662(.S(n_59354), .A(to_acu1[179]), .B(n_43759), .Z(n_39231
		));
	notech_reg to_acu1_reg_180(.CP(n_63127), .D(n_39237), .CD(n_62524), .Q(to_acu1
		[180]));
	notech_mux2 i_42670(.S(n_59349), .A(to_acu1[180]), .B(n_43761), .Z(n_39237
		));
	notech_reg to_acu1_reg_181(.CP(n_63124), .D(n_39243), .CD(n_62524), .Q(to_acu1
		[181]));
	notech_mux2 i_42678(.S(n_59349), .A(to_acu1[181]), .B(n_43764), .Z(n_39243
		));
	notech_reg to_acu1_reg_182(.CP(n_63127), .D(n_39249), .CD(n_62529), .Q(to_acu1
		[182]));
	notech_mux2 i_42686(.S(n_59349), .A(to_acu1[182]), .B(n_43766), .Z(n_39249
		));
	notech_reg to_acu1_reg_183(.CP(n_63127), .D(n_39255), .CD(n_62529), .Q(to_acu1
		[183]));
	notech_mux2 i_42694(.S(n_59349), .A(to_acu1[183]), .B(n_43260), .Z(n_39255
		));
	notech_reg to_acu1_reg_184(.CP(n_63127), .D(n_39261), .CD(n_62529), .Q(to_acu1
		[184]));
	notech_mux2 i_42702(.S(n_59349), .A(to_acu1[184]), .B(n_43262), .Z(n_39261
		));
	notech_reg to_acu1_reg_185(.CP(n_63127), .D(n_39267), .CD(n_62526), .Q(to_acu1
		[185]));
	notech_mux2 i_42710(.S(n_59349), .A(to_acu1[185]), .B(n_43265), .Z(n_39267
		));
	notech_reg to_acu1_reg_186(.CP(n_63127), .D(n_39273), .CD(n_62529), .Q(to_acu1
		[186]));
	notech_mux2 i_42718(.S(n_59349), .A(to_acu1[186]), .B(n_43267), .Z(n_39273
		));
	notech_reg to_acu1_reg_187(.CP(n_63127), .D(n_39279), .CD(n_62529), .Q(to_acu1
		[187]));
	notech_mux2 i_42726(.S(n_59349), .A(to_acu1[187]), .B(n_43269), .Z(n_39279
		));
	notech_reg to_acu1_reg_188(.CP(n_63124), .D(n_39285), .CD(n_62529), .Q(to_acu1
		[188]));
	notech_mux2 i_42734(.S(n_59354), .A(to_acu1[188]), .B(n_43272), .Z(n_39285
		));
	notech_reg to_acu1_reg_189(.CP(n_63124), .D(n_39291), .CD(n_62529), .Q(to_acu1
		[189]));
	notech_mux2 i_42742(.S(n_59354), .A(to_acu1[189]), .B(n_43273), .Z(n_39291
		));
	notech_reg to_acu1_reg_190(.CP(n_63124), .D(n_39297), .CD(n_62529), .Q(to_acu1
		[190]));
	notech_mux2 i_42750(.S(n_59349), .A(to_acu1[190]), .B(n_44117), .Z(n_39297
		));
	notech_reg to_acu1_reg_191(.CP(n_63124), .D(n_39303), .CD(n_62529), .Q(to_acu1
		[191]));
	notech_mux2 i_42758(.S(n_59349), .A(to_acu1[191]), .B(n_44120), .Z(n_39303
		));
	notech_reg to_acu1_reg_192(.CP(n_63124), .D(n_39309), .CD(n_62526), .Q(to_acu1
		[192]));
	notech_mux2 i_42766(.S(n_59349), .A(to_acu1[192]), .B(n_44122), .Z(n_39309
		));
	notech_reg to_acu1_reg_193(.CP(n_63124), .D(n_39315), .CD(n_62526), .Q(to_acu1
		[193]));
	notech_mux2 i_42774(.S(n_59332), .A(to_acu1[193]), .B(n_43274), .Z(n_39315
		));
	notech_reg to_acu1_reg_194(.CP(n_63124), .D(n_39321), .CD(n_62526), .Q(to_acu1
		[194]));
	notech_mux2 i_42782(.S(n_59332), .A(to_acu1[194]), .B(n_43275), .Z(n_39321
		));
	notech_reg to_acu1_reg_195(.CP(n_63124), .D(n_39327), .CD(n_62526), .Q(to_acu1
		[195]));
	notech_mux2 i_42790(.S(n_59332), .A(to_acu1[195]), .B(n_43277), .Z(n_39327
		));
	notech_reg to_acu1_reg_196(.CP(n_63124), .D(n_39333), .CD(n_62526), .Q(to_acu1
		[196]));
	notech_mux2 i_42798(.S(n_59332), .A(to_acu1[196]), .B(n_43278), .Z(n_39333
		));
	notech_reg to_acu1_reg_197(.CP(n_63124), .D(n_39339), .CD(n_62526), .Q(to_acu1
		[197]));
	notech_mux2 i_42806(.S(n_59332), .A(to_acu1[197]), .B(n_43279), .Z(n_39339
		));
	notech_reg to_acu1_reg_198(.CP(n_63124), .D(n_39345), .CD(n_62526), .Q(to_acu1
		[198]));
	notech_mux2 i_42814(.S(n_59332), .A(to_acu1[198]), .B(n_43280), .Z(n_39345
		));
	notech_reg to_acu1_reg_199(.CP(n_63092), .D(n_39351), .CD(n_62526), .Q(to_acu1
		[199]));
	notech_mux2 i_42822(.S(n_59332), .A(to_acu1[199]), .B(n_43281), .Z(n_39351
		));
	notech_reg to_acu1_reg_200(.CP(n_63092), .D(n_39357), .CD(n_62526), .Q(to_acu1
		[200]));
	notech_mux2 i_42830(.S(n_59332), .A(to_acu1[200]), .B(n_43284), .Z(n_39357
		));
	notech_reg to_acu1_reg_201(.CP(n_63092), .D(n_39363), .CD(n_62526), .Q(to_acu1
		[201]));
	notech_mux2 i_42838(.S(n_59332), .A(to_acu1[201]), .B(n_43286), .Z(n_39363
		));
	notech_reg to_acu1_reg_202(.CP(n_63092), .D(n_39369), .CD(n_62526), .Q(to_acu1
		[202]));
	notech_mux2 i_42846(.S(n_59332), .A(to_acu1[202]), .B(n_43289), .Z(n_39369
		));
	notech_reg to_acu1_reg_203(.CP(n_63092), .D(n_39375), .CD(n_62510), .Q(to_acu1
		[203]));
	notech_mux2 i_42854(.S(n_59332), .A(to_acu1[203]), .B(n_43291), .Z(n_39375
		));
	notech_reg to_acu1_reg_204(.CP(n_63092), .D(n_39381), .CD(n_62494), .Q(to_acu1
		[204]));
	notech_mux2 i_42862(.S(n_59332), .A(to_acu1[204]), .B(n_43293), .Z(n_39381
		));
	notech_reg to_acu1_reg_205(.CP(n_63092), .D(n_39387), .CD(n_62494), .Q(to_acu1
		[205]));
	notech_mux2 i_42870(.S(n_59332), .A(to_acu1[205]), .B(n_43296), .Z(n_39387
		));
	notech_reg to_acu1_reg_206(.CP(n_63092), .D(n_39393), .CD(n_62494), .Q(to_acu1
		[206]));
	notech_mux2 i_42878(.S(n_59331), .A(to_acu1[206]), .B(n_43298), .Z(n_39393
		));
	notech_reg to_acu1_reg_207(.CP(n_63092), .D(n_39399), .CD(n_62492), .Q(to_acu1
		[207]));
	notech_mux2 i_42886(.S(n_59331), .A(to_acu1[207]), .B(n_44141), .Z(n_39399
		));
	notech_reg to_acu1_reg_208(.CP(n_63092), .D(n_39405), .CD(n_62494), .Q(to_acu1
		[208]));
	notech_mux2 i_42894(.S(n_59331), .A(to_acu1[208]), .B(n_43301), .Z(n_39405
		));
	notech_reg to_acu1_reg_209(.CP(n_63090), .D(n_39411), .CD(n_62494), .Q(to_acu1
		[209]));
	notech_mux2 i_42902(.S(n_59331), .A(to_acu1[209]), .B(n_44145), .Z(n_39411
		));
	notech_reg to_acu1_reg_210(.CP(n_63090), .D(n_39417), .CD(n_62494), .Q(to_acu1
		[210]));
	notech_mux2 i_42910(.S(n_59331), .A(to_acu1[210]), .B(n_43769), .Z(n_39417
		));
	notech_reg pfx_sz_reg_0(.CP(n_63090), .D(n_39423), .CD(n_62494), .Q(pfx_sz
		[0]));
	notech_mux2 i_42918(.S(\nbus_13538[0] ), .A(pfx_sz[0]), .B(n_42604), .Z(n_39423
		));
	notech_reg pfx_sz_reg_1(.CP(n_63090), .D(n_39429), .CD(n_62494), .Q(pfx_sz
		[1]));
	notech_mux2 i_42926(.S(\nbus_13538[0] ), .A(pfx_sz[1]), .B(n_44149), .Z(n_39429
		));
	notech_reg pfx_sz_reg_2(.CP(n_63090), .D(n_39435), .CD(n_62494), .Q(pfx_sz
		[2]));
	notech_mux2 i_42934(.S(\nbus_13538[0] ), .A(pfx_sz[2]), .B(n_1623100928)
		, .Z(n_39435));
	notech_reg pfx_sz_reg_3(.CP(n_63090), .D(n_39441), .CD(n_62492), .Q(pfx_sz
		[3]));
	notech_mux2 i_42942(.S(\nbus_13538[0] ), .A(pfx_sz[3]), .B(n_1624100929)
		, .Z(n_39441));
	notech_reg pfx_sz_reg_4(.CP(n_63090), .D(n_39447), .CD(n_62492), .Q(pfx_sz
		[4]));
	notech_mux2 i_42950(.S(\nbus_13538[0] ), .A(pfx_sz[4]), .B(n_1625100930)
		, .Z(n_39447));
	notech_reg lenpc2_reg_0(.CP(n_63090), .D(n_39453), .CD(n_62492), .Q(lenpc2
		[0]));
	notech_mux2 i_42958(.S(n_56475), .A(lenpc2[0]), .B(n_1914), .Z(n_39453)
		);
	notech_reg lenpc2_reg_1(.CP(n_63090), .D(n_39459), .CD(n_62492), .Q(lenpc2
		[1]));
	notech_mux2 i_42966(.S(n_56475), .A(lenpc2[1]), .B(n_1516100822), .Z(n_39459
		));
	notech_reg lenpc2_reg_2(.CP(n_63090), .D(n_39465), .CD(n_62492), .Q(lenpc2
		[2]));
	notech_mux2 i_42974(.S(n_56475), .A(lenpc2[2]), .B(n_1518100823), .Z(n_39465
		));
	notech_reg lenpc2_reg_3(.CP(n_63090), .D(n_39471), .CD(n_62492), .Q(lenpc2
		[3]));
	notech_mux2 i_42982(.S(n_56475), .A(lenpc2[3]), .B(n_1519100824), .Z(n_39471
		));
	notech_reg lenpc2_reg_4(.CP(n_63095), .D(n_39477), .CD(n_62492), .Q(lenpc2
		[4]));
	notech_mux2 i_42990(.S(n_56475), .A(lenpc2[4]), .B(n_1520100825), .Z(n_39477
		));
	notech_reg lenpc2_reg_5(.CP(n_63095), .D(n_39483), .CD(n_62492), .Q(lenpc2
		[5]));
	notech_mux2 i_42998(.S(n_56476), .A(lenpc2[5]), .B(n_1559100864), .Z(n_39483
		));
	notech_reg lenpc2_reg_6(.CP(n_63095), .D(n_39493), .CD(n_62492), .Q(lenpc2
		[6]));
	notech_ao3 i_43010(.A(lenpc2[6]), .B(1'b1), .C(n_56487), .Z(n_39493));
	notech_reg lenpc2_reg_7(.CP(n_63095), .D(n_39499), .CD(n_62492), .Q(lenpc2
		[7]));
	notech_ao3 i_43018(.A(lenpc2[7]), .B(1'b1), .C(n_56487), .Z(n_39499));
	notech_reg lenpc2_reg_8(.CP(n_63095), .D(n_39505), .CD(n_62492), .Q(lenpc2
		[8]));
	notech_ao3 i_43026(.A(lenpc2[8]), .B(1'b1), .C(n_56487), .Z(n_39505));
	notech_reg lenpc2_reg_9(.CP(n_63095), .D(n_39511), .CD(n_62497), .Q(lenpc2
		[9]));
	notech_ao3 i_43034(.A(lenpc2[9]), .B(1'b1), .C(n_56482), .Z(n_39511));
	notech_reg lenpc2_reg_10(.CP(n_63095), .D(n_39517), .CD(n_62497), .Q(lenpc2
		[10]));
	notech_ao3 i_43042(.A(lenpc2[10]), .B(1'b1), .C(n_56482), .Z(n_39517));
	notech_reg lenpc2_reg_11(.CP(n_63095), .D(n_39523), .CD(n_62497), .Q(lenpc2
		[11]));
	notech_ao3 i_43050(.A(lenpc2[11]), .B(1'b1), .C(n_56482), .Z(n_39523));
	notech_reg lenpc2_reg_12(.CP(n_63095), .D(n_39529), .CD(n_62497), .Q(lenpc2
		[12]));
	notech_ao3 i_43058(.A(lenpc2[12]), .B(1'b1), .C(n_56487), .Z(n_39529));
	notech_reg lenpc2_reg_13(.CP(n_63095), .D(n_39535), .CD(n_62497), .Q(lenpc2
		[13]));
	notech_ao3 i_43066(.A(lenpc2[13]), .B(1'b1), .C(n_56487), .Z(n_39535));
	notech_reg lenpc2_reg_14(.CP(n_63095), .D(n_39541), .CD(n_62497), .Q(lenpc2
		[14]));
	notech_ao3 i_43074(.A(lenpc2[14]), .B(1'b1), .C(n_56487), .Z(n_39541));
	notech_reg lenpc2_reg_15(.CP(n_63092), .D(n_39547), .CD(n_62497), .Q(lenpc2
		[15]));
	notech_ao3 i_43082(.A(lenpc2[15]), .B(1'b1), .C(n_56487), .Z(n_39547));
	notech_reg lenpc2_reg_16(.CP(n_63092), .D(n_39553), .CD(n_62497), .Q(lenpc2
		[16]));
	notech_ao3 i_43090(.A(lenpc2[16]), .B(1'b1), .C(n_56487), .Z(n_39553));
	notech_reg lenpc2_reg_17(.CP(n_63092), .D(n_39559), .CD(n_62497), .Q(lenpc2
		[17]));
	notech_ao3 i_43098(.A(lenpc2[17]), .B(1'b1), .C(n_56487), .Z(n_39559));
	notech_reg lenpc2_reg_18(.CP(n_63092), .D(n_39565), .CD(n_62497), .Q(lenpc2
		[18]));
	notech_ao3 i_43106(.A(lenpc2[18]), .B(1'b1), .C(n_56487), .Z(n_39565));
	notech_reg lenpc2_reg_19(.CP(n_63092), .D(n_39571), .CD(n_62497), .Q(lenpc2
		[19]));
	notech_ao3 i_43114(.A(lenpc2[19]), .B(1'b1), .C(n_56476), .Z(n_39571));
	notech_reg lenpc2_reg_20(.CP(n_63095), .D(n_39577), .CD(n_62494), .Q(lenpc2
		[20]));
	notech_ao3 i_43122(.A(lenpc2[20]), .B(1'b1), .C(n_56482), .Z(n_39577));
	notech_reg lenpc2_reg_21(.CP(n_63095), .D(n_39583), .CD(n_62494), .Q(lenpc2
		[21]));
	notech_ao3 i_43130(.A(lenpc2[21]), .B(1'b1), .C(n_56482), .Z(n_39583));
	notech_reg lenpc2_reg_22(.CP(n_63092), .D(n_39589), .CD(n_62494), .Q(lenpc2
		[22]));
	notech_ao3 i_43138(.A(lenpc2[22]), .B(1'b1), .C(n_56476), .Z(n_39589));
	notech_reg lenpc2_reg_23(.CP(n_63092), .D(n_39595), .CD(n_62494), .Q(lenpc2
		[23]));
	notech_ao3 i_43146(.A(lenpc2[23]), .B(1'b1), .C(n_56476), .Z(n_39595));
	notech_reg lenpc2_reg_24(.CP(n_63092), .D(n_39601), .CD(n_62494), .Q(lenpc2
		[24]));
	notech_ao3 i_43154(.A(lenpc2[24]), .B(1'b1), .C(n_56476), .Z(n_39601));
	notech_reg lenpc2_reg_25(.CP(n_63090), .D(n_39607), .CD(n_62494), .Q(lenpc2
		[25]));
	notech_ao3 i_43162(.A(lenpc2[25]), .B(1'b1), .C(n_56482), .Z(n_39607));
	notech_reg lenpc2_reg_26(.CP(n_63085), .D(n_39613), .CD(n_62497), .Q(lenpc2
		[26]));
	notech_ao3 i_43170(.A(lenpc2[26]), .B(1'b1), .C(n_56482), .Z(n_39613));
	notech_reg lenpc2_reg_27(.CP(n_63085), .D(n_39619), .CD(n_62494), .Q(lenpc2
		[27]));
	notech_ao3 i_43178(.A(lenpc2[27]), .B(1'b1), .C(n_56482), .Z(n_39619));
	notech_reg lenpc2_reg_28(.CP(n_63085), .D(n_39625), .CD(n_62494), .Q(lenpc2
		[28]));
	notech_ao3 i_43186(.A(lenpc2[28]), .B(1'b1), .C(n_56482), .Z(n_39625));
	notech_reg lenpc2_reg_29(.CP(n_63085), .D(n_39631), .CD(n_62494), .Q(lenpc2
		[29]));
	notech_ao3 i_43194(.A(lenpc2[29]), .B(1'b1), .C(n_56482), .Z(n_39631));
	notech_reg lenpc2_reg_30(.CP(n_63085), .D(n_39637), .CD(n_62487), .Q(lenpc2
		[30]));
	notech_ao3 i_43202(.A(lenpc2[30]), .B(1'b1), .C(n_56482), .Z(n_39637));
	notech_reg lenpc2_reg_31(.CP(n_63087), .D(n_39643), .CD(n_62487), .Q(lenpc2
		[31]));
	notech_ao3 i_43210(.A(lenpc2[31]), .B(1'b1), .C(n_56482), .Z(n_39643));
	notech_reg iack_reg(.CP(n_63087), .D(n_42602), .CD(n_62487), .Q(iack));
	notech_reg over_seg0_reg_5(.CP(n_63087), .D(n_39647), .CD(n_62487), .Q(\over_seg0[5] 
		));
	notech_mux2 i_43218(.S(n_56670), .A(n_42577), .B(\over_seg0[5] ), .Z(n_39647
		));
	notech_reg imm0_reg_0(.CP(n_63085), .D(n_39653), .CD(n_62487), .Q(\imm0[0] 
		));
	notech_mux2 i_43226(.S(n_56670), .A(n_42852), .B(\imm0[0] ), .Z(n_39653)
		);
	notech_reg imm0_reg_1(.CP(n_63085), .D(n_39659), .CD(n_62489), .Q(\imm0[1] 
		));
	notech_mux2 i_43234(.S(n_56640), .A(n_42854), .B(\imm0[1] ), .Z(n_39659)
		);
	notech_reg imm0_reg_2(.CP(n_63085), .D(n_39665), .CD(n_62489), .Q(\imm0[2] 
		));
	notech_mux2 i_43242(.S(n_56640), .A(n_43632), .B(\imm0[2] ), .Z(n_39665)
		);
	notech_reg imm0_reg_3(.CP(n_63085), .D(n_39671), .CD(n_62489), .Q(\imm0[3] 
		));
	notech_mux2 i_43250(.S(n_56670), .A(n_42857), .B(\imm0[3] ), .Z(n_39671)
		);
	notech_reg imm0_reg_4(.CP(n_63085), .D(n_39677), .CD(n_62487), .Q(\imm0[4] 
		));
	notech_mux2 i_43258(.S(n_56670), .A(n_43634), .B(\imm0[4] ), .Z(n_39677)
		);
	notech_reg imm0_reg_5(.CP(n_63085), .D(n_39683), .CD(n_62487), .Q(\imm0[5] 
		));
	notech_mux2 i_43266(.S(n_56670), .A(n_42860), .B(\imm0[5] ), .Z(n_39683)
		);
	notech_reg imm0_reg_6(.CP(n_63085), .D(n_39689), .CD(n_62487), .Q(\imm0[6] 
		));
	notech_mux2 i_43274(.S(n_56670), .A(n_42864), .B(\imm0[6] ), .Z(n_39689)
		);
	notech_reg imm0_reg_7(.CP(n_63085), .D(n_39695), .CD(n_62487), .Q(\imm0[7] 
		));
	notech_mux2 i_43282(.S(n_56640), .A(n_42867), .B(\imm0[7] ), .Z(n_39695)
		);
	notech_reg imm0_reg_8(.CP(n_63085), .D(n_39701), .CD(n_62487), .Q(\imm0[8] 
		));
	notech_mux2 i_43290(.S(n_56640), .A(n_43637), .B(\imm0[8] ), .Z(n_39701)
		);
	notech_reg imm0_reg_9(.CP(n_63085), .D(n_39707), .CD(n_62487), .Q(\imm0[9] 
		));
	notech_mux2 i_43298(.S(n_56640), .A(n_42871), .B(\imm0[9] ), .Z(n_39707)
		);
	notech_reg imm0_reg_10(.CP(n_63085), .D(n_39713), .CD(n_62487), .Q(\imm0[10] 
		));
	notech_mux2 i_43306(.S(n_56640), .A(n_42875), .B(\imm0[10] ), .Z(n_39713
		));
	notech_reg imm0_reg_11(.CP(n_63085), .D(n_39719), .CD(n_62487), .Q(\imm0[11] 
		));
	notech_mux2 i_43314(.S(n_56640), .A(n_43639), .B(\imm0[11] ), .Z(n_39719
		));
	notech_reg imm0_reg_12(.CP(n_63085), .D(n_39725), .CD(n_62487), .Q(\imm0[12] 
		));
	notech_mux2 i_43322(.S(n_56640), .A(n_43641), .B(\imm0[12] ), .Z(n_39725
		));
	notech_reg imm0_reg_13(.CP(n_63087), .D(n_39731), .CD(n_62487), .Q(\imm0[13] 
		));
	notech_mux2 i_43330(.S(n_56640), .A(n_42878), .B(\imm0[13] ), .Z(n_39731
		));
	notech_reg imm0_reg_14(.CP(n_63090), .D(n_39737), .CD(n_62487), .Q(\imm0[14] 
		));
	notech_mux2 i_43338(.S(n_56640), .A(n_42882), .B(\imm0[14] ), .Z(n_39737
		));
	notech_reg imm0_reg_15(.CP(n_63087), .D(n_39743), .CD(n_62487), .Q(\imm0[15] 
		));
	notech_mux2 i_43346(.S(n_56670), .A(n_43644), .B(\imm0[15] ), .Z(n_39743
		));
	notech_reg imm0_reg_16(.CP(n_63087), .D(n_39749), .CD(n_62487), .Q(\imm0[16] 
		));
	notech_mux2 i_43354(.S(n_56674), .A(n_43646), .B(\imm0[16] ), .Z(n_39749
		));
	notech_reg imm0_reg_17(.CP(n_63087), .D(n_39755), .CD(n_62489), .Q(\imm0[17] 
		));
	notech_mux2 i_43362(.S(n_56674), .A(n_43649), .B(\imm0[17] ), .Z(n_39755
		));
	notech_reg imm0_reg_18(.CP(n_63090), .D(n_39761), .CD(n_62492), .Q(\imm0[18] 
		));
	notech_mux2 i_43370(.S(n_56674), .A(n_42885), .B(\imm0[18] ), .Z(n_39761
		));
	notech_reg imm0_reg_19(.CP(n_63090), .D(n_39767), .CD(n_62489), .Q(\imm0[19] 
		));
	notech_mux2 i_43378(.S(n_56674), .A(n_43651), .B(\imm0[19] ), .Z(n_39767
		));
	notech_reg imm0_reg_20(.CP(n_63090), .D(n_39773), .CD(n_62489), .Q(\imm0[20] 
		));
	notech_mux2 i_43386(.S(n_56674), .A(n_42889), .B(\imm0[20] ), .Z(n_39773
		));
	notech_reg imm0_reg_21(.CP(n_63090), .D(n_39779), .CD(n_62489), .Q(\imm0[21] 
		));
	notech_mux2 i_43394(.S(n_56674), .A(n_42893), .B(\imm0[21] ), .Z(n_39779
		));
	notech_reg imm0_reg_22(.CP(n_63090), .D(n_39785), .CD(n_62492), .Q(\imm0[22] 
		));
	notech_mux2 i_43402(.S(n_56674), .A(n_43653), .B(\imm0[22] ), .Z(n_39785
		));
	notech_reg imm0_reg_23(.CP(n_63087), .D(n_39791), .CD(n_62492), .Q(\imm0[23] 
		));
	notech_mux2 i_43410(.S(n_56674), .A(n_42896), .B(\imm0[23] ), .Z(n_39791
		));
	notech_reg imm0_reg_24(.CP(n_63087), .D(n_39797), .CD(n_62492), .Q(\imm0[24] 
		));
	notech_mux2 i_43418(.S(n_56670), .A(n_43656), .B(\imm0[24] ), .Z(n_39797
		));
	notech_reg imm0_reg_25(.CP(n_63087), .D(n_39803), .CD(n_62492), .Q(\imm0[25] 
		));
	notech_mux2 i_43426(.S(n_56670), .A(n_42900), .B(\imm0[25] ), .Z(n_39803
		));
	notech_reg imm0_reg_26(.CP(n_63087), .D(n_39809), .CD(n_62492), .Q(\imm0[26] 
		));
	notech_mux2 i_43434(.S(n_56670), .A(n_43658), .B(\imm0[26] ), .Z(n_39809
		));
	notech_reg imm0_reg_27(.CP(n_63087), .D(n_39815), .CD(n_62489), .Q(\imm0[27] 
		));
	notech_mux2 i_43442(.S(n_56670), .A(n_43661), .B(\imm0[27] ), .Z(n_39815
		));
	notech_reg imm0_reg_28(.CP(n_63087), .D(n_39821), .CD(n_62489), .Q(\imm0[28] 
		));
	notech_mux2 i_43450(.S(n_56670), .A(n_43663), .B(\imm0[28] ), .Z(n_39821
		));
	notech_reg imm0_reg_29(.CP(n_63087), .D(n_39827), .CD(n_62489), .Q(\imm0[29] 
		));
	notech_mux2 i_43458(.S(n_56670), .A(n_43665), .B(\imm0[29] ), .Z(n_39827
		));
	notech_reg imm0_reg_30(.CP(n_63087), .D(n_39833), .CD(n_62489), .Q(\imm0[30] 
		));
	notech_mux2 i_43466(.S(n_56670), .A(n_43668), .B(\imm0[30] ), .Z(n_39833
		));
	notech_reg imm0_reg_31(.CP(n_63087), .D(n_39839), .CD(n_62489), .Q(\imm0[31] 
		));
	notech_mux2 i_43474(.S(n_56670), .A(n_43670), .B(\imm0[31] ), .Z(n_39839
		));
	notech_reg imm0_reg_32(.CP(n_63087), .D(n_39845), .CD(n_62489), .Q(\imm0[32] 
		));
	notech_mux2 i_43482(.S(n_56655), .A(n_43673), .B(\imm0[32] ), .Z(n_39845
		));
	notech_reg imm0_reg_33(.CP(n_63087), .D(n_39851), .CD(n_62489), .Q(\imm0[33] 
		));
	notech_mux2 i_43490(.S(n_56655), .A(n_43675), .B(\imm0[33] ), .Z(n_39851
		));
	notech_reg imm0_reg_34(.CP(n_63103), .D(n_39857), .CD(n_62489), .Q(\imm0[34] 
		));
	notech_mux2 i_43498(.S(n_56655), .A(n_43677), .B(\imm0[34] ), .Z(n_39857
		));
	notech_reg imm0_reg_35(.CP(n_63103), .D(n_39863), .CD(n_62489), .Q(\imm0[35] 
		));
	notech_mux2 i_43506(.S(n_56655), .A(n_43680), .B(\imm0[35] ), .Z(n_39863
		));
	notech_reg imm0_reg_36(.CP(n_63103), .D(n_39869), .CD(n_62489), .Q(\imm0[36] 
		));
	notech_mux2 i_43514(.S(n_56660), .A(n_43682), .B(\imm0[36] ), .Z(n_39869
		));
	notech_reg imm0_reg_37(.CP(n_63103), .D(n_39875), .CD(n_62489), .Q(\imm0[37] 
		));
	notech_mux2 i_43522(.S(n_56660), .A(n_43685), .B(\imm0[37] ), .Z(n_39875
		));
	notech_reg imm0_reg_38(.CP(n_63103), .D(n_39881), .CD(n_62497), .Q(\imm0[38] 
		));
	notech_mux2 i_43530(.S(n_56655), .A(n_42575), .B(\imm0[38] ), .Z(n_39881
		));
	notech_reg imm0_reg_39(.CP(n_63106), .D(n_39887), .CD(n_62505), .Q(\imm0[39] 
		));
	notech_mux2 i_43538(.S(n_56660), .A(n_43687), .B(\imm0[39] ), .Z(n_39887
		));
	notech_reg imm0_reg_40(.CP(n_63106), .D(n_39893), .CD(n_62505), .Q(\imm0[40] 
		));
	notech_mux2 i_43546(.S(n_56655), .A(n_43689), .B(\imm0[40] ), .Z(n_39893
		));
	notech_reg imm0_reg_41(.CP(n_63106), .D(n_39899), .CD(n_62505), .Q(\imm0[41] 
		));
	notech_mux2 i_43554(.S(n_56655), .A(n_43692), .B(\imm0[41] ), .Z(n_39899
		));
	notech_reg imm0_reg_42(.CP(n_63106), .D(n_39905), .CD(n_62505), .Q(\imm0[42] 
		));
	notech_mux2 i_43562(.S(n_56655), .A(n_43694), .B(\imm0[42] ), .Z(n_39905
		));
	notech_reg imm0_reg_43(.CP(n_63106), .D(n_39911), .CD(n_62505), .Q(\imm0[43] 
		));
	notech_mux2 i_43570(.S(n_56655), .A(n_43697), .B(\imm0[43] ), .Z(n_39911
		));
	notech_reg imm0_reg_44(.CP(n_63103), .D(n_39917), .CD(n_62508), .Q(\imm0[44] 
		));
	notech_mux2 i_43578(.S(n_56655), .A(n_43699), .B(\imm0[44] ), .Z(n_39917
		));
	notech_reg imm0_reg_45(.CP(n_63103), .D(n_39923), .CD(n_62508), .Q(\imm0[45] 
		));
	notech_mux2 i_43586(.S(n_56655), .A(n_43701), .B(\imm0[45] ), .Z(n_39923
		));
	notech_reg imm0_reg_46(.CP(n_63103), .D(n_39929), .CD(n_62508), .Q(\imm0[46] 
		));
	notech_mux2 i_43594(.S(n_56655), .A(n_43704), .B(\imm0[46] ), .Z(n_39929
		));
	notech_reg imm0_reg_47(.CP(n_63103), .D(n_39935), .CD(n_62505), .Q(\imm0[47] 
		));
	notech_mux2 i_43602(.S(n_56655), .A(n_43706), .B(\imm0[47] ), .Z(n_39935
		));
	notech_reg lenpc1_reg_0(.CP(n_63103), .D(n_39941), .CD(n_62508), .Q(lenpc1
		[0]));
	notech_mux2 i_43610(.S(n_59331), .A(lenpc1[0]), .B(n_42574), .Z(n_39941)
		);
	notech_reg lenpc1_reg_1(.CP(n_63103), .D(n_39947), .CD(n_62505), .Q(lenpc1
		[1]));
	notech_mux2 i_43618(.S(n_59331), .A(lenpc1[1]), .B(n_44173), .Z(n_39947)
		);
	notech_reg lenpc1_reg_2(.CP(n_63103), .D(n_39953), .CD(n_62505), .Q(lenpc1
		[2]));
	notech_mux2 i_43626(.S(n_59331), .A(lenpc1[2]), .B(n_44175), .Z(n_39953)
		);
	notech_reg lenpc1_reg_3(.CP(n_63103), .D(n_39959), .CD(n_62505), .Q(lenpc1
		[3]));
	notech_mux2 i_43634(.S(n_59331), .A(lenpc1[3]), .B(n_44177), .Z(n_39959)
		);
	notech_reg lenpc1_reg_4(.CP(n_63103), .D(n_39965), .CD(n_62505), .Q(lenpc1
		[4]));
	notech_mux2 i_43642(.S(n_59331), .A(lenpc1[4]), .B(n_44180), .Z(n_39965)
		);
	notech_reg lenpc1_reg_5(.CP(n_63103), .D(n_39971), .CD(n_62505), .Q(lenpc1
		[5]));
	notech_mux2 i_43650(.S(n_59331), .A(lenpc1[5]), .B(n_44182), .Z(n_39971)
		);
	notech_reg lenpc1_reg_6(.CP(n_63103), .D(n_39977), .CD(n_62505), .Q(lenpc1
		[6]));
	notech_mux2 i_43658(.S(n_59331), .A(lenpc1[6]), .B(n_1493100799), .Z(n_39977
		));
	notech_reg lenpc1_reg_7(.CP(n_63108), .D(n_39983), .CD(n_62505), .Q(lenpc1
		[7]));
	notech_mux2 i_43666(.S(n_59331), .A(lenpc1[7]), .B(n_44100), .Z(n_39983)
		);
	notech_reg lenpc1_reg_8(.CP(n_63108), .D(n_39989), .CD(n_62505), .Q(lenpc1
		[8]));
	notech_mux2 i_43674(.S(n_59332), .A(lenpc1[8]), .B(n_1494100800), .Z(n_39989
		));
	notech_reg lenpc1_reg_9(.CP(n_63108), .D(n_39995), .CD(n_62505), .Q(lenpc1
		[9]));
	notech_mux2 i_43682(.S(n_59343), .A(lenpc1[9]), .B(n_1495100801), .Z(n_39995
		));
	notech_reg lenpc1_reg_10(.CP(n_63106), .D(n_40001), .CD(n_62505), .Q(lenpc1
		[10]));
	notech_mux2 i_43690(.S(n_59343), .A(lenpc1[10]), .B(n_44118), .Z(n_40001
		));
	notech_reg lenpc1_reg_11(.CP(n_63106), .D(n_40007), .CD(n_62505), .Q(lenpc1
		[11]));
	notech_mux2 i_43698(.S(n_59343), .A(lenpc1[11]), .B(n_1496100802), .Z(n_40007
		));
	notech_reg lenpc1_reg_12(.CP(n_63108), .D(n_40013), .CD(n_62510), .Q(lenpc1
		[12]));
	notech_mux2 i_43706(.S(n_59338), .A(lenpc1[12]), .B(n_1497100803), .Z(n_40013
		));
	notech_reg lenpc1_reg_13(.CP(n_63108), .D(n_40019), .CD(n_62510), .Q(lenpc1
		[13]));
	notech_mux2 i_43714(.S(n_59338), .A(lenpc1[13]), .B(n_1498100804), .Z(n_40019
		));
	notech_reg lenpc1_reg_14(.CP(n_63108), .D(n_40025), .CD(n_62508), .Q(lenpc1
		[14]));
	notech_mux2 i_43722(.S(n_59338), .A(lenpc1[14]), .B(n_1499100805), .Z(n_40025
		));
	notech_reg lenpc1_reg_15(.CP(n_63108), .D(n_40031), .CD(n_62508), .Q(lenpc1
		[15]));
	notech_mux2 i_43730(.S(n_59343), .A(lenpc1[15]), .B(n_1500100806), .Z(n_40031
		));
	notech_reg lenpc1_reg_16(.CP(n_63108), .D(n_40037), .CD(n_62508), .Q(lenpc1
		[16]));
	notech_mux2 i_43738(.S(n_59343), .A(lenpc1[16]), .B(n_1501100807), .Z(n_40037
		));
	notech_reg lenpc1_reg_17(.CP(n_63106), .D(n_40043), .CD(n_62510), .Q(lenpc1
		[17]));
	notech_mux2 i_43746(.S(n_59343), .A(lenpc1[17]), .B(n_1502100808), .Z(n_40043
		));
	notech_reg lenpc1_reg_18(.CP(n_63106), .D(n_40049), .CD(n_62510), .Q(lenpc1
		[18]));
	notech_mux2 i_43754(.S(n_59343), .A(lenpc1[18]), .B(n_1503100809), .Z(n_40049
		));
	notech_reg lenpc1_reg_19(.CP(n_63106), .D(n_40055), .CD(n_62510), .Q(lenpc1
		[19]));
	notech_mux2 i_43762(.S(n_59343), .A(lenpc1[19]), .B(n_1504100810), .Z(n_40055
		));
	notech_reg lenpc1_reg_20(.CP(n_63106), .D(n_40061), .CD(n_62510), .Q(lenpc1
		[20]));
	notech_mux2 i_43770(.S(n_59343), .A(lenpc1[20]), .B(n_1505100811), .Z(n_40061
		));
	notech_reg lenpc1_reg_21(.CP(n_63106), .D(n_40067), .CD(n_62510), .Q(lenpc1
		[21]));
	notech_mux2 i_43778(.S(n_59343), .A(lenpc1[21]), .B(n_1506100812), .Z(n_40067
		));
	notech_reg lenpc1_reg_22(.CP(n_63106), .D(n_40073), .CD(n_62508), .Q(lenpc1
		[22]));
	notech_mux2 i_43786(.S(n_59332), .A(lenpc1[22]), .B(n_1507100813), .Z(n_40073
		));
	notech_reg lenpc1_reg_23(.CP(n_63106), .D(n_40079), .CD(n_62508), .Q(lenpc1
		[23]));
	notech_mux2 i_43794(.S(n_59338), .A(lenpc1[23]), .B(n_1508100814), .Z(n_40079
		));
	notech_nao3 i_22678823(.A(n_60854), .B(n_44744), .C(n_229999378), .Z(n_194199020
		));
	notech_reg lenpc1_reg_24(.CP(n_63106), .D(n_40085), .CD(n_62508), .Q(lenpc1
		[24]));
	notech_mux2 i_43802(.S(n_59338), .A(lenpc1[24]), .B(n_1509100815), .Z(n_40085
		));
	notech_nao3 i_3179010(.A(n_2997), .B(n_42611), .C(n_2975), .Z(n_194099019
		));
	notech_reg lenpc1_reg_25(.CP(n_63106), .D(n_40091), .CD(n_62508), .Q(lenpc1
		[25]));
	notech_mux2 i_43810(.S(n_59332), .A(lenpc1[25]), .B(n_1510100816), .Z(n_40091
		));
	notech_ao4 i_126479397(.A(n_59153), .B(n_43079), .C(n_60127), .D(n_44374
		), .Z(n_193999018));
	notech_reg lenpc1_reg_26(.CP(n_63106), .D(n_40097), .CD(n_62508), .Q(lenpc1
		[26]));
	notech_mux2 i_43818(.S(n_59332), .A(lenpc1[26]), .B(n_1511100817), .Z(n_40097
		));
	notech_ao4 i_126579396(.A(n_59153), .B(n_43081), .C(n_60127), .D(n_44376
		), .Z(n_193899017));
	notech_reg lenpc1_reg_27(.CP(n_63106), .D(n_40103), .CD(n_62508), .Q(lenpc1
		[27]));
	notech_mux2 i_43826(.S(n_59332), .A(lenpc1[27]), .B(n_1512100818), .Z(n_40103
		));
	notech_ao4 i_126679395(.A(n_59153), .B(n_43083), .C(n_60127), .D(n_44377
		), .Z(n_193799016));
	notech_reg lenpc1_reg_28(.CP(n_63103), .D(n_40109), .CD(n_62508), .Q(lenpc1
		[28]));
	notech_mux2 i_43834(.S(n_59338), .A(lenpc1[28]), .B(n_1513100819), .Z(n_40109
		));
	notech_ao4 i_126779394(.A(n_59153), .B(n_43086), .C(n_60127), .D(n_44378
		), .Z(n_193699015));
	notech_reg lenpc1_reg_29(.CP(n_63097), .D(n_40115), .CD(n_62508), .Q(lenpc1
		[29]));
	notech_mux2 i_43842(.S(n_59338), .A(lenpc1[29]), .B(n_1514100820), .Z(n_40115
		));
	notech_ao4 i_126879393(.A(n_59151), .B(n_43088), .C(n_60127), .D(n_44379
		), .Z(n_193599014));
	notech_reg lenpc1_reg_30(.CP(n_63097), .D(n_40121), .CD(n_62508), .Q(lenpc1
		[30]));
	notech_mux2 i_43850(.S(n_59338), .A(lenpc1[30]), .B(n_1515100821), .Z(n_40121
		));
	notech_ao4 i_126979392(.A(n_59151), .B(n_43092), .C(n_60127), .D(n_44380
		), .Z(n_193499013));
	notech_reg lenpc1_reg_31(.CP(n_63097), .D(n_40127), .CD(n_62508), .Q(lenpc1
		[31]));
	notech_mux2 i_43858(.S(n_59338), .A(lenpc1[31]), .B(n_1195100503), .Z(n_40127
		));
	notech_ao4 i_127079391(.A(n_59151), .B(n_43094), .C(n_60127), .D(n_44382
		), .Z(n_193399012));
	notech_reg lenpc_reg_0(.CP(n_63097), .D(n_40133), .CD(n_62508), .Q(lenpc
		[0]));
	notech_mux2 i_43866(.S(n_3303), .A(n_44189), .B(lenpc[0]), .Z(n_40133)
		);
	notech_ao4 i_127179390(.A(n_59151), .B(n_43097), .C(n_60125), .D(n_44383
		), .Z(n_193299011));
	notech_reg lenpc_reg_1(.CP(n_63097), .D(n_40139), .CD(n_62499), .Q(lenpc
		[1]));
	notech_mux2 i_43874(.S(n_3303), .A(n_44191), .B(lenpc[1]), .Z(n_40139)
		);
	notech_ao4 i_127979382(.A(n_59151), .B(n_43117), .C(n_60125), .D(n_44392
		), .Z(n_193199010));
	notech_reg lenpc_reg_2(.CP(n_63097), .D(n_40145), .CD(n_62499), .Q(lenpc
		[2]));
	notech_mux2 i_43882(.S(n_3303), .A(n_44192), .B(lenpc[2]), .Z(n_40145)
		);
	notech_ao4 i_128379378(.A(n_59151), .B(n_43128), .C(n_60125), .D(n_44398
		), .Z(n_193099009));
	notech_reg lenpc_reg_3(.CP(n_63097), .D(n_40151), .CD(n_62499), .Q(lenpc
		[3]));
	notech_mux2 i_43890(.S(n_3303), .A(n_44193), .B(lenpc[3]), .Z(n_40151)
		);
	notech_ao4 i_128679375(.A(n_59151), .B(n_43136), .C(n_60125), .D(n_44403
		), .Z(n_192999008));
	notech_reg lenpc_reg_4(.CP(n_63097), .D(n_40157), .CD(n_62499), .Q(lenpc
		[4]));
	notech_mux2 i_43898(.S(n_3303), .A(n_44194), .B(lenpc[4]), .Z(n_40157)
		);
	notech_ao4 i_128779374(.A(n_59151), .B(n_43139), .C(n_60125), .D(n_44404
		), .Z(n_192899007));
	notech_reg lenpc_reg_5(.CP(n_63097), .D(n_40163), .CD(n_62499), .Q(lenpc
		[5]));
	notech_mux2 i_43906(.S(n_3303), .A(n_44195), .B(lenpc[5]), .Z(n_40163)
		);
	notech_ao4 i_128879373(.A(n_59151), .B(n_43141), .C(n_60125), .D(n_44406
		), .Z(n_192799006));
	notech_reg lenpc_reg_6(.CP(n_63097), .D(n_40169), .CD(n_62499), .Q(lenpc
		[6]));
	notech_mux2 i_43914(.S(n_3303), .A(n_1181100489), .B(lenpc[6]), .Z(n_40169
		));
	notech_ao4 i_128979372(.A(n_59153), .B(n_43143), .C(n_60125), .D(n_44407
		), .Z(n_192699005));
	notech_reg lenpc_reg_7(.CP(n_63097), .D(n_40175), .CD(n_62499), .Q(lenpc
		[7]));
	notech_mux2 i_43922(.S(n_3303), .A(n_1182100490), .B(lenpc[7]), .Z(n_40175
		));
	notech_ao4 i_129079371(.A(n_59151), .B(n_43146), .C(n_60125), .D(n_44408
		), .Z(n_192599004));
	notech_reg lenpc_reg_8(.CP(n_63095), .D(n_40181), .CD(n_62499), .Q(lenpc
		[8]));
	notech_mux2 i_43930(.S(n_3303), .A(n_1183100491), .B(lenpc[8]), .Z(n_40181
		));
	notech_ao4 i_129179370(.A(n_59151), .B(n_43148), .C(n_60125), .D(n_44409
		), .Z(n_192499003));
	notech_reg lenpc_reg_9(.CP(n_63095), .D(n_40187), .CD(n_62499), .Q(lenpc
		[9]));
	notech_mux2 i_43938(.S(n_3303), .A(n_1184100492), .B(lenpc[9]), .Z(n_40187
		));
	notech_ao4 i_129279369(.A(n_59151), .B(n_43151), .C(n_60125), .D(n_44410
		), .Z(n_192399002));
	notech_reg lenpc_reg_10(.CP(n_63095), .D(n_40193), .CD(n_62499), .Q(lenpc
		[10]));
	notech_mux2 i_43946(.S(n_3303), .A(n_1185100493), .B(lenpc[10]), .Z(n_40193
		));
	notech_ao4 i_129479367(.A(n_59151), .B(n_43155), .C(n_60125), .D(n_44413
		), .Z(n_192299001));
	notech_reg lenpc_reg_11(.CP(n_63095), .D(n_40199), .CD(n_62499), .Q(lenpc
		[11]));
	notech_mux2 i_43954(.S(n_3303), .A(n_1186100494), .B(lenpc[11]), .Z(n_40199
		));
	notech_ao4 i_129979362(.A(n_59146), .B(n_43167), .C(n_60125), .D(n_44419
		), .Z(n_192199000));
	notech_reg lenpc_reg_12(.CP(n_63095), .D(n_40205), .CD(n_62497), .Q(lenpc
		[12]));
	notech_mux2 i_43962(.S(n_3303), .A(n_1187100495), .B(lenpc[12]), .Z(n_40205
		));
	notech_ao4 i_130579356(.A(n_59139), .B(n_43183), .C(n_60125), .D(n_44426
		), .Z(n_192098999));
	notech_reg lenpc_reg_13(.CP(n_63097), .D(n_40211), .CD(n_62497), .Q(lenpc
		[13]));
	notech_mux2 i_43970(.S(n_3303), .A(n_1188100496), .B(lenpc[13]), .Z(n_40211
		));
	notech_ao4 i_130879353(.A(n_59139), .B(n_43191), .C(n_60125), .D(n_44429
		), .Z(n_191998998));
	notech_reg lenpc_reg_14(.CP(n_63097), .D(n_40217), .CD(n_62497), .Q(lenpc
		[14]));
	notech_mux2 i_43978(.S(n_3303), .A(n_1189100497), .B(lenpc[14]), .Z(n_40217
		));
	notech_ao4 i_130979352(.A(n_59141), .B(n_43194), .C(n_60125), .D(n_44430
		), .Z(n_191898997));
	notech_reg lenpc_reg_15(.CP(n_63097), .D(n_40223), .CD(n_62497), .Q(lenpc
		[15]));
	notech_mux2 i_43986(.S(n_3303), .A(n_1190100498), .B(lenpc[15]), .Z(n_40223
		));
	notech_ao4 i_131279349(.A(n_59139), .B(n_43201), .C(n_60125), .D(n_44433
		), .Z(n_1917));
	notech_reg lenpc_reg_16(.CP(n_63097), .D(n_40229), .CD(n_62497), .Q(lenpc
		[16]));
	notech_mux2 i_43994(.S(n_55782), .A(n_1191100499), .B(lenpc[16]), .Z(n_40229
		));
	notech_ao4 i_131779344(.A(n_59139), .B(n_43213), .C(n_60112), .D(n_44439
		), .Z(n_1916));
	notech_reg lenpc_reg_17(.CP(n_63097), .D(n_40235), .CD(n_62499), .Q(lenpc
		[17]));
	notech_mux2 i_44002(.S(n_55782), .A(n_1192100500), .B(lenpc[17]), .Z(n_40235
		));
	notech_ao4 i_132079341(.A(n_59139), .B(n_43220), .C(n_60112), .D(n_44443
		), .Z(n_1911));
	notech_reg lenpc_reg_18(.CP(n_63101), .D(n_40241), .CD(n_62499), .Q(lenpc
		[18]));
	notech_mux2 i_44010(.S(n_55782), .A(n_1193100501), .B(lenpc[18]), .Z(n_40241
		));
	notech_ao4 i_132779334(.A(n_59139), .B(n_43237), .C(n_60112), .D(n_44451
		), .Z(n_1897));
	notech_reg lenpc_reg_19(.CP(n_63101), .D(n_40247), .CD(n_62499), .Q(lenpc
		[19]));
	notech_mux2 i_44018(.S(n_55782), .A(n_1622100927), .B(lenpc[19]), .Z(n_40247
		));
	notech_ao4 i_132879333(.A(n_59141), .B(n_43239), .C(n_60112), .D(n_44452
		), .Z(n_1896));
	notech_reg lenpc_reg_20(.CP(n_63101), .D(n_40253), .CD(n_62499), .Q(lenpc
		[20]));
	notech_mux2 i_44026(.S(n_55782), .A(n_1194100502), .B(lenpc[20]), .Z(n_40253
		));
	notech_ao4 i_132979332(.A(n_59141), .B(n_43242), .C(n_60112), .D(n_44453
		), .Z(n_1895));
	notech_reg lenpc_reg_21(.CP(n_63101), .D(n_40259), .CD(n_62499), .Q(lenpc
		[21]));
	notech_mux2 i_44034(.S(n_55782), .A(n_1482100788), .B(lenpc[21]), .Z(n_40259
		));
	notech_ao4 i_133079331(.A(n_59141), .B(n_43244), .C(n_60112), .D(n_44454
		), .Z(n_1894));
	notech_reg lenpc_reg_22(.CP(n_63101), .D(n_40265), .CD(n_62503), .Q(lenpc
		[22]));
	notech_mux2 i_44042(.S(n_55782), .A(n_1483100789), .B(lenpc[22]), .Z(n_40265
		));
	notech_ao4 i_133179330(.A(n_59141), .B(n_43247), .C(n_60112), .D(n_44455
		), .Z(n_1893));
	notech_reg lenpc_reg_23(.CP(n_63101), .D(n_40271), .CD(n_62503), .Q(lenpc
		[23]));
	notech_mux2 i_44050(.S(n_55782), .A(n_1484100790), .B(lenpc[23]), .Z(n_40271
		));
	notech_ao4 i_133279329(.A(n_59141), .B(n_43249), .C(n_60112), .D(n_44456
		), .Z(n_1891));
	notech_reg lenpc_reg_24(.CP(n_63103), .D(n_40277), .CD(n_62503), .Q(lenpc
		[24]));
	notech_mux2 i_44058(.S(n_55782), .A(n_1485100791), .B(lenpc[24]), .Z(n_40277
		));
	notech_ao4 i_133379328(.A(n_59141), .B(n_43251), .C(n_60112), .D(n_44457
		), .Z(n_1890));
	notech_reg lenpc_reg_25(.CP(n_63101), .D(n_40283), .CD(n_62503), .Q(lenpc
		[25]));
	notech_mux2 i_44066(.S(n_55782), .A(n_1486100792), .B(lenpc[25]), .Z(n_40283
		));
	notech_ao4 i_133479327(.A(n_59141), .B(n_43254), .C(n_60112), .D(n_44458
		), .Z(n_1889));
	notech_reg lenpc_reg_26(.CP(n_63101), .D(n_40289), .CD(n_62503), .Q(lenpc
		[26]));
	notech_mux2 i_44074(.S(n_55782), .A(n_1487100793), .B(lenpc[26]), .Z(n_40289
		));
	notech_ao4 i_133579326(.A(n_59139), .B(n_43256), .C(n_60112), .D(n_44459
		), .Z(n_1888));
	notech_reg lenpc_reg_27(.CP(n_63101), .D(n_40295), .CD(n_62503), .Q(lenpc
		[27]));
	notech_mux2 i_44082(.S(n_55782), .A(n_1488100794), .B(lenpc[27]), .Z(n_40295
		));
	notech_ao4 i_133779324(.A(n_59138), .B(n_43261), .C(n_60112), .D(n_44461
		), .Z(n_1887));
	notech_reg lenpc_reg_28(.CP(n_63101), .D(n_40301), .CD(n_62505), .Q(lenpc
		[28]));
	notech_mux2 i_44090(.S(n_55782), .A(n_1489100795), .B(lenpc[28]), .Z(n_40301
		));
	notech_ao4 i_133879323(.A(n_59138), .B(n_43263), .C(n_60112), .D(n_44462
		), .Z(n_1886));
	notech_reg lenpc_reg_29(.CP(n_63101), .D(n_40307), .CD(n_62503), .Q(lenpc
		[29]));
	notech_mux2 i_44098(.S(n_55782), .A(n_1490100796), .B(lenpc[29]), .Z(n_40307
		));
	notech_ao4 i_133979322(.A(n_59138), .B(n_43266), .C(n_60112), .D(n_44463
		), .Z(n_1885));
	notech_reg lenpc_reg_30(.CP(n_63101), .D(n_40313), .CD(n_62503), .Q(lenpc
		[30]));
	notech_mux2 i_44106(.S(n_55782), .A(n_1491100797), .B(lenpc[30]), .Z(n_40313
		));
	notech_ao4 i_134079321(.A(n_59138), .B(n_43268), .C(n_60112), .D(n_44464
		), .Z(n_188498996));
	notech_reg lenpc_reg_31(.CP(n_63101), .D(n_40319), .CD(n_62503), .Q(lenpc
		[31]));
	notech_mux2 i_44114(.S(n_55782), .A(n_1492100798), .B(lenpc[31]), .Z(n_40319
		));
	notech_ao4 i_134179320(.A(n_59138), .B(n_43271), .C(n_60112), .D(n_44466
		), .Z(n_188398995));
	notech_reg opz1_reg_0(.CP(n_63097), .D(n_40325), .CD(n_62503), .Q(opz1[0
		]));
	notech_mux2 i_44122(.S(n_59338), .A(opz1[0]), .B(n_43627), .Z(n_40325)
		);
	notech_reg opz1_reg_1(.CP(n_63097), .D(n_40331), .CD(n_62503), .Q(opz1[1
		]));
	notech_mux2 i_44130(.S(n_59338), .A(opz1[1]), .B(n_43629), .Z(n_40331)
		);
	notech_ao4 i_134379318(.A(n_60110), .B(n_44467), .C(n_1912), .D(n_43399)
		, .Z(n_188198993));
	notech_reg_set opz1_reg_2(.CP(n_63101), .D(n_40337), .SD(n_62503), .Q(opz1
		[2]));
	notech_mux2 i_44138(.S(n_59338), .A(opz1[2]), .B(n_2906), .Z(n_40337));
	notech_reg_set inst_deco_reg_0(.CP(n_63101), .D(n_40343), .SD(n_62503), 
		.Q(inst_deco[0]));
	notech_mux2 i_44146(.S(n_60143), .A(n_3465), .B(inst_deco[0]), .Z(n_40343
		));
	notech_ao4 i_134579316(.A(n_60110), .B(n_44468), .C(n_1912), .D(n_43401)
		, .Z(n_1877));
	notech_reg_set inst_deco_reg_1(.CP(n_63101), .D(n_40349), .SD(n_62499), 
		.Q(inst_deco[1]));
	notech_mux2 i_44154(.S(n_60143), .A(n_3464), .B(inst_deco[1]), .Z(n_40349
		));
	notech_reg_set inst_deco_reg_2(.CP(n_63101), .D(n_40355), .SD(n_62499), 
		.Q(inst_deco[2]));
	notech_mux2 i_44162(.S(n_60143), .A(n_3463), .B(inst_deco[2]), .Z(n_40355
		));
	notech_ao4 i_134779314(.A(n_60110), .B(n_44469), .C(n_1912), .D(n_43403)
		, .Z(n_1875));
	notech_reg_set inst_deco_reg_3(.CP(n_63101), .D(n_40361), .SD(n_62503), 
		.Q(inst_deco[3]));
	notech_mux2 i_44170(.S(n_60143), .A(n_3462), .B(inst_deco[3]), .Z(n_40361
		));
	notech_reg_set inst_deco_reg_4(.CP(n_63133), .D(n_40367), .SD(n_62503), 
		.Q(inst_deco[4]));
	notech_mux2 i_44178(.S(n_60143), .A(n_3461), .B(inst_deco[4]), .Z(n_40367
		));
	notech_ao4 i_134979312(.A(n_60110), .B(n_44470), .C(n_1912), .D(n_43405)
		, .Z(n_1873));
	notech_reg_set inst_deco_reg_5(.CP(n_63168), .D(n_40373), .SD(n_62503), 
		.Q(inst_deco[5]));
	notech_mux2 i_44186(.S(n_60143), .A(n_3460), .B(inst_deco[5]), .Z(n_40373
		));
	notech_reg_set inst_deco_reg_6(.CP(n_63168), .D(n_40379), .SD(n_62503), 
		.Q(inst_deco[6]));
	notech_mux2 i_44194(.S(n_60143), .A(n_3459), .B(inst_deco[6]), .Z(n_40379
		));
	notech_ao4 i_135179310(.A(n_60110), .B(n_44472), .C(n_1912), .D(n_43406)
		, .Z(n_1871));
	notech_reg_set inst_deco_reg_7(.CP(n_63168), .D(n_40385), .SD(n_62503), 
		.Q(inst_deco[7]));
	notech_mux2 i_44202(.S(n_60143), .A(n_3458), .B(inst_deco[7]), .Z(n_40385
		));
	notech_reg_set inst_deco_reg_8(.CP(n_63168), .D(n_40391), .SD(n_62570), 
		.Q(inst_deco[8]));
	notech_mux2 i_44210(.S(n_60143), .A(n_44817), .B(inst_deco[8]), .Z(n_40391
		));
	notech_ao4 i_135379308(.A(n_60110), .B(n_44473), .C(n_1912), .D(n_43409)
		, .Z(n_1869));
	notech_reg_set inst_deco_reg_9(.CP(n_63168), .D(n_40397), .SD(n_62570), 
		.Q(inst_deco[9]));
	notech_mux2 i_44218(.S(n_60143), .A(n_44823), .B(inst_deco[9]), .Z(n_40397
		));
	notech_reg_set inst_deco_reg_10(.CP(n_63168), .D(n_40403), .SD(n_62570),
		 .Q(inst_deco[10]));
	notech_mux2 i_44226(.S(n_60143), .A(n_44829), .B(inst_deco[10]), .Z(n_40403
		));
	notech_ao4 i_135579306(.A(n_60110), .B(n_44474), .C(n_1912), .D(n_43410)
		, .Z(n_1867));
	notech_reg_set inst_deco_reg_11(.CP(n_63168), .D(n_40409), .SD(n_62570),
		 .Q(inst_deco[11]));
	notech_mux2 i_44234(.S(n_60143), .A(n_44835), .B(inst_deco[11]), .Z(n_40409
		));
	notech_reg_set inst_deco_reg_12(.CP(n_63168), .D(n_40415), .SD(n_62570),
		 .Q(inst_deco[12]));
	notech_mux2 i_44242(.S(n_60143), .A(n_44841), .B(inst_deco[12]), .Z(n_40415
		));
	notech_ao4 i_135779304(.A(n_60110), .B(n_44475), .C(n_1912), .D(n_43412)
		, .Z(n_1865));
	notech_reg_set inst_deco_reg_13(.CP(n_63168), .D(n_40421), .SD(n_62570),
		 .Q(inst_deco[13]));
	notech_mux2 i_44250(.S(n_60143), .A(n_44847), .B(inst_deco[13]), .Z(n_40421
		));
	notech_ao4 i_135879303(.A(n_59138), .B(n_43283), .C(n_60110), .D(n_44476
		), .Z(n_1864));
	notech_reg_set inst_deco_reg_14(.CP(n_63168), .D(n_40427), .SD(n_62570),
		 .Q(inst_deco[14]));
	notech_mux2 i_44258(.S(n_60143), .A(n_44853), .B(inst_deco[14]), .Z(n_40427
		));
	notech_ao4 i_135979302(.A(n_59138), .B(n_43285), .C(n_60110), .D(n_44478
		), .Z(n_1863));
	notech_reg_set inst_deco_reg_15(.CP(n_63168), .D(n_40433), .SD(n_62570),
		 .Q(inst_deco[15]));
	notech_mux2 i_44266(.S(n_60143), .A(n_3457), .B(inst_deco[15]), .Z(n_40433
		));
	notech_ao4 i_136079301(.A(n_59139), .B(n_43287), .C(n_60110), .D(n_44479
		), .Z(n_1862));
	notech_reg_set inst_deco_reg_16(.CP(n_63166), .D(n_40439), .SD(n_62570),
		 .Q(inst_deco[16]));
	notech_mux2 i_44274(.S(n_60141), .A(n_44865), .B(inst_deco[16]), .Z(n_40439
		));
	notech_ao4 i_136179300(.A(n_59139), .B(n_43290), .C(n_60110), .D(n_44480
		), .Z(n_1861));
	notech_reg_set inst_deco_reg_17(.CP(n_63168), .D(n_40445), .SD(n_62570),
		 .Q(inst_deco[17]));
	notech_mux2 i_44282(.S(n_60141), .A(n_2913), .B(inst_deco[17]), .Z(n_40445
		));
	notech_ao4 i_136279299(.A(n_59139), .B(n_43292), .C(n_60110), .D(n_44481
		), .Z(n_1860));
	notech_reg_set inst_deco_reg_18(.CP(n_63166), .D(n_40451), .SD(n_62570),
		 .Q(inst_deco[18]));
	notech_mux2 i_44290(.S(n_60141), .A(n_44877), .B(inst_deco[18]), .Z(n_40451
		));
	notech_ao4 i_136379298(.A(n_59139), .B(n_43295), .C(n_60110), .D(n_44482
		), .Z(n_1859));
	notech_reg_set inst_deco_reg_19(.CP(n_63166), .D(n_40457), .SD(n_62568),
		 .Q(inst_deco[19]));
	notech_mux2 i_44298(.S(n_60141), .A(n_44883), .B(inst_deco[19]), .Z(n_40457
		));
	notech_ao4 i_136479297(.A(n_59139), .B(n_43297), .C(n_60110), .D(n_44484
		), .Z(n_1858));
	notech_reg_set inst_deco_reg_20(.CP(n_63166), .D(n_40463), .SD(n_62568),
		 .Q(inst_deco[20]));
	notech_mux2 i_44306(.S(n_60141), .A(n_3456), .B(inst_deco[20]), .Z(n_40463
		));
	notech_ao4 i_136579296(.A(n_59139), .B(n_43299), .C(n_60110), .D(n_44485
		), .Z(n_1857));
	notech_reg_set inst_deco_reg_21(.CP(n_63168), .D(n_40469), .SD(n_62568),
		 .Q(inst_deco[21]));
	notech_mux2 i_44314(.S(n_60141), .A(n_2909), .B(inst_deco[21]), .Z(n_40469
		));
	notech_ao4 i_136679295(.A(n_59139), .B(n_43302), .C(n_60117), .D(n_44486
		), .Z(n_1856));
	notech_reg_set inst_deco_reg_22(.CP(n_63168), .D(n_40475), .SD(n_62568),
		 .Q(inst_deco[22]));
	notech_mux2 i_44322(.S(n_60141), .A(n_44901), .B(inst_deco[22]), .Z(n_40475
		));
	notech_ao4 i_136779294(.A(n_59144), .B(n_43304), .C(n_60117), .D(n_44487
		), .Z(n_1855));
	notech_reg_set inst_deco_reg_23(.CP(n_63168), .D(n_40481), .SD(n_62568),
		 .Q(inst_deco[23]));
	notech_mux2 i_44330(.S(n_60141), .A(n_44907), .B(inst_deco[23]), .Z(n_40481
		));
	notech_ao4 i_136879293(.A(n_59144), .B(n_43307), .C(n_60117), .D(n_44488
		), .Z(n_1854));
	notech_reg_set inst_deco_reg_24(.CP(n_63168), .D(n_40487), .SD(n_62570),
		 .Q(inst_deco[24]));
	notech_mux2 i_44338(.S(n_60141), .A(n_3455), .B(inst_deco[24]), .Z(n_40487
		));
	notech_ao4 i_136979292(.A(n_59144), .B(n_43309), .C(n_60117), .D(n_44490
		), .Z(n_1853));
	notech_reg_set inst_deco_reg_25(.CP(n_63168), .D(n_40493), .SD(n_62570),
		 .Q(inst_deco[25]));
	notech_mux2 i_44346(.S(n_60141), .A(n_3454), .B(inst_deco[25]), .Z(n_40493
		));
	notech_ao4 i_137079291(.A(n_59144), .B(n_43311), .C(n_60117), .D(n_44491
		), .Z(n_1852));
	notech_reg_set inst_deco_reg_26(.CP(n_63171), .D(n_40499), .SD(n_62570),
		 .Q(inst_deco[26]));
	notech_mux2 i_44354(.S(n_60141), .A(n_3453), .B(inst_deco[26]), .Z(n_40499
		));
	notech_ao4 i_137179290(.A(n_59144), .B(n_43314), .C(n_60117), .D(n_44492
		), .Z(n_1851));
	notech_reg_set inst_deco_reg_27(.CP(n_63171), .D(n_40505), .SD(n_62570),
		 .Q(inst_deco[27]));
	notech_mux2 i_44362(.S(n_60141), .A(n_3452), .B(inst_deco[27]), .Z(n_40505
		));
	notech_ao4 i_137279289(.A(n_59144), .B(n_43316), .C(n_60117), .D(n_44493
		), .Z(n_1850));
	notech_reg_set inst_deco_reg_28(.CP(n_63171), .D(n_40511), .SD(n_62570),
		 .Q(inst_deco[28]));
	notech_mux2 i_44370(.S(n_60141), .A(n_3451), .B(inst_deco[28]), .Z(n_40511
		));
	notech_ao4 i_137379288(.A(n_59144), .B(n_43319), .C(n_60117), .D(n_44494
		), .Z(n_1849));
	notech_reg_set inst_deco_reg_29(.CP(n_63171), .D(n_40517), .SD(n_62573),
		 .Q(inst_deco[29]));
	notech_mux2 i_44378(.S(n_60141), .A(n_3450), .B(inst_deco[29]), .Z(n_40517
		));
	notech_ao4 i_137479287(.A(n_59146), .B(n_43321), .C(n_60117), .D(n_44496
		), .Z(n_1848));
	notech_reg_set inst_deco_reg_30(.CP(n_63171), .D(n_40523), .SD(n_62573),
		 .Q(inst_deco[30]));
	notech_mux2 i_44386(.S(n_60141), .A(n_3449), .B(inst_deco[30]), .Z(n_40523
		));
	notech_ao4 i_137579286(.A(n_59146), .B(n_43323), .C(n_60117), .D(n_44497
		), .Z(n_1847));
	notech_reg_set inst_deco_reg_31(.CP(n_63173), .D(n_40529), .SD(n_62573),
		 .Q(inst_deco[31]));
	notech_mux2 i_44394(.S(n_60141), .A(n_44955), .B(inst_deco[31]), .Z(n_40529
		));
	notech_reg_set inst_deco_reg_32(.CP(n_63173), .D(n_40535), .SD(n_62573),
		 .Q(inst_deco[32]));
	notech_mux2 i_44402(.S(n_60148), .A(n_3448), .B(inst_deco[32]), .Z(n_40535
		));
	notech_ao4 i_137779284(.A(n_60117), .B(n_44498), .C(n_42555), .D(n_44744
		), .Z(n_1845));
	notech_reg_set inst_deco_reg_33(.CP(n_63171), .D(n_40541), .SD(n_62573),
		 .Q(inst_deco[33]));
	notech_mux2 i_44410(.S(n_60148), .A(n_44967), .B(inst_deco[33]), .Z(n_40541
		));
	notech_ao4 i_137879283(.A(n_59146), .B(n_43327), .C(n_60117), .D(n_44499
		), .Z(n_1844));
	notech_reg_set inst_deco_reg_34(.CP(n_63171), .D(n_40547), .SD(n_62573),
		 .Q(inst_deco[34]));
	notech_mux2 i_44418(.S(n_60148), .A(n_44973), .B(inst_deco[34]), .Z(n_40547
		));
	notech_ao4 i_137979282(.A(n_59146), .B(n_43329), .C(n_60117), .D(n_44500
		), .Z(n_1843));
	notech_reg_set inst_deco_reg_35(.CP(n_63171), .D(n_40553), .SD(n_62575),
		 .Q(inst_deco[35]));
	notech_mux2 i_44426(.S(n_60148), .A(n_44979), .B(inst_deco[35]), .Z(n_40553
		));
	notech_ao4 i_138079281(.A(n_59144), .B(n_43332), .C(n_60117), .D(n_44501
		), .Z(n_1842));
	notech_reg_set inst_deco_reg_36(.CP(n_63171), .D(n_40559), .SD(n_62573),
		 .Q(inst_deco[36]));
	notech_mux2 i_44434(.S(n_60148), .A(n_44985), .B(inst_deco[36]), .Z(n_40559
		));
	notech_ao4 i_138179280(.A(n_59144), .B(n_43334), .C(n_60117), .D(n_44502
		), .Z(n_1841));
	notech_reg_set inst_deco_reg_37(.CP(n_63171), .D(n_40565), .SD(n_62573),
		 .Q(inst_deco[37]));
	notech_mux2 i_44442(.S(n_60148), .A(n_3447), .B(inst_deco[37]), .Z(n_40565
		));
	notech_ao4 i_138279279(.A(n_59146), .B(n_43337), .C(n_60117), .D(n_44503
		), .Z(n_1840));
	notech_reg_set inst_deco_reg_38(.CP(n_63171), .D(n_40571), .SD(n_62573),
		 .Q(inst_deco[38]));
	notech_mux2 i_44450(.S(n_60148), .A(n_44997), .B(inst_deco[38]), .Z(n_40571
		));
	notech_reg_set inst_deco_reg_39(.CP(n_63171), .D(n_40577), .SD(n_62573),
		 .Q(inst_deco[39]));
	notech_mux2 i_44458(.S(n_60148), .A(n_45003), .B(inst_deco[39]), .Z(n_40577
		));
	notech_ao4 i_138479277(.A(n_59144), .B(n_43339), .C(n_60115), .D(n_44504
		), .Z(n_1838));
	notech_reg_set inst_deco_reg_40(.CP(n_63168), .D(n_40583), .SD(n_62573),
		 .Q(inst_deco[40]));
	notech_mux2 i_44466(.S(n_60148), .A(n_45009), .B(inst_deco[40]), .Z(n_40583
		));
	notech_mux2 i_10980631(.S(pg_fault), .A(n_60854), .B(n_160356214), .Z(n_12254735
		));
	notech_reg_set inst_deco_reg_41(.CP(n_63171), .D(n_40589), .SD(n_62573),
		 .Q(inst_deco[41]));
	notech_mux2 i_44474(.S(n_60148), .A(n_45015), .B(inst_deco[41]), .Z(n_40589
		));
	notech_ao4 i_138779274(.A(n_59141), .B(n_43343), .C(n_60115), .D(n_44506
		), .Z(n_1837));
	notech_reg_set inst_deco_reg_42(.CP(n_63171), .D(n_40595), .SD(n_62573),
		 .Q(inst_deco[42]));
	notech_mux2 i_44482(.S(n_60148), .A(n_45021), .B(inst_deco[42]), .Z(n_40595
		));
	notech_reg_set inst_deco_reg_43(.CP(n_63171), .D(n_40601), .SD(n_62570),
		 .Q(inst_deco[43]));
	notech_mux2 i_44490(.S(n_60148), .A(n_3446), .B(inst_deco[43]), .Z(n_40601
		));
	notech_ao4 i_138879273(.A(n_59141), .B(n_43345), .C(n_60115), .D(n_44508
		), .Z(n_1835));
	notech_reg_set inst_deco_reg_44(.CP(n_63171), .D(n_40607), .SD(n_62570),
		 .Q(inst_deco[44]));
	notech_mux2 i_44498(.S(n_60148), .A(n_45033), .B(inst_deco[44]), .Z(n_40607
		));
	notech_ao4 i_138979272(.A(n_59141), .B(n_43347), .C(n_60115), .D(n_44509
		), .Z(n_1834));
	notech_reg_set inst_deco_reg_45(.CP(n_63171), .D(n_40613), .SD(n_62573),
		 .Q(inst_deco[45]));
	notech_mux2 i_44506(.S(n_60148), .A(n_45039), .B(inst_deco[45]), .Z(n_40613
		));
	notech_ao4 i_139079271(.A(n_59141), .B(n_43350), .C(n_60115), .D(n_44510
		), .Z(n_1833));
	notech_reg_set inst_deco_reg_46(.CP(n_63171), .D(n_40619), .SD(n_62573),
		 .Q(inst_deco[46]));
	notech_mux2 i_44514(.S(n_60148), .A(n_3445), .B(inst_deco[46]), .Z(n_40619
		));
	notech_ao4 i_139179270(.A(n_59141), .B(n_43352), .C(n_60115), .D(n_44511
		), .Z(n_1832));
	notech_reg_set inst_deco_reg_47(.CP(n_63166), .D(n_40625), .SD(n_62573),
		 .Q(inst_deco[47]));
	notech_mux2 i_44522(.S(n_60148), .A(n_3444), .B(inst_deco[47]), .Z(n_40625
		));
	notech_ao4 i_139279269(.A(n_59141), .B(n_43355), .C(n_60115), .D(n_44512
		), .Z(n_1831));
	notech_reg_set inst_deco_reg_48(.CP(n_63162), .D(n_40631), .SD(n_62573),
		 .Q(inst_deco[48]));
	notech_mux2 i_44530(.S(n_60146), .A(n_45057), .B(inst_deco[48]), .Z(n_40631
		));
	notech_ao4 i_139379268(.A(n_59141), .B(n_43357), .C(n_60115), .D(n_44514
		), .Z(n_1830));
	notech_reg_set inst_deco_reg_49(.CP(n_63162), .D(n_40637), .SD(n_62573),
		 .Q(inst_deco[49]));
	notech_mux2 i_44538(.S(n_60146), .A(n_45063), .B(inst_deco[49]), .Z(n_40637
		));
	notech_ao4 i_139479267(.A(n_59144), .B(n_43359), .C(n_60115), .D(n_44515
		), .Z(n_1829));
	notech_reg_set inst_deco_reg_50(.CP(n_63162), .D(n_40643), .SD(n_62564),
		 .Q(inst_deco[50]));
	notech_mux2 i_44546(.S(n_60146), .A(n_3443), .B(inst_deco[50]), .Z(n_40643
		));
	notech_ao4 i_139579266(.A(n_59144), .B(n_43362), .C(n_60115), .D(n_44516
		), .Z(n_1828));
	notech_reg_set inst_deco_reg_51(.CP(n_63162), .D(n_40649), .SD(n_62564),
		 .Q(inst_deco[51]));
	notech_mux2 i_44554(.S(n_60146), .A(n_45075), .B(inst_deco[51]), .Z(n_40649
		));
	notech_ao4 i_139679265(.A(n_59144), .B(n_43364), .C(n_60115), .D(n_44517
		), .Z(n_1827));
	notech_reg_set inst_deco_reg_52(.CP(n_63162), .D(n_40655), .SD(n_62564),
		 .Q(inst_deco[52]));
	notech_mux2 i_44562(.S(n_60146), .A(n_45081), .B(inst_deco[52]), .Z(n_40655
		));
	notech_ao4 i_139779264(.A(n_59144), .B(n_43367), .C(n_60115), .D(n_44518
		), .Z(n_1826));
	notech_reg_set inst_deco_reg_53(.CP(n_63162), .D(n_40661), .SD(n_62564),
		 .Q(inst_deco[53]));
	notech_mux2 i_44570(.S(n_60146), .A(n_45087), .B(inst_deco[53]), .Z(n_40661
		));
	notech_ao4 i_139879263(.A(n_59141), .B(n_43369), .C(n_60115), .D(n_44520
		), .Z(n_1825));
	notech_reg_set inst_deco_reg_54(.CP(n_63162), .D(n_40667), .SD(n_62564),
		 .Q(inst_deco[54]));
	notech_mux2 i_44578(.S(n_60146), .A(n_45093), .B(inst_deco[54]), .Z(n_40667
		));
	notech_ao4 i_139979262(.A(n_59144), .B(n_43371), .C(n_60115), .D(n_44521
		), .Z(n_1824));
	notech_reg_set inst_deco_reg_55(.CP(n_63162), .D(n_40673), .SD(n_62564),
		 .Q(inst_deco[55]));
	notech_mux2 i_44586(.S(n_60146), .A(n_3442), .B(inst_deco[55]), .Z(n_40673
		));
	notech_reg_set inst_deco_reg_56(.CP(n_63162), .D(n_40679), .SD(n_62564),
		 .Q(inst_deco[56]));
	notech_mux2 i_44594(.S(n_60146), .A(n_45105), .B(inst_deco[56]), .Z(n_40679
		));
	notech_ao4 i_140079261(.A(n_59144), .B(n_43374), .C(n_60115), .D(n_44522
		), .Z(n_1823));
	notech_reg_set inst_deco_reg_57(.CP(n_63162), .D(n_40685), .SD(n_62564),
		 .Q(inst_deco[57]));
	notech_mux2 i_44602(.S(n_60146), .A(n_45111), .B(inst_deco[57]), .Z(n_40685
		));
	notech_reg_set inst_deco_reg_58(.CP(n_63160), .D(n_40691), .SD(n_62564),
		 .Q(inst_deco[58]));
	notech_mux2 i_44610(.S(n_60146), .A(n_3441), .B(inst_deco[58]), .Z(n_40691
		));
	notech_reg_set inst_deco_reg_59(.CP(n_63160), .D(n_40697), .SD(n_62564),
		 .Q(inst_deco[59]));
	notech_mux2 i_44618(.S(n_60146), .A(n_45123), .B(inst_deco[59]), .Z(n_40697
		));
	notech_reg_set inst_deco_reg_60(.CP(n_63160), .D(n_40703), .SD(n_62562),
		 .Q(inst_deco[60]));
	notech_mux2 i_44626(.S(n_60146), .A(n_45129), .B(inst_deco[60]), .Z(n_40703
		));
	notech_reg_set inst_deco_reg_61(.CP(n_63160), .D(n_40709), .SD(n_62562),
		 .Q(inst_deco[61]));
	notech_mux2 i_44634(.S(n_60146), .A(n_45135), .B(inst_deco[61]), .Z(n_40709
		));
	notech_reg_set inst_deco_reg_62(.CP(n_63160), .D(n_40715), .SD(n_62562),
		 .Q(inst_deco[62]));
	notech_mux2 i_44642(.S(n_60146), .A(n_45141), .B(inst_deco[62]), .Z(n_40715
		));
	notech_reg_set inst_deco_reg_63(.CP(n_63160), .D(n_40721), .SD(n_62562),
		 .Q(inst_deco[63]));
	notech_mux2 i_44650(.S(n_60146), .A(n_45147), .B(inst_deco[63]), .Z(n_40721
		));
	notech_and4 i_142679235(.A(n_60937), .B(n_60115), .C(n_2384), .D(n_44200
		), .Z(n_1817));
	notech_reg_set inst_deco_reg_64(.CP(n_63160), .D(n_40727), .SD(n_62562),
		 .Q(inst_deco[64]));
	notech_mux2 i_44658(.S(n_60133), .A(n_45153), .B(inst_deco[64]), .Z(n_40727
		));
	notech_reg_set inst_deco_reg_65(.CP(n_63160), .D(n_40733), .SD(n_62562),
		 .Q(inst_deco[65]));
	notech_mux2 i_44666(.S(n_60133), .A(n_3440), .B(inst_deco[65]), .Z(n_40733
		));
	notech_reg_set inst_deco_reg_66(.CP(n_63160), .D(n_40739), .SD(n_62562),
		 .Q(inst_deco[66]));
	notech_mux2 i_44674(.S(n_60133), .A(n_3439), .B(inst_deco[66]), .Z(n_40739
		));
	notech_reg_set inst_deco_reg_67(.CP(n_63160), .D(n_40745), .SD(n_62562),
		 .Q(inst_deco[67]));
	notech_mux2 i_44682(.S(n_60133), .A(n_3438), .B(inst_deco[67]), .Z(n_40745
		));
	notech_ao4 i_9880632(.A(n_42549), .B(n_2402), .C(n_42724), .D(n_44170), 
		.Z(n_1813));
	notech_reg_set inst_deco_reg_68(.CP(n_63160), .D(n_40751), .SD(n_62562),
		 .Q(inst_deco[68]));
	notech_mux2 i_44690(.S(n_60133), .A(n_3437), .B(inst_deco[68]), .Z(n_40751
		));
	notech_ao4 i_142879233(.A(n_42549), .B(n_44169), .C(n_2336), .D(n_1811),
		 .Z(n_1812));
	notech_reg_set inst_deco_reg_69(.CP(n_63166), .D(n_40757), .SD(n_62562),
		 .Q(inst_deco[69]));
	notech_mux2 i_44698(.S(n_60133), .A(n_3436), .B(inst_deco[69]), .Z(n_40757
		));
	notech_or4 i_143079231(.A(ipg_fault), .B(n_57724), .C(n_2997), .D(n_44170
		), .Z(n_1811));
	notech_reg_set inst_deco_reg_70(.CP(n_63166), .D(n_40763), .SD(n_62562),
		 .Q(inst_deco[70]));
	notech_mux2 i_44706(.S(n_60133), .A(n_3435), .B(inst_deco[70]), .Z(n_40763
		));
	notech_reg_set inst_deco_reg_71(.CP(n_63166), .D(n_40769), .SD(n_62568),
		 .Q(inst_deco[71]));
	notech_mux2 i_44714(.S(n_60133), .A(n_3434), .B(inst_deco[71]), .Z(n_40769
		));
	notech_reg_set inst_deco_reg_72(.CP(n_63166), .D(n_40775), .SD(n_62568),
		 .Q(inst_deco[72]));
	notech_mux2 i_44722(.S(n_60133), .A(n_3433), .B(inst_deco[72]), .Z(n_40775
		));
	notech_reg_set inst_deco_reg_73(.CP(n_63166), .D(n_40781), .SD(n_62568),
		 .Q(inst_deco[73]));
	notech_mux2 i_44730(.S(n_60133), .A(n_3432), .B(inst_deco[73]), .Z(n_40781
		));
	notech_reg_set inst_deco_reg_74(.CP(n_63166), .D(n_40787), .SD(n_62568),
		 .Q(inst_deco[74]));
	notech_mux2 i_44738(.S(n_60133), .A(n_45213), .B(inst_deco[74]), .Z(n_40787
		));
	notech_reg_set inst_deco_reg_75(.CP(n_63166), .D(n_40793), .SD(n_62568),
		 .Q(inst_deco[75]));
	notech_mux2 i_44746(.S(n_60133), .A(n_3431), .B(inst_deco[75]), .Z(n_40793
		));
	notech_reg_set inst_deco_reg_76(.CP(n_63166), .D(n_40799), .SD(n_62568),
		 .Q(inst_deco[76]));
	notech_mux2 i_44754(.S(n_60133), .A(n_3430), .B(inst_deco[76]), .Z(n_40799
		));
	notech_and4 i_125679405(.A(n_2379), .B(db67), .C(\fpu_indrm[0] ), .D(fpu
		), .Z(n_1804));
	notech_reg_set inst_deco_reg_77(.CP(n_63166), .D(n_40805), .SD(n_62568),
		 .Q(inst_deco[77]));
	notech_mux2 i_44762(.S(n_60133), .A(n_3429), .B(inst_deco[77]), .Z(n_40805
		));
	notech_and4 i_125579406(.A(n_2859), .B(db67), .C(n_5712), .D(n_2942), .Z
		(n_1803));
	notech_reg_set inst_deco_reg_78(.CP(n_63166), .D(n_40811), .SD(n_62568),
		 .Q(inst_deco[78]));
	notech_mux2 i_44770(.S(n_60133), .A(n_3428), .B(inst_deco[78]), .Z(n_40811
		));
	notech_reg_set inst_deco_reg_79(.CP(n_63166), .D(n_40817), .SD(n_62568),
		 .Q(inst_deco[79]));
	notech_mux2 i_44778(.S(n_60133), .A(n_3427), .B(inst_deco[79]), .Z(n_40817
		));
	notech_reg_set inst_deco_reg_80(.CP(n_63162), .D(n_40823), .SD(n_62568),
		 .Q(inst_deco[80]));
	notech_mux2 i_44786(.S(n_60131), .A(n_3426), .B(inst_deco[80]), .Z(n_40823
		));
	notech_nao3 i_125179410(.A(ipg_fault), .B(n_2995), .C(n_57724), .Z(n_1800
		));
	notech_reg_set inst_deco_reg_81(.CP(n_63162), .D(n_40829), .SD(n_62568),
		 .Q(inst_deco[81]));
	notech_mux2 i_44794(.S(n_60131), .A(n_3425), .B(inst_deco[81]), .Z(n_40829
		));
	notech_ao3 i_2786(.A(n_2395), .B(n_1599), .C(n_2981), .Z(useq_ptr[3]));
	notech_reg_set inst_deco_reg_82(.CP(n_63162), .D(n_40835), .SD(n_62564),
		 .Q(inst_deco[82]));
	notech_mux2 i_44802(.S(n_60131), .A(n_3424), .B(inst_deco[82]), .Z(n_40835
		));
	notech_and3 i_2787(.A(n_2395), .B(n_1599), .C(n_2983), .Z(useq_ptr[2])
		);
	notech_reg_set inst_deco_reg_83(.CP(n_63162), .D(n_40841), .SD(n_62564),
		 .Q(inst_deco[83]));
	notech_mux2 i_44810(.S(n_60131), .A(n_3423), .B(inst_deco[83]), .Z(n_40841
		));
	notech_and3 i_2788(.A(n_2395), .B(n_1599), .C(n_2985), .Z(useq_ptr[1])
		);
	notech_reg_set inst_deco_reg_84(.CP(n_63162), .D(n_40847), .SD(n_62564),
		 .Q(inst_deco[84]));
	notech_mux2 i_44818(.S(n_60131), .A(n_3422), .B(inst_deco[84]), .Z(n_40847
		));
	notech_and3 i_2789(.A(n_2395), .B(n_1599), .C(n_2358), .Z(useq_ptr[0])
		);
	notech_reg_set inst_deco_reg_85(.CP(n_63166), .D(n_40853), .SD(n_62564),
		 .Q(inst_deco[85]));
	notech_mux2 i_44826(.S(n_60131), .A(n_3421), .B(inst_deco[85]), .Z(n_40853
		));
	notech_reg_set inst_deco_reg_86(.CP(n_63166), .D(n_40859), .SD(n_62564),
		 .Q(inst_deco[86]));
	notech_mux2 i_44834(.S(n_60131), .A(n_3420), .B(inst_deco[86]), .Z(n_40859
		));
	notech_reg_set inst_deco_reg_87(.CP(n_63162), .D(n_40865), .SD(n_62568),
		 .Q(inst_deco[87]));
	notech_mux2 i_44842(.S(n_60131), .A(n_3419), .B(inst_deco[87]), .Z(n_40865
		));
	notech_reg_set inst_deco_reg_88(.CP(n_63162), .D(n_40871), .SD(n_62568),
		 .Q(inst_deco[88]));
	notech_mux2 i_44850(.S(n_60131), .A(n_3418), .B(inst_deco[88]), .Z(n_40871
		));
	notech_reg_set inst_deco_reg_89(.CP(n_63162), .D(n_40877), .SD(n_62564),
		 .Q(inst_deco[89]));
	notech_mux2 i_44858(.S(n_60131), .A(n_3417), .B(inst_deco[89]), .Z(n_40877
		));
	notech_reg_set inst_deco_reg_90(.CP(n_63182), .D(n_40883), .SD(n_62564),
		 .Q(inst_deco[90]));
	notech_mux2 i_44866(.S(n_60131), .A(n_3416), .B(inst_deco[90]), .Z(n_40883
		));
	notech_reg_set inst_deco_reg_91(.CP(n_63182), .D(n_40889), .SD(n_62564),
		 .Q(inst_deco[91]));
	notech_mux2 i_44874(.S(n_60131), .A(n_3415), .B(inst_deco[91]), .Z(n_40889
		));
	notech_reg_set inst_deco_reg_92(.CP(n_63182), .D(n_40895), .SD(n_62575),
		 .Q(inst_deco[92]));
	notech_mux2 i_44882(.S(n_60131), .A(n_3414), .B(inst_deco[92]), .Z(n_40895
		));
	notech_reg_set inst_deco_reg_93(.CP(n_63182), .D(n_40901), .SD(n_62584),
		 .Q(inst_deco[93]));
	notech_mux2 i_44890(.S(n_60131), .A(n_3413), .B(inst_deco[93]), .Z(n_40901
		));
	notech_reg_set inst_deco_reg_94(.CP(n_63182), .D(n_40907), .SD(n_62584),
		 .Q(inst_deco[94]));
	notech_mux2 i_44898(.S(n_60131), .A(n_3412), .B(inst_deco[94]), .Z(n_40907
		));
	notech_reg_set inst_deco_reg_95(.CP(n_63182), .D(n_40913), .SD(n_62584),
		 .Q(inst_deco[95]));
	notech_mux2 i_44906(.S(n_60131), .A(n_3411), .B(inst_deco[95]), .Z(n_40913
		));
	notech_reg_set inst_deco_reg_96(.CP(n_63182), .D(n_40919), .SD(n_62584),
		 .Q(inst_deco[96]));
	notech_mux2 i_44914(.S(n_60138), .A(n_3410), .B(inst_deco[96]), .Z(n_40919
		));
	notech_reg_set inst_deco_reg_97(.CP(n_63182), .D(n_40925), .SD(n_62584),
		 .Q(inst_deco[97]));
	notech_mux2 i_44922(.S(n_60138), .A(n_3409), .B(inst_deco[97]), .Z(n_40925
		));
	notech_reg_set inst_deco_reg_98(.CP(n_63182), .D(n_40931), .SD(n_62584),
		 .Q(inst_deco[98]));
	notech_mux2 i_44930(.S(n_60138), .A(n_3408), .B(inst_deco[98]), .Z(n_40931
		));
	notech_reg_set inst_deco_reg_99(.CP(n_63182), .D(n_40937), .SD(n_62584),
		 .Q(inst_deco[99]));
	notech_mux2 i_44938(.S(n_60138), .A(n_3407), .B(inst_deco[99]), .Z(n_40937
		));
	notech_reg_set inst_deco_reg_100(.CP(n_63182), .D(n_40943), .SD(n_62584)
		, .Q(inst_deco[100]));
	notech_mux2 i_44946(.S(n_60138), .A(n_3406), .B(inst_deco[100]), .Z(n_40943
		));
	notech_reg_set inst_deco_reg_101(.CP(n_63178), .D(n_40949), .SD(n_62584)
		, .Q(inst_deco[101]));
	notech_mux2 i_44954(.S(n_60138), .A(n_3405), .B(inst_deco[101]), .Z(n_40949
		));
	notech_reg_set inst_deco_reg_102(.CP(n_63178), .D(n_40955), .SD(n_62584)
		, .Q(inst_deco[102]));
	notech_mux2 i_44962(.S(n_60138), .A(n_3404), .B(inst_deco[102]), .Z(n_40955
		));
	notech_reg_set inst_deco_reg_103(.CP(n_63178), .D(n_40961), .SD(n_62584)
		, .Q(inst_deco[103]));
	notech_mux2 i_44970(.S(n_60138), .A(n_3403), .B(inst_deco[103]), .Z(n_40961
		));
	notech_reg_set inst_deco_reg_104(.CP(n_63178), .D(n_40967), .SD(n_62580)
		, .Q(inst_deco[104]));
	notech_mux2 i_44978(.S(n_60138), .A(n_3402), .B(inst_deco[104]), .Z(n_40967
		));
	notech_reg_set inst_deco_reg_105(.CP(n_63178), .D(n_40973), .SD(n_62580)
		, .Q(inst_deco[105]));
	notech_mux2 i_44986(.S(n_60138), .A(n_3401), .B(inst_deco[105]), .Z(n_40973
		));
	notech_reg_set inst_deco_reg_106(.CP(n_63178), .D(n_40979), .SD(n_62580)
		, .Q(inst_deco[106]));
	notech_mux2 i_44994(.S(n_60138), .A(n_3400), .B(inst_deco[106]), .Z(n_40979
		));
	notech_reg_set inst_deco_reg_107(.CP(n_63182), .D(n_40985), .SD(n_62580)
		, .Q(inst_deco[107]));
	notech_mux2 i_45002(.S(n_60138), .A(n_3399), .B(inst_deco[107]), .Z(n_40985
		));
	notech_reg_set inst_deco_reg_108(.CP(n_63178), .D(n_40991), .SD(n_62580)
		, .Q(inst_deco[108]));
	notech_mux2 i_45010(.S(n_60138), .A(n_3398), .B(inst_deco[108]), .Z(n_40991
		));
	notech_reg_set inst_deco_reg_109(.CP(n_63178), .D(n_40997), .SD(n_62580)
		, .Q(inst_deco[109]));
	notech_mux2 i_45018(.S(n_60138), .A(n_3397), .B(inst_deco[109]), .Z(n_40997
		));
	notech_reg_set inst_deco_reg_110(.CP(n_63178), .D(n_41003), .SD(n_62580)
		, .Q(inst_deco[110]));
	notech_mux2 i_45026(.S(n_60138), .A(n_3396), .B(inst_deco[110]), .Z(n_41003
		));
	notech_reg_set inst_deco_reg_111(.CP(n_63184), .D(n_41009), .SD(n_62580)
		, .Q(inst_deco[111]));
	notech_mux2 i_45034(.S(n_60138), .A(n_3395), .B(inst_deco[111]), .Z(n_41009
		));
	notech_reg_set inst_deco_reg_112(.CP(n_63184), .D(n_41015), .SD(n_62580)
		, .Q(inst_deco[112]));
	notech_mux2 i_45042(.S(n_60136), .A(n_3394), .B(inst_deco[112]), .Z(n_41015
		));
	notech_reg_set inst_deco_reg_113(.CP(n_63184), .D(n_41021), .SD(n_62580)
		, .Q(inst_deco[113]));
	notech_mux2 i_45050(.S(n_60136), .A(n_45447), .B(inst_deco[113]), .Z(n_41021
		));
	notech_reg_set inst_deco_reg_114(.CP(n_63184), .D(n_41027), .SD(n_62586)
		, .Q(inst_deco[114]));
	notech_mux2 i_45058(.S(n_60136), .A(n_3393), .B(inst_deco[114]), .Z(n_41027
		));
	notech_reg_set inst_deco_reg_115(.CP(n_63184), .D(n_41033), .SD(n_62586)
		, .Q(inst_deco[115]));
	notech_mux2 i_45066(.S(n_60136), .A(n_3392), .B(inst_deco[115]), .Z(n_41033
		));
	notech_reg_set inst_deco_reg_116(.CP(n_63184), .D(n_41039), .SD(n_62586)
		, .Q(inst_deco[116]));
	notech_mux2 i_45074(.S(n_60136), .A(n_3391), .B(inst_deco[116]), .Z(n_41039
		));
	notech_reg_set inst_deco_reg_117(.CP(n_63184), .D(n_41045), .SD(n_62586)
		, .Q(inst_deco[117]));
	notech_mux2 i_45082(.S(n_60136), .A(n_3390), .B(inst_deco[117]), .Z(n_41045
		));
	notech_reg_set inst_deco_reg_118(.CP(n_63184), .D(n_41051), .SD(n_62586)
		, .Q(inst_deco[118]));
	notech_mux2 i_45090(.S(n_60136), .A(n_3389), .B(inst_deco[118]), .Z(n_41051
		));
	notech_reg_set inst_deco_reg_119(.CP(n_63184), .D(n_41057), .SD(n_62586)
		, .Q(inst_deco[119]));
	notech_mux2 i_45098(.S(n_60136), .A(n_3388), .B(inst_deco[119]), .Z(n_41057
		));
	notech_reg_set inst_deco_reg_120(.CP(n_63184), .D(n_41063), .SD(n_62586)
		, .Q(inst_deco[120]));
	notech_mux2 i_45106(.S(n_60136), .A(n_3387), .B(inst_deco[120]), .Z(n_41063
		));
	notech_reg_set inst_deco_reg_121(.CP(n_63184), .D(n_41069), .SD(n_62586)
		, .Q(inst_deco[121]));
	notech_mux2 i_45114(.S(n_60136), .A(n_3386), .B(inst_deco[121]), .Z(n_41069
		));
	notech_reg_set inst_deco_reg_122(.CP(n_63182), .D(n_41075), .SD(n_62586)
		, .Q(inst_deco[122]));
	notech_mux2 i_45122(.S(n_60136), .A(n_3385), .B(inst_deco[122]), .Z(n_41075
		));
	notech_reg_set inst_deco_reg_123(.CP(n_63182), .D(n_41081), .SD(n_62586)
		, .Q(inst_deco[123]));
	notech_mux2 i_45130(.S(n_60136), .A(n_3384), .B(inst_deco[123]), .Z(n_41081
		));
	notech_reg_set inst_deco_reg_124(.CP(n_63182), .D(n_41087), .SD(n_62586)
		, .Q(inst_deco[124]));
	notech_mux2 i_45138(.S(n_60136), .A(n_3383), .B(inst_deco[124]), .Z(n_41087
		));
	notech_reg_set inst_deco_reg_125(.CP(n_63182), .D(n_41093), .SD(n_62584)
		, .Q(inst_deco[125]));
	notech_mux2 i_45146(.S(n_60136), .A(n_3382), .B(inst_deco[125]), .Z(n_41093
		));
	notech_reg_set inst_deco_reg_126(.CP(n_63182), .D(n_41099), .SD(n_62584)
		, .Q(inst_deco[126]));
	notech_mux2 i_45154(.S(n_60136), .A(n_3381), .B(inst_deco[126]), .Z(n_41099
		));
	notech_reg_set inst_deco_reg_127(.CP(n_63184), .D(n_41105), .SD(n_62584)
		, .Q(inst_deco[127]));
	notech_mux2 i_45162(.S(n_60136), .A(n_3380), .B(inst_deco[127]), .Z(n_41105
		));
	notech_nand3 i_26580391(.A(n_2995), .B(inst_deco1[106]), .C(n_59405), .Z
		(n_1757));
	notech_reg to_acu0_reg_0(.CP(n_63184), .D(n_41111), .CD(n_62584), .Q(to_acu0
		[0]));
	notech_mux2 i_45170(.S(n_56660), .A(n_42565), .B(to_acu0[0]), .Z(n_41111
		));
	notech_reg to_acu0_reg_1(.CP(n_63184), .D(n_41117), .CD(n_62584), .Q(to_acu0
		[1]));
	notech_mux2 i_45178(.S(n_56660), .A(n_42566), .B(to_acu0[1]), .Z(n_41117
		));
	notech_reg to_acu0_reg_2(.CP(n_63182), .D(n_41123), .CD(n_62586), .Q(to_acu0
		[2]));
	notech_mux2 i_45186(.S(n_56640), .A(n_42567), .B(to_acu0[2]), .Z(n_41123
		));
	notech_reg to_acu0_reg_3(.CP(n_63184), .D(n_41129), .CD(n_62586), .Q(to_acu0
		[3]));
	notech_mux2 i_45194(.S(n_56660), .A(n_42568), .B(to_acu0[3]), .Z(n_41129
		));
	notech_reg to_acu0_reg_4(.CP(n_63178), .D(n_41135), .CD(n_62586), .Q(to_acu0
		[4]));
	notech_mux2 i_45202(.S(n_56660), .A(n_42569), .B(to_acu0[4]), .Z(n_41135
		));
	notech_reg to_acu0_reg_5(.CP(n_63173), .D(n_41141), .CD(n_62584), .Q(to_acu0
		[5]));
	notech_mux2 i_45210(.S(n_56640), .A(n_42571), .B(to_acu0[5]), .Z(n_41141
		));
	notech_reg to_acu0_reg_6(.CP(n_63173), .D(n_41147), .CD(n_62584), .Q(to_acu0
		[6]));
	notech_mux2 i_45218(.S(n_56640), .A(n_42572), .B(to_acu0[6]), .Z(n_41147
		));
	notech_reg to_acu0_reg_7(.CP(n_63173), .D(n_41153), .CD(n_62575), .Q(to_acu0
		[7]));
	notech_mux2 i_45226(.S(n_56640), .A(n_44201), .B(to_acu0[7]), .Z(n_41153
		));
	notech_reg to_acu0_reg_8(.CP(n_63173), .D(n_41159), .CD(n_62575), .Q(to_acu0
		[8]));
	notech_mux2 i_45234(.S(n_56640), .A(n_44203), .B(to_acu0[8]), .Z(n_41159
		));
	notech_reg to_acu0_reg_9(.CP(n_63173), .D(n_41165), .CD(n_62575), .Q(to_acu0
		[9]));
	notech_mux2 i_45242(.S(n_56660), .A(n_44204), .B(to_acu0[9]), .Z(n_41165
		));
	notech_reg to_acu0_reg_10(.CP(n_63176), .D(n_41171), .CD(n_62575), .Q(to_acu0
		[10]));
	notech_mux2 i_45250(.S(n_56660), .A(n_44205), .B(to_acu0[10]), .Z(n_41171
		));
	notech_reg to_acu0_reg_11(.CP(n_63176), .D(n_41177), .CD(n_62575), .Q(to_acu0
		[11]));
	notech_mux2 i_45258(.S(n_56660), .A(n_44206), .B(to_acu0[11]), .Z(n_41177
		));
	notech_reg to_acu0_reg_12(.CP(n_63176), .D(n_41183), .CD(n_62578), .Q(to_acu0
		[12]));
	notech_mux2 i_45266(.S(n_56660), .A(n_44207), .B(to_acu0[12]), .Z(n_41183
		));
	notech_reg to_acu0_reg_13(.CP(n_63176), .D(n_41189), .CD(n_62578), .Q(to_acu0
		[13]));
	notech_mux2 i_45274(.S(n_56660), .A(n_44209), .B(to_acu0[13]), .Z(n_41189
		));
	notech_reg to_acu0_reg_14(.CP(n_63176), .D(n_41195), .CD(n_62578), .Q(to_acu0
		[14]));
	notech_mux2 i_45282(.S(n_56660), .A(n_44210), .B(to_acu0[14]), .Z(n_41195
		));
	notech_reg to_acu0_reg_15(.CP(n_63173), .D(n_41201), .CD(n_62578), .Q(to_acu0
		[15]));
	notech_mux2 i_45290(.S(n_56660), .A(n_44211), .B(to_acu0[15]), .Z(n_41201
		));
	notech_reg to_acu0_reg_16(.CP(n_63173), .D(n_41207), .CD(n_62578), .Q(to_acu0
		[16]));
	notech_mux2 i_45298(.S(n_56660), .A(n_44212), .B(to_acu0[16]), .Z(n_41207
		));
	notech_reg to_acu0_reg_17(.CP(n_63173), .D(n_41213), .CD(n_62575), .Q(to_acu0
		[17]));
	notech_mux2 i_45306(.S(n_56674), .A(n_44213), .B(to_acu0[17]), .Z(n_41213
		));
	notech_reg to_acu0_reg_18(.CP(n_63173), .D(n_41219), .CD(n_62575), .Q(to_acu0
		[18]));
	notech_mux2 i_45314(.S(n_56688), .A(n_44215), .B(to_acu0[18]), .Z(n_41219
		));
	notech_reg to_acu0_reg_19(.CP(n_63173), .D(n_41225), .CD(n_62575), .Q(to_acu0
		[19]));
	notech_mux2 i_45322(.S(n_56688), .A(n_42727), .B(to_acu0[19]), .Z(n_41225
		));
	notech_reg to_acu0_reg_20(.CP(n_63173), .D(n_41231), .CD(n_62575), .Q(to_acu0
		[20]));
	notech_mux2 i_45330(.S(n_56688), .A(n_44216), .B(to_acu0[20]), .Z(n_41231
		));
	notech_reg to_acu0_reg_21(.CP(n_63173), .D(n_41237), .CD(n_62575), .Q(to_acu0
		[21]));
	notech_mux2 i_45338(.S(n_56688), .A(n_42730), .B(to_acu0[21]), .Z(n_41237
		));
	notech_reg to_acu0_reg_22(.CP(n_63173), .D(n_41243), .CD(n_62575), .Q(to_acu0
		[22]));
	notech_mux2 i_45346(.S(n_56688), .A(n_42732), .B(to_acu0[22]), .Z(n_41243
		));
	notech_reg to_acu0_reg_23(.CP(n_63173), .D(n_41249), .CD(n_62575), .Q(to_acu0
		[23]));
	notech_mux2 i_45354(.S(n_56688), .A(n_42735), .B(to_acu0[23]), .Z(n_41249
		));
	notech_reg to_acu0_reg_24(.CP(n_63173), .D(n_41255), .CD(n_62575), .Q(to_acu0
		[24]));
	notech_mux2 i_45362(.S(n_56688), .A(n_42737), .B(to_acu0[24]), .Z(n_41255
		));
	notech_reg to_acu0_reg_25(.CP(n_63173), .D(n_41261), .CD(n_62575), .Q(to_acu0
		[25]));
	notech_mux2 i_45370(.S(n_56688), .A(n_42739), .B(to_acu0[25]), .Z(n_41261
		));
	notech_reg to_acu0_reg_26(.CP(n_63178), .D(n_41267), .CD(n_62575), .Q(to_acu0
		[26]));
	notech_mux2 i_45378(.S(n_56683), .A(n_42742), .B(to_acu0[26]), .Z(n_41267
		));
	notech_reg to_acu0_reg_27(.CP(n_63178), .D(n_41273), .CD(n_62575), .Q(to_acu0
		[27]));
	notech_mux2 i_45386(.S(n_56688), .A(n_42744), .B(to_acu0[27]), .Z(n_41273
		));
	notech_reg to_acu0_reg_28(.CP(n_63178), .D(n_41279), .CD(n_62580), .Q(to_acu0
		[28]));
	notech_mux2 i_45394(.S(n_56683), .A(n_42746), .B(to_acu0[28]), .Z(n_41279
		));
	notech_reg to_acu0_reg_29(.CP(n_63176), .D(n_41285), .CD(n_62580), .Q(to_acu0
		[29]));
	notech_mux2 i_45402(.S(n_56683), .A(n_44217), .B(to_acu0[29]), .Z(n_41285
		));
	notech_reg to_acu0_reg_30(.CP(n_63176), .D(n_41291), .CD(n_62580), .Q(to_acu0
		[30]));
	notech_mux2 i_45410(.S(n_56688), .A(n_44218), .B(to_acu0[30]), .Z(n_41291
		));
	notech_reg to_acu0_reg_31(.CP(n_63178), .D(n_41297), .CD(n_62578), .Q(to_acu0
		[31]));
	notech_mux2 i_45418(.S(n_56688), .A(n_44219), .B(to_acu0[31]), .Z(n_41297
		));
	notech_reg to_acu0_reg_32(.CP(n_63178), .D(n_41303), .CD(n_62578), .Q(to_acu0
		[32]));
	notech_mux2 i_45426(.S(n_56688), .A(n_44221), .B(to_acu0[32]), .Z(n_41303
		));
	notech_reg to_acu0_reg_33(.CP(n_63178), .D(n_41309), .CD(n_62580), .Q(to_acu0
		[33]));
	notech_mux2 i_45434(.S(n_56688), .A(n_42748), .B(to_acu0[33]), .Z(n_41309
		));
	notech_reg to_acu0_reg_34(.CP(n_63178), .D(n_41315), .CD(n_62580), .Q(to_acu0
		[34]));
	notech_mux2 i_45442(.S(n_56688), .A(n_42750), .B(to_acu0[34]), .Z(n_41315
		));
	notech_reg to_acu0_reg_35(.CP(n_63178), .D(n_41321), .CD(n_62580), .Q(to_acu0
		[35]));
	notech_mux2 i_45450(.S(n_3302), .A(n_44222), .B(to_acu0[35]), .Z(n_41321
		));
	notech_reg to_acu0_reg_36(.CP(n_63176), .D(n_41327), .CD(n_62580), .Q(to_acu0
		[36]));
	notech_mux2 i_45458(.S(n_3302), .A(n_44223), .B(to_acu0[36]), .Z(n_41327
		));
	notech_reg to_acu0_reg_37(.CP(n_63176), .D(n_41333), .CD(n_62580), .Q(to_acu0
		[37]));
	notech_mux2 i_45466(.S(n_3302), .A(n_44224), .B(to_acu0[37]), .Z(n_41333
		));
	notech_reg to_acu0_reg_38(.CP(n_63176), .D(n_41339), .CD(n_62578), .Q(to_acu0
		[38]));
	notech_mux2 i_45474(.S(n_3302), .A(n_44225), .B(to_acu0[38]), .Z(n_41339
		));
	notech_nand3 i_21980430(.A(n_2995), .B(inst_deco1[87]), .C(n_59405), .Z(n_1710
		));
	notech_reg to_acu0_reg_39(.CP(n_63176), .D(n_41345), .CD(n_62578), .Q(to_acu0
		[39]));
	notech_mux2 i_45482(.S(n_3302), .A(n_1099100407), .B(to_acu0[39]), .Z(n_41345
		));
	notech_reg to_acu0_reg_40(.CP(n_63176), .D(n_41351), .CD(n_62578), .Q(to_acu0
		[40]));
	notech_mux2 i_45490(.S(n_3302), .A(n_42752), .B(to_acu0[40]), .Z(n_41351
		));
	notech_reg to_acu0_reg_41(.CP(n_63176), .D(n_41357), .CD(n_62578), .Q(to_acu0
		[41]));
	notech_mux2 i_45498(.S(n_3302), .A(n_42754), .B(to_acu0[41]), .Z(n_41357
		));
	notech_nand3 i_21680433(.A(n_2995), .B(inst_deco1[86]), .C(n_59405), .Z(n_1707
		));
	notech_reg to_acu0_reg_42(.CP(n_63176), .D(n_41363), .CD(n_62578), .Q(to_acu0
		[42]));
	notech_mux2 i_45506(.S(n_3302), .A(n_44227), .B(to_acu0[42]), .Z(n_41363
		));
	notech_reg to_acu0_reg_43(.CP(n_63176), .D(n_41369), .CD(n_62578), .Q(to_acu0
		[43]));
	notech_mux2 i_45514(.S(n_3302), .A(n_44228), .B(to_acu0[43]), .Z(n_41369
		));
	notech_reg to_acu0_reg_44(.CP(n_63176), .D(n_41375), .CD(n_62578), .Q(to_acu0
		[44]));
	notech_mux2 i_45522(.S(n_3302), .A(n_44229), .B(to_acu0[44]), .Z(n_41375
		));
	notech_nand3 i_21380436(.A(n_2995), .B(inst_deco1[85]), .C(n_59405), .Z(n_1704
		));
	notech_reg to_acu0_reg_45(.CP(n_63176), .D(n_41381), .CD(n_62578), .Q(to_acu0
		[45]));
	notech_mux2 i_45530(.S(n_56688), .A(n_44230), .B(to_acu0[45]), .Z(n_41381
		));
	notech_reg to_acu0_reg_46(.CP(n_63176), .D(n_41387), .CD(n_62578), .Q(to_acu0
		[46]));
	notech_mux2 i_45538(.S(n_3302), .A(n_44231), .B(to_acu0[46]), .Z(n_41387
		));
	notech_reg to_acu0_reg_47(.CP(n_63143), .D(n_41393), .CD(n_62578), .Q(to_acu0
		[47]));
	notech_mux2 i_45546(.S(n_3302), .A(n_44233), .B(to_acu0[47]), .Z(n_41393
		));
	notech_nand3 i_21080439(.A(n_2995), .B(inst_deco1[84]), .C(n_59405), .Z(n_1701
		));
	notech_reg to_acu0_reg_48(.CP(n_63143), .D(n_41399), .CD(n_62578), .Q(to_acu0
		[48]));
	notech_mux2 i_45554(.S(n_3302), .A(n_44234), .B(to_acu0[48]), .Z(n_41399
		));
	notech_reg to_acu0_reg_49(.CP(n_63143), .D(n_41405), .CD(n_62562), .Q(to_acu0
		[49]));
	notech_mux2 i_45562(.S(n_3302), .A(n_42757), .B(to_acu0[49]), .Z(n_41405
		));
	notech_reg to_acu0_reg_50(.CP(n_63140), .D(n_41411), .CD(n_62542), .Q(to_acu0
		[50]));
	notech_mux2 i_45570(.S(n_3302), .A(n_42760), .B(to_acu0[50]), .Z(n_41411
		));
	notech_nand3 i_20780442(.A(n_2995), .B(inst_deco1[83]), .C(n_59405), .Z(n_1698
		));
	notech_reg to_acu0_reg_51(.CP(n_63143), .D(n_41417), .CD(n_62545), .Q(to_acu0
		[51]));
	notech_mux2 i_45578(.S(n_56679), .A(n_42762), .B(to_acu0[51]), .Z(n_41417
		));
	notech_reg to_acu0_reg_52(.CP(n_63143), .D(n_41423), .CD(n_62542), .Q(to_acu0
		[52]));
	notech_mux2 i_45586(.S(n_56679), .A(n_42764), .B(to_acu0[52]), .Z(n_41423
		));
	notech_reg to_acu0_reg_53(.CP(n_63143), .D(n_41429), .CD(n_62542), .Q(to_acu0
		[53]));
	notech_mux2 i_45594(.S(n_56679), .A(n_44235), .B(to_acu0[53]), .Z(n_41429
		));
	notech_nand3 i_20480445(.A(n_2995), .B(inst_deco1[82]), .C(n_59405), .Z(n_1695
		));
	notech_reg to_acu0_reg_54(.CP(n_63143), .D(n_41435), .CD(n_62542), .Q(to_acu0
		[54]));
	notech_mux2 i_45602(.S(n_56679), .A(n_42573), .B(to_acu0[54]), .Z(n_41435
		));
	notech_reg to_acu0_reg_55(.CP(n_63143), .D(n_41441), .CD(n_62545), .Q(to_acu0
		[55]));
	notech_mux2 i_45610(.S(n_56679), .A(n_42766), .B(to_acu0[55]), .Z(n_41441
		));
	notech_reg to_acu0_reg_56(.CP(n_63143), .D(n_41447), .CD(n_62545), .Q(to_acu0
		[56]));
	notech_mux2 i_45618(.S(n_56679), .A(n_42768), .B(to_acu0[56]), .Z(n_41447
		));
	notech_nand3 i_20180448(.A(n_2995), .B(inst_deco1[81]), .C(n_59405), .Z(n_1692
		));
	notech_reg to_acu0_reg_57(.CP(n_63140), .D(n_41453), .CD(n_62545), .Q(to_acu0
		[57]));
	notech_mux2 i_45626(.S(n_56679), .A(n_42770), .B(to_acu0[57]), .Z(n_41453
		));
	notech_reg to_acu0_reg_58(.CP(n_63140), .D(n_41459), .CD(n_62545), .Q(to_acu0
		[58]));
	notech_mux2 i_45634(.S(n_56679), .A(n_44236), .B(to_acu0[58]), .Z(n_41459
		));
	notech_reg to_acu0_reg_59(.CP(n_63140), .D(n_41465), .CD(n_62545), .Q(to_acu0
		[59]));
	notech_mux2 i_45642(.S(n_56674), .A(n_44237), .B(to_acu0[59]), .Z(n_41465
		));
	notech_nand3 i_19880451(.A(n_2995), .B(inst_deco1[80]), .C(n_59405), .Z(n_1689
		));
	notech_reg to_acu0_reg_60(.CP(n_63140), .D(n_41471), .CD(n_62542), .Q(to_acu0
		[60]));
	notech_mux2 i_45650(.S(n_56674), .A(n_42773), .B(to_acu0[60]), .Z(n_41471
		));
	notech_reg to_acu0_reg_61(.CP(n_63140), .D(n_41477), .CD(n_62542), .Q(to_acu0
		[61]));
	notech_mux2 i_45658(.S(n_56674), .A(n_42775), .B(to_acu0[61]), .Z(n_41477
		));
	notech_reg to_acu0_reg_62(.CP(n_63140), .D(n_41483), .CD(n_62542), .Q(to_acu0
		[62]));
	notech_mux2 i_45666(.S(n_56674), .A(n_44239), .B(to_acu0[62]), .Z(n_41483
		));
	notech_reg to_acu0_reg_63(.CP(n_63140), .D(n_41489), .CD(n_62542), .Q(to_acu0
		[63]));
	notech_mux2 i_45674(.S(n_56679), .A(n_42777), .B(to_acu0[63]), .Z(n_41489
		));
	notech_reg to_acu0_reg_64(.CP(n_63140), .D(n_41495), .CD(n_62542), .Q(to_acu0
		[64]));
	notech_mux2 i_45682(.S(n_56679), .A(n_44240), .B(to_acu0[64]), .Z(n_41495
		));
	notech_reg to_acu0_reg_65(.CP(n_63140), .D(n_41501), .CD(n_62542), .Q(to_acu0
		[65]));
	notech_mux2 i_45690(.S(n_56674), .A(n_44241), .B(to_acu0[65]), .Z(n_41501
		));
	notech_reg to_acu0_reg_66(.CP(n_63140), .D(n_41507), .CD(n_62542), .Q(to_acu0
		[66]));
	notech_mux2 i_45698(.S(n_56674), .A(n_42780), .B(to_acu0[66]), .Z(n_41507
		));
	notech_reg to_acu0_reg_67(.CP(n_63140), .D(n_41513), .CD(n_62542), .Q(to_acu0
		[67]));
	notech_mux2 i_45706(.S(n_56679), .A(n_44242), .B(to_acu0[67]), .Z(n_41513
		));
	notech_reg to_acu0_reg_68(.CP(n_63145), .D(n_41519), .CD(n_62542), .Q(to_acu0
		[68]));
	notech_mux2 i_45714(.S(n_56683), .A(n_44243), .B(to_acu0[68]), .Z(n_41519
		));
	notech_reg to_acu0_reg_69(.CP(n_63145), .D(n_41525), .CD(n_62542), .Q(to_acu0
		[69]));
	notech_mux2 i_45722(.S(n_56683), .A(n_44245), .B(to_acu0[69]), .Z(n_41525
		));
	notech_reg to_acu0_reg_70(.CP(n_63145), .D(n_41531), .CD(n_62542), .Q(to_acu0
		[70]));
	notech_mux2 i_45730(.S(n_56683), .A(n_44246), .B(to_acu0[70]), .Z(n_41531
		));
	notech_reg to_acu0_reg_71(.CP(n_63145), .D(n_41537), .CD(n_62547), .Q(to_acu0
		[71]));
	notech_mux2 i_45738(.S(n_56683), .A(n_44247), .B(to_acu0[71]), .Z(n_41537
		));
	notech_reg to_acu0_reg_72(.CP(n_63145), .D(n_41545), .CD(n_62547), .Q(to_acu0
		[72]));
	notech_mux2 i_45746(.S(n_56683), .A(n_44248), .B(to_acu0[72]), .Z(n_41545
		));
	notech_reg to_acu0_reg_73(.CP(n_63145), .D(n_41551), .CD(n_62547), .Q(to_acu0
		[73]));
	notech_mux2 i_45754(.S(n_56683), .A(n_44249), .B(to_acu0[73]), .Z(n_41551
		));
	notech_reg to_acu0_reg_74(.CP(n_63145), .D(n_41557), .CD(n_62545), .Q(to_acu0
		[74]));
	notech_mux2 i_45762(.S(n_56683), .A(n_44250), .B(to_acu0[74]), .Z(n_41557
		));
	notech_reg to_acu0_reg_75(.CP(n_63145), .D(n_41563), .CD(n_62547), .Q(to_acu0
		[75]));
	notech_mux2 i_45770(.S(n_56683), .A(n_44251), .B(to_acu0[75]), .Z(n_41563
		));
	notech_reg to_acu0_reg_76(.CP(n_63145), .D(n_41569), .CD(n_62547), .Q(to_acu0
		[76]));
	notech_mux2 i_45778(.S(n_56679), .A(n_44252), .B(to_acu0[76]), .Z(n_41569
		));
	notech_reg to_acu0_reg_77(.CP(n_63145), .D(n_41575), .CD(n_62547), .Q(to_acu0
		[77]));
	notech_mux2 i_45786(.S(n_56679), .A(n_44253), .B(to_acu0[77]), .Z(n_41575
		));
	notech_reg to_acu0_reg_78(.CP(n_63145), .D(n_41581), .CD(n_62547), .Q(to_acu0
		[78]));
	notech_mux2 i_45794(.S(n_56679), .A(n_44254), .B(to_acu0[78]), .Z(n_41581
		));
	notech_reg to_acu0_reg_79(.CP(n_63143), .D(n_41588), .CD(n_62547), .Q(to_acu0
		[79]));
	notech_mux2 i_45802(.S(n_56679), .A(n_44255), .B(to_acu0[79]), .Z(n_41588
		));
	notech_reg to_acu0_reg_80(.CP(n_63143), .D(n_41595), .CD(n_62547), .Q(to_acu0
		[80]));
	notech_mux2 i_45810(.S(n_56683), .A(n_44256), .B(to_acu0[80]), .Z(n_41595
		));
	notech_reg to_acu0_reg_81(.CP(n_63143), .D(n_41601), .CD(n_62545), .Q(to_acu0
		[81]));
	notech_mux2 i_45818(.S(n_56683), .A(n_44257), .B(to_acu0[81]), .Z(n_41601
		));
	notech_reg to_acu0_reg_82(.CP(n_63143), .D(n_41608), .CD(n_62545), .Q(to_acu0
		[82]));
	notech_mux2 i_45826(.S(n_56683), .A(n_44258), .B(to_acu0[82]), .Z(n_41608
		));
	notech_reg to_acu0_reg_83(.CP(n_63143), .D(n_41615), .CD(n_62545), .Q(to_acu0
		[83]));
	notech_mux2 i_45834(.S(n_56683), .A(n_44259), .B(to_acu0[83]), .Z(n_41615
		));
	notech_reg to_acu0_reg_84(.CP(n_63143), .D(n_41621), .CD(n_62545), .Q(to_acu0
		[84]));
	notech_mux2 i_45842(.S(n_56627), .A(n_43530), .B(to_acu0[84]), .Z(n_41621
		));
	notech_reg to_acu0_reg_85(.CP(n_63145), .D(n_41627), .CD(n_62545), .Q(to_acu0
		[85]));
	notech_mux2 i_45850(.S(n_56627), .A(n_44260), .B(to_acu0[85]), .Z(n_41627
		));
	notech_reg to_acu0_reg_86(.CP(n_63143), .D(n_41635), .CD(n_62545), .Q(to_acu0
		[86]));
	notech_mux2 i_45858(.S(n_56627), .A(n_44261), .B(to_acu0[86]), .Z(n_41635
		));
	notech_reg to_acu0_reg_87(.CP(n_63143), .D(n_41641), .CD(n_62545), .Q(to_acu0
		[87]));
	notech_mux2 i_45866(.S(n_56627), .A(n_44262), .B(to_acu0[87]), .Z(n_41641
		));
	notech_reg to_acu0_reg_88(.CP(n_63143), .D(n_41647), .CD(n_62545), .Q(to_acu0
		[88]));
	notech_mux2 i_45874(.S(n_56627), .A(n_44263), .B(to_acu0[88]), .Z(n_41647
		));
	notech_reg to_acu0_reg_89(.CP(n_63140), .D(n_41653), .CD(n_62545), .Q(to_acu0
		[89]));
	notech_mux2 i_45882(.S(n_56627), .A(n_44264), .B(to_acu0[89]), .Z(n_41653
		));
	notech_reg to_acu0_reg_90(.CP(n_63135), .D(n_41659), .CD(n_62545), .Q(to_acu0
		[90]));
	notech_mux2 i_45890(.S(n_56627), .A(n_44265), .B(to_acu0[90]), .Z(n_41659
		));
	notech_reg to_acu0_reg_91(.CP(n_63135), .D(n_41665), .CD(n_62545), .Q(to_acu0
		[91]));
	notech_mux2 i_45898(.S(n_56627), .A(n_44266), .B(to_acu0[91]), .Z(n_41665
		));
	notech_reg to_acu0_reg_92(.CP(n_63135), .D(n_41672), .CD(n_62537), .Q(to_acu0
		[92]));
	notech_mux2 i_45906(.S(n_56623), .A(n_42782), .B(to_acu0[92]), .Z(n_41672
		));
	notech_reg to_acu0_reg_93(.CP(n_63135), .D(n_41680), .CD(n_62537), .Q(to_acu0
		[93]));
	notech_mux2 i_45914(.S(n_56623), .A(n_42785), .B(to_acu0[93]), .Z(n_41680
		));
	notech_reg to_acu0_reg_94(.CP(n_63135), .D(n_41686), .CD(n_62537), .Q(to_acu0
		[94]));
	notech_mux2 i_45922(.S(n_56623), .A(n_42789), .B(to_acu0[94]), .Z(n_41686
		));
	notech_reg to_acu0_reg_95(.CP(n_63138), .D(n_41692), .CD(n_62537), .Q(to_acu0
		[95]));
	notech_mux2 i_45930(.S(n_56623), .A(n_42792), .B(to_acu0[95]), .Z(n_41692
		));
	notech_reg to_acu0_reg_96(.CP(n_63138), .D(n_41698), .CD(n_62537), .Q(to_acu0
		[96]));
	notech_mux2 i_45938(.S(n_56623), .A(n_42794), .B(to_acu0[96]), .Z(n_41698
		));
	notech_reg to_acu0_reg_97(.CP(n_63135), .D(n_41705), .CD(n_62537), .Q(to_acu0
		[97]));
	notech_mux2 i_45946(.S(n_56623), .A(n_44267), .B(to_acu0[97]), .Z(n_41705
		));
	notech_reg to_acu0_reg_98(.CP(n_63135), .D(n_41712), .CD(n_62537), .Q(to_acu0
		[98]));
	notech_mux2 i_45954(.S(n_56623), .A(n_44268), .B(to_acu0[98]), .Z(n_41712
		));
	notech_reg to_acu0_reg_99(.CP(n_63135), .D(n_41719), .CD(n_62537), .Q(to_acu0
		[99]));
	notech_mux2 i_45962(.S(n_56623), .A(n_44269), .B(to_acu0[99]), .Z(n_41719
		));
	notech_reg to_acu0_reg_100(.CP(n_63135), .D(n_41725), .CD(n_62537), .Q(to_acu0
		[100]));
	notech_mux2 i_45970(.S(n_56627), .A(n_42797), .B(to_acu0[100]), .Z(n_41725
		));
	notech_reg to_acu0_reg_101(.CP(n_63135), .D(n_41732), .CD(n_62537), .Q(to_acu0
		[101]));
	notech_mux2 i_45978(.S(n_56632), .A(n_42799), .B(to_acu0[101]), .Z(n_41732
		));
	notech_reg to_acu0_reg_102(.CP(n_63135), .D(n_41739), .CD(n_62537), .Q(to_acu0
		[102]));
	notech_mux2 i_45986(.S(n_56632), .A(n_42801), .B(to_acu0[102]), .Z(n_41739
		));
	notech_reg to_acu0_reg_103(.CP(n_63135), .D(n_41746), .CD(n_62537), .Q(to_acu0
		[103]));
	notech_mux2 i_45994(.S(n_56632), .A(n_42804), .B(to_acu0[103]), .Z(n_41746
		));
	notech_reg to_acu0_reg_104(.CP(n_63133), .D(n_41753), .CD(n_62537), .Q(to_acu0
		[104]));
	notech_mux2 i_46002(.S(n_56632), .A(n_42806), .B(to_acu0[104]), .Z(n_41753
		));
	notech_reg to_acu0_reg_105(.CP(n_63135), .D(n_41760), .CD(n_62535), .Q(to_acu0
		[105]));
	notech_mux2 i_46010(.S(n_56632), .A(n_42809), .B(to_acu0[105]), .Z(n_41760
		));
	notech_reg to_acu0_reg_106(.CP(n_63135), .D(n_41766), .CD(n_62535), .Q(to_acu0
		[106]));
	notech_mux2 i_46018(.S(n_56632), .A(n_44270), .B(to_acu0[106]), .Z(n_41766
		));
	notech_reg to_acu0_reg_107(.CP(n_63135), .D(n_41772), .CD(n_62535), .Q(to_acu0
		[107]));
	notech_mux2 i_46026(.S(n_56632), .A(n_42811), .B(to_acu0[107]), .Z(n_41772
		));
	notech_reg to_acu0_reg_108(.CP(n_63135), .D(n_41778), .CD(n_62537), .Q(to_acu0
		[108]));
	notech_mux2 i_46034(.S(n_56632), .A(n_44271), .B(to_acu0[108]), .Z(n_41778
		));
	notech_reg to_acu0_reg_109(.CP(n_63135), .D(n_41784), .CD(n_62537), .Q(to_acu0
		[109]));
	notech_mux2 i_46042(.S(n_56627), .A(n_42813), .B(to_acu0[109]), .Z(n_41784
		));
	notech_reg to_acu0_reg_110(.CP(n_63135), .D(n_41790), .CD(n_62537), .Q(to_acu0
		[110]));
	notech_mux2 i_46050(.S(n_56627), .A(n_44272), .B(to_acu0[110]), .Z(n_41790
		));
	notech_reg to_acu0_reg_111(.CP(n_63138), .D(n_41796), .CD(n_62537), .Q(to_acu0
		[111]));
	notech_mux2 i_46058(.S(n_56627), .A(n_42816), .B(to_acu0[111]), .Z(n_41796
		));
	notech_reg to_acu0_reg_112(.CP(n_63138), .D(n_41803), .CD(n_62537), .Q(to_acu0
		[112]));
	notech_mux2 i_46066(.S(n_56627), .A(n_42818), .B(to_acu0[112]), .Z(n_41803
		));
	notech_reg to_acu0_reg_113(.CP(n_63138), .D(n_41810), .CD(n_62540), .Q(to_acu0
		[113]));
	notech_mux2 i_46074(.S(n_56632), .A(n_42821), .B(to_acu0[113]), .Z(n_41810
		));
	notech_reg to_acu0_reg_114(.CP(n_63138), .D(n_41817), .CD(n_62540), .Q(to_acu0
		[114]));
	notech_mux2 i_46082(.S(n_56632), .A(n_42823), .B(to_acu0[114]), .Z(n_41817
		));
	notech_reg to_acu0_reg_115(.CP(n_63138), .D(n_41823), .CD(n_62540), .Q(to_acu0
		[115]));
	notech_mux2 i_46090(.S(n_56627), .A(n_42825), .B(to_acu0[115]), .Z(n_41823
		));
	notech_reg to_acu0_reg_116(.CP(n_63140), .D(n_41829), .CD(n_62540), .Q(to_acu0
		[116]));
	notech_mux2 i_46098(.S(n_56627), .A(n_42828), .B(to_acu0[116]), .Z(n_41829
		));
	notech_reg to_acu0_reg_117(.CP(n_63140), .D(n_41835), .CD(n_62540), .Q(to_acu0
		[117]));
	notech_mux2 i_46106(.S(n_56614), .A(n_42830), .B(to_acu0[117]), .Z(n_41835
		));
	notech_reg to_acu0_reg_118(.CP(n_63140), .D(n_41841), .CD(n_62542), .Q(to_acu0
		[118]));
	notech_mux2 i_46114(.S(n_56614), .A(n_42833), .B(to_acu0[118]), .Z(n_41841
		));
	notech_reg to_acu0_reg_119(.CP(n_63140), .D(n_41848), .CD(n_62542), .Q(to_acu0
		[119]));
	notech_mux2 i_46122(.S(n_56614), .A(n_42835), .B(to_acu0[119]), .Z(n_41848
		));
	notech_reg to_acu0_reg_120(.CP(n_63140), .D(n_41854), .CD(n_62542), .Q(to_acu0
		[120]));
	notech_mux2 i_46130(.S(n_56614), .A(n_42837), .B(to_acu0[120]), .Z(n_41854
		));
	notech_reg to_acu0_reg_121(.CP(n_63138), .D(n_41860), .CD(n_62540), .Q(to_acu0
		[121]));
	notech_mux2 i_46138(.S(n_56618), .A(n_42840), .B(to_acu0[121]), .Z(n_41860
		));
	notech_reg to_acu0_reg_122(.CP(n_63138), .D(n_41866), .CD(n_62540), .Q(to_acu0
		[122]));
	notech_mux2 i_46146(.S(n_56618), .A(n_42842), .B(to_acu0[122]), .Z(n_41866
		));
	notech_reg to_acu0_reg_123(.CP(n_63138), .D(n_41872), .CD(n_62540), .Q(to_acu0
		[123]));
	notech_mux2 i_46154(.S(n_56618), .A(n_42846), .B(to_acu0[123]), .Z(n_41872
		));
	notech_reg to_acu0_reg_124(.CP(n_63138), .D(n_41878), .CD(n_62540), .Q(to_acu0
		[124]));
	notech_mux2 i_46162(.S(n_56618), .A(n_44273), .B(to_acu0[124]), .Z(n_41878
		));
	notech_reg to_acu0_reg_125(.CP(n_63138), .D(n_41885), .CD(n_62540), .Q(to_acu0
		[125]));
	notech_mux2 i_46170(.S(n_56614), .A(n_44274), .B(to_acu0[125]), .Z(n_41885
		));
	notech_reg to_acu0_reg_126(.CP(n_63138), .D(n_41893), .CD(n_62540), .Q(to_acu0
		[126]));
	notech_mux2 i_46178(.S(n_56614), .A(n_44275), .B(to_acu0[126]), .Z(n_41893
		));
	notech_reg to_acu0_reg_127(.CP(n_63138), .D(n_41900), .CD(n_62540), .Q(to_acu0
		[127]));
	notech_mux2 i_46186(.S(n_56614), .A(n_44276), .B(to_acu0[127]), .Z(n_41900
		));
	notech_reg to_acu0_reg_128(.CP(n_63138), .D(n_41907), .CD(n_62540), .Q(to_acu0
		[128]));
	notech_mux2 i_46194(.S(n_56614), .A(n_44277), .B(to_acu0[128]), .Z(n_41907
		));
	notech_reg to_acu0_reg_129(.CP(n_63138), .D(n_41914), .CD(n_62540), .Q(to_acu0
		[129]));
	notech_mux2 i_46202(.S(n_56614), .A(n_44279), .B(to_acu0[129]), .Z(n_41914
		));
	notech_reg to_acu0_reg_130(.CP(n_63138), .D(n_41921), .CD(n_62540), .Q(to_acu0
		[130]));
	notech_mux2 i_46210(.S(n_56614), .A(n_44280), .B(to_acu0[130]), .Z(n_41921
		));
	notech_reg to_acu0_reg_131(.CP(n_63138), .D(n_41929), .CD(n_62540), .Q(to_acu0
		[131]));
	notech_mux2 i_46218(.S(n_56614), .A(n_44281), .B(to_acu0[131]), .Z(n_41929
		));
	notech_reg to_acu0_reg_132(.CP(n_63155), .D(n_41936), .CD(n_62540), .Q(to_acu0
		[132]));
	notech_mux2 i_46226(.S(n_56614), .A(n_44282), .B(to_acu0[132]), .Z(n_41936
		));
	notech_reg to_acu0_reg_133(.CP(n_63155), .D(n_41943), .CD(n_62540), .Q(to_acu0
		[133]));
	notech_mux2 i_46234(.S(n_56618), .A(n_44283), .B(to_acu0[133]), .Z(n_41943
		));
	notech_reg to_acu0_reg_134(.CP(n_63155), .D(n_41950), .CD(n_62547), .Q(to_acu0
		[134]));
	notech_mux2 i_46242(.S(n_56623), .A(n_42849), .B(to_acu0[134]), .Z(n_41950
		));
	notech_reg to_acu0_reg_135(.CP(n_63155), .D(n_41957), .CD(n_62557), .Q(to_acu0
		[135]));
	notech_mux2 i_46250(.S(n_56623), .A(n_44285), .B(to_acu0[135]), .Z(n_41957
		));
	notech_reg to_acu0_reg_136(.CP(n_63155), .D(n_41965), .CD(n_62557), .Q(to_acu0
		[136]));
	notech_mux2 i_46258(.S(n_56618), .A(n_44286), .B(to_acu0[136]), .Z(n_41965
		));
	notech_reg to_acu0_reg_137(.CP(n_63157), .D(n_41972), .CD(n_62557), .Q(to_acu0
		[137]));
	notech_mux2 i_46266(.S(n_56623), .A(n_44287), .B(to_acu0[137]), .Z(n_41972
		));
	notech_reg to_acu0_reg_138(.CP(n_63157), .D(n_41979), .CD(n_62557), .Q(to_acu0
		[138]));
	notech_mux2 i_46274(.S(n_56623), .A(n_44288), .B(to_acu0[138]), .Z(n_41979
		));
	notech_and4 i_126279399(.A(n_1676), .B(n_44165), .C(n_2379), .D(n_3012),
		 .Z(n_1608));
	notech_reg to_acu0_reg_139(.CP(n_63157), .D(n_41986), .CD(n_62557), .Q(to_acu0
		[139]));
	notech_mux2 i_46282(.S(n_56623), .A(n_44289), .B(to_acu0[139]), .Z(n_41986
		));
	notech_and2 i_125979402(.A(n_62559), .B(n_42554), .Z(n_1607));
	notech_reg to_acu0_reg_140(.CP(n_63155), .D(n_41993), .CD(n_62559), .Q(to_acu0
		[140]));
	notech_mux2 i_46290(.S(n_56623), .A(n_44290), .B(to_acu0[140]), .Z(n_41993
		));
	notech_and4 i_125879403(.A(n_1676), .B(n_2379), .C(n_62557), .D(n_3009),
		 .Z(n_1606));
	notech_reg to_acu0_reg_141(.CP(n_63157), .D(n_42001), .CD(n_62557), .Q(to_acu0
		[141]));
	notech_mux2 i_46298(.S(n_56623), .A(n_44291), .B(to_acu0[141]), .Z(n_42001
		));
	notech_and4 i_125779404(.A(n_2379), .B(n_2859), .C(n_44729), .D(n_3014),
		 .Z(n_1605));
	notech_reg to_acu0_reg_142(.CP(n_63155), .D(n_42008), .CD(n_62557), .Q(to_acu0
		[142]));
	notech_mux2 i_46306(.S(n_56618), .A(n_44293), .B(to_acu0[142]), .Z(n_42008
		));
	notech_nand2 i_125479407(.A(n_2379), .B(n_2383), .Z(n_1604));
	notech_reg to_acu0_reg_143(.CP(n_63155), .D(n_42015), .CD(n_62557), .Q(to_acu0
		[143]));
	notech_mux2 i_46314(.S(n_56618), .A(n_44294), .B(to_acu0[143]), .Z(n_42015
		));
	notech_reg to_acu0_reg_144(.CP(n_63155), .D(n_42022), .CD(n_62557), .Q(to_acu0
		[144]));
	notech_mux2 i_46322(.S(n_56618), .A(n_44295), .B(to_acu0[144]), .Z(n_42022
		));
	notech_reg to_acu0_reg_145(.CP(n_63155), .D(n_42029), .CD(n_62557), .Q(to_acu0
		[145]));
	notech_mux2 i_46330(.S(n_56618), .A(n_44296), .B(to_acu0[145]), .Z(n_42029
		));
	notech_or4 i_124879413(.A(in128[1]), .B(n_17054783), .C(n_44728), .D(n_44659
		), .Z(n_1601));
	notech_reg to_acu0_reg_146(.CP(n_63155), .D(n_42037), .CD(n_62557), .Q(to_acu0
		[146]));
	notech_mux2 i_46338(.S(n_56618), .A(n_44297), .B(to_acu0[146]), .Z(n_42037
		));
	notech_nao3 i_39280268(.A(n_43434), .B(n_43431), .C(n_5767), .Z(n_1600)
		);
	notech_reg to_acu0_reg_147(.CP(n_63155), .D(n_42044), .CD(n_62554), .Q(to_acu0
		[147]));
	notech_mux2 i_46346(.S(n_56618), .A(n_44299), .B(to_acu0[147]), .Z(n_42044
		));
	notech_or4 i_39080270(.A(i_ptr[1]), .B(i_ptr[0]), .C(i_ptr[3]), .D(i_ptr
		[2]), .Z(n_1599));
	notech_reg to_acu0_reg_148(.CP(n_63155), .D(n_42051), .CD(n_62554), .Q(to_acu0
		[148]));
	notech_mux2 i_46354(.S(n_56618), .A(n_44300), .B(to_acu0[148]), .Z(n_42051
		));
	notech_reg to_acu0_reg_149(.CP(n_63155), .D(n_42058), .CD(n_62557), .Q(to_acu0
		[149]));
	notech_mux2 i_46362(.S(n_56618), .A(n_44301), .B(to_acu0[149]), .Z(n_42058
		));
	notech_reg to_acu0_reg_150(.CP(n_63155), .D(n_42065), .CD(n_62557), .Q(to_acu0
		[150]));
	notech_mux2 i_46370(.S(n_56632), .A(n_44302), .B(to_acu0[150]), .Z(n_42065
		));
	notech_reg to_acu0_reg_151(.CP(n_63155), .D(n_42073), .CD(n_62557), .Q(to_acu0
		[151]));
	notech_mux2 i_46378(.S(n_56646), .A(n_44303), .B(to_acu0[151]), .Z(n_42073
		));
	notech_reg to_acu0_reg_152(.CP(n_63155), .D(n_42080), .CD(n_62557), .Q(to_acu0
		[152]));
	notech_mux2 i_46386(.S(n_56646), .A(n_44305), .B(to_acu0[152]), .Z(n_42080
		));
	notech_reg to_acu0_reg_153(.CP(n_63160), .D(n_42087), .CD(n_62557), .Q(to_acu0
		[153]));
	notech_mux2 i_46394(.S(n_56646), .A(n_44306), .B(to_acu0[153]), .Z(n_42087
		));
	notech_reg to_acu0_reg_154(.CP(n_63160), .D(n_42094), .CD(n_62559), .Q(to_acu0
		[154]));
	notech_mux2 i_46402(.S(n_56646), .A(n_44307), .B(to_acu0[154]), .Z(n_42094
		));
	notech_reg to_acu0_reg_155(.CP(n_63157), .D(n_42101), .CD(n_62562), .Q(to_acu0
		[155]));
	notech_mux2 i_46410(.S(n_56646), .A(n_44308), .B(to_acu0[155]), .Z(n_42101
		));
	notech_reg to_acu0_reg_156(.CP(n_63157), .D(n_42109), .CD(n_62559), .Q(to_acu0
		[156]));
	notech_mux2 i_46418(.S(n_56646), .A(n_44309), .B(to_acu0[156]), .Z(n_42109
		));
	notech_reg to_acu0_reg_157(.CP(n_63157), .D(n_42116), .CD(n_62559), .Q(to_acu0
		[157]));
	notech_mux2 i_46426(.S(n_56646), .A(n_44311), .B(to_acu0[157]), .Z(n_42116
		));
	notech_reg to_acu0_reg_158(.CP(n_63160), .D(n_42123), .CD(n_62559), .Q(to_acu0
		[158]));
	notech_mux2 i_46434(.S(n_56646), .A(n_44312), .B(to_acu0[158]), .Z(n_42123
		));
	notech_reg to_acu0_reg_159(.CP(n_63160), .D(n_42130), .CD(n_62562), .Q(to_acu0
		[159]));
	notech_mux2 i_46442(.S(n_56646), .A(n_44313), .B(to_acu0[159]), .Z(n_42130
		));
	notech_reg to_acu0_reg_160(.CP(n_63160), .D(n_42137), .CD(n_62562), .Q(to_acu0
		[160]));
	notech_mux2 i_46450(.S(n_56646), .A(n_44314), .B(to_acu0[160]), .Z(n_42137
		));
	notech_reg to_acu0_reg_161(.CP(n_63160), .D(n_42145), .CD(n_62562), .Q(to_acu0
		[161]));
	notech_mux2 i_46458(.S(n_56642), .A(n_44315), .B(to_acu0[161]), .Z(n_42145
		));
	notech_reg to_acu0_reg_162(.CP(n_63160), .D(n_42152), .CD(n_62562), .Q(to_acu0
		[162]));
	notech_mux2 i_46466(.S(n_56646), .A(n_44317), .B(to_acu0[162]), .Z(n_42152
		));
	notech_reg to_acu0_reg_163(.CP(n_63157), .D(n_42159), .CD(n_62562), .Q(to_acu0
		[163]));
	notech_mux2 i_46474(.S(n_56646), .A(n_44318), .B(to_acu0[163]), .Z(n_42159
		));
	notech_reg to_acu0_reg_164(.CP(n_63157), .D(n_42166), .CD(n_62559), .Q(to_acu0
		[164]));
	notech_mux2 i_46482(.S(n_56646), .A(n_44319), .B(to_acu0[164]), .Z(n_42166
		));
	notech_reg to_acu0_reg_165(.CP(n_63157), .D(n_42173), .CD(n_62559), .Q(to_acu0
		[165]));
	notech_mux2 i_46490(.S(n_56646), .A(n_44320), .B(to_acu0[165]), .Z(n_42173
		));
	notech_reg to_acu0_reg_166(.CP(n_63157), .D(n_42181), .CD(n_62559), .Q(to_acu0
		[166]));
	notech_mux2 i_46498(.S(n_56646), .A(n_44321), .B(to_acu0[166]), .Z(n_42181
		));
	notech_reg to_acu0_reg_167(.CP(n_63157), .D(n_42188), .CD(n_62559), .Q(to_acu0
		[167]));
	notech_mux2 i_46506(.S(n_56651), .A(n_44323), .B(to_acu0[167]), .Z(n_42188
		));
	notech_reg to_acu0_reg_168(.CP(n_63157), .D(n_42195), .CD(n_62559), .Q(to_acu0
		[168]));
	notech_mux2 i_46514(.S(n_56651), .A(n_44324), .B(to_acu0[168]), .Z(n_42195
		));
	notech_reg to_acu0_reg_169(.CP(n_63157), .D(n_42202), .CD(n_62559), .Q(to_acu0
		[169]));
	notech_mux2 i_46522(.S(n_56651), .A(n_44325), .B(to_acu0[169]), .Z(n_42202
		));
	notech_reg to_acu0_reg_170(.CP(n_63157), .D(n_42209), .CD(n_62559), .Q(to_acu0
		[170]));
	notech_mux2 i_46530(.S(n_56651), .A(n_44326), .B(to_acu0[170]), .Z(n_42209
		));
	notech_reg to_acu0_reg_171(.CP(n_63157), .D(n_42217), .CD(n_62559), .Q(to_acu0
		[171]));
	notech_mux2 i_46538(.S(n_56651), .A(n_44327), .B(to_acu0[171]), .Z(n_42217
		));
	notech_reg to_acu0_reg_172(.CP(n_63157), .D(n_42224), .CD(n_62559), .Q(to_acu0
		[172]));
	notech_mux2 i_46546(.S(n_56655), .A(n_44329), .B(to_acu0[172]), .Z(n_42224
		));
	notech_reg to_acu0_reg_173(.CP(n_63157), .D(n_42231), .CD(n_62559), .Q(to_acu0
		[173]));
	notech_mux2 i_46554(.S(n_56655), .A(n_44330), .B(to_acu0[173]), .Z(n_42231
		));
	notech_reg to_acu0_reg_174(.CP(n_63155), .D(n_42238), .CD(n_62559), .Q(to_acu0
		[174]));
	notech_mux2 i_46562(.S(n_56651), .A(n_44331), .B(to_acu0[174]), .Z(n_42238
		));
	notech_reg to_acu0_reg_175(.CP(n_63150), .D(n_42245), .CD(n_62552), .Q(to_acu0
		[175]));
	notech_mux2 i_46570(.S(n_56651), .A(n_44332), .B(to_acu0[175]), .Z(n_42245
		));
	notech_reg to_acu0_reg_176(.CP(n_63150), .D(n_42253), .CD(n_62552), .Q(to_acu0
		[176]));
	notech_mux2 i_46578(.S(n_56651), .A(n_44333), .B(to_acu0[176]), .Z(n_42253
		));
	notech_reg to_acu0_reg_177(.CP(n_63150), .D(n_42260), .CD(n_62552), .Q(to_acu0
		[177]));
	notech_mux2 i_46586(.S(n_56651), .A(n_44335), .B(to_acu0[177]), .Z(n_42260
		));
	notech_reg to_acu0_reg_178(.CP(n_63150), .D(n_42267), .CD(n_62552), .Q(to_acu0
		[178]));
	notech_mux2 i_46594(.S(n_56651), .A(n_44336), .B(to_acu0[178]), .Z(n_42267
		));
	notech_reg to_acu0_reg_179(.CP(n_63150), .D(n_42274), .CD(n_62552), .Q(to_acu0
		[179]));
	notech_mux2 i_46602(.S(n_56651), .A(n_44337), .B(to_acu0[179]), .Z(n_42274
		));
	notech_reg to_acu0_reg_180(.CP(n_63150), .D(n_42281), .CD(n_62552), .Q(to_acu0
		[180]));
	notech_mux2 i_46610(.S(n_56651), .A(n_44338), .B(to_acu0[180]), .Z(n_42281
		));
	notech_reg to_acu0_reg_181(.CP(n_63150), .D(n_42289), .CD(n_62552), .Q(to_acu0
		[181]));
	notech_mux2 i_46618(.S(n_56651), .A(n_44339), .B(to_acu0[181]), .Z(n_42289
		));
	notech_reg to_acu0_reg_182(.CP(n_63150), .D(n_42296), .CD(n_62552), .Q(to_acu0
		[182]));
	notech_mux2 i_46626(.S(n_56651), .A(n_44340), .B(to_acu0[182]), .Z(n_42296
		));
	notech_reg to_acu0_reg_183(.CP(n_63150), .D(n_42303), .CD(n_62552), .Q(to_acu0
		[183]));
	notech_mux2 i_46634(.S(n_56651), .A(n_44341), .B(to_acu0[183]), .Z(n_42303
		));
	notech_reg to_acu0_reg_184(.CP(n_63150), .D(n_42310), .CD(n_62552), .Q(to_acu0
		[184]));
	notech_mux2 i_46642(.S(n_56612), .A(n_44342), .B(to_acu0[184]), .Z(n_42310
		));
	notech_reg to_acu0_reg_185(.CP(n_63150), .D(n_42317), .CD(n_62552), .Q(to_acu0
		[185]));
	notech_mux2 i_46650(.S(n_56612), .A(n_44343), .B(to_acu0[185]), .Z(n_42317
		));
	notech_reg to_acu0_reg_186(.CP(n_63145), .D(n_42325), .CD(n_62547), .Q(to_acu0
		[186]));
	notech_mux2 i_46658(.S(n_56612), .A(n_44344), .B(to_acu0[186]), .Z(n_42325
		));
	notech_reg to_acu0_reg_187(.CP(n_63145), .D(n_42332), .CD(n_62547), .Q(to_acu0
		[187]));
	notech_mux2 i_46666(.S(n_56612), .A(n_44345), .B(to_acu0[187]), .Z(n_42332
		));
	notech_reg to_acu0_reg_188(.CP(n_63145), .D(n_42339), .CD(n_62547), .Q(to_acu0
		[188]));
	notech_mux2 i_46674(.S(n_56612), .A(n_44346), .B(to_acu0[188]), .Z(n_42339
		));
	notech_reg to_acu0_reg_189(.CP(n_63145), .D(n_42346), .CD(n_62547), .Q(to_acu0
		[189]));
	notech_mux2 i_46682(.S(n_56612), .A(n_44347), .B(to_acu0[189]), .Z(n_42346
		));
	notech_reg to_acu0_reg_190(.CP(n_63145), .D(n_42353), .CD(n_62547), .Q(to_acu0
		[190]));
	notech_mux2 i_46690(.S(n_56612), .A(n_44348), .B(to_acu0[190]), .Z(n_42353
		));
	notech_reg to_acu0_reg_191(.CP(n_63150), .D(n_42361), .CD(n_62552), .Q(to_acu0
		[191]));
	notech_mux2 i_46698(.S(n_56612), .A(n_44349), .B(to_acu0[191]), .Z(n_42361
		));
	notech_reg to_acu0_reg_192(.CP(n_63150), .D(n_42368), .CD(n_62552), .Q(to_acu0
		[192]));
	notech_mux2 i_46706(.S(n_56632), .A(n_44350), .B(to_acu0[192]), .Z(n_42368
		));
	notech_reg to_acu0_reg_193(.CP(n_63150), .D(n_42375), .CD(n_62547), .Q(to_acu0
		[193]));
	notech_mux2 i_46714(.S(n_56632), .A(n_44351), .B(to_acu0[193]), .Z(n_42375
		));
	notech_reg to_acu0_reg_194(.CP(n_63145), .D(n_42382), .CD(n_62547), .Q(to_acu0
		[194]));
	notech_mux2 i_46722(.S(n_56632), .A(n_44352), .B(to_acu0[194]), .Z(n_42382
		));
	notech_reg to_acu0_reg_195(.CP(n_63150), .D(n_42389), .CD(n_62547), .Q(to_acu0
		[195]));
	notech_mux2 i_46730(.S(n_56632), .A(n_44353), .B(to_acu0[195]), .Z(n_42389
		));
	notech_reg to_acu0_reg_196(.CP(n_63152), .D(n_42397), .CD(n_62554), .Q(to_acu0
		[196]));
	notech_mux2 i_46738(.S(n_56612), .A(n_44354), .B(to_acu0[196]), .Z(n_42397
		));
	notech_reg to_acu0_reg_197(.CP(n_63152), .D(n_42404), .CD(n_62554), .Q(to_acu0
		[197]));
	notech_mux2 i_46746(.S(n_56612), .A(n_44355), .B(to_acu0[197]), .Z(n_42404
		));
	notech_reg to_acu0_reg_198(.CP(n_63152), .D(n_42411), .CD(n_62554), .Q(to_acu0
		[198]));
	notech_mux2 i_46754(.S(n_56612), .A(n_44356), .B(to_acu0[198]), .Z(n_42411
		));
	notech_reg to_acu0_reg_199(.CP(n_63152), .D(n_42418), .CD(n_62554), .Q(to_acu0
		[199]));
	notech_mux2 i_46762(.S(n_56612), .A(n_44357), .B(to_acu0[199]), .Z(n_42418
		));
	notech_reg to_acu0_reg_200(.CP(n_63152), .D(n_42425), .CD(n_62554), .Q(to_acu0
		[200]));
	notech_mux2 i_46770(.S(n_56612), .A(n_44358), .B(to_acu0[200]), .Z(n_42425
		));
	notech_reg to_acu0_reg_201(.CP(n_63152), .D(n_42433), .CD(n_62554), .Q(to_acu0
		[201]));
	notech_mux2 i_46778(.S(n_56642), .A(n_44359), .B(to_acu0[201]), .Z(n_42433
		));
	notech_reg to_acu0_reg_202(.CP(n_63152), .D(n_42440), .CD(n_62554), .Q(to_acu0
		[202]));
	notech_mux2 i_46786(.S(n_56642), .A(n_44361), .B(to_acu0[202]), .Z(n_42440
		));
	notech_reg to_acu0_reg_203(.CP(n_63152), .D(n_42447), .CD(n_62554), .Q(to_acu0
		[203]));
	notech_mux2 i_46794(.S(n_56642), .A(n_44362), .B(to_acu0[203]), .Z(n_42447
		));
	notech_reg to_acu0_reg_204(.CP(n_63152), .D(n_42454), .CD(n_62554), .Q(to_acu0
		[204]));
	notech_mux2 i_46802(.S(n_56642), .A(n_44363), .B(to_acu0[204]), .Z(n_42454
		));
	notech_reg to_acu0_reg_205(.CP(n_63152), .D(n_42461), .CD(n_62554), .Q(to_acu0
		[205]));
	notech_mux2 i_46810(.S(n_56642), .A(n_44364), .B(to_acu0[205]), .Z(n_42461
		));
	notech_reg to_acu0_reg_206(.CP(n_63152), .D(n_42469), .CD(n_62554), .Q(to_acu0
		[206]));
	notech_mux2 i_46818(.S(n_56642), .A(n_44365), .B(to_acu0[206]), .Z(n_42469
		));
	notech_reg to_acu0_reg_207(.CP(n_63152), .D(n_42476), .CD(n_62552), .Q(to_acu0
		[207]));
	notech_mux2 i_46826(.S(n_56642), .A(n_44366), .B(to_acu0[207]), .Z(n_42476
		));
	notech_reg to_acu0_reg_208(.CP(n_63152), .D(n_42483), .CD(n_62552), .Q(to_acu0
		[208]));
	notech_mux2 i_46834(.S(n_56642), .A(n_44367), .B(to_acu0[208]), .Z(n_42483
		));
	notech_nor2 i_31180346(.A(n_59157), .B(n_42555), .Z(n_1538));
	notech_reg to_acu0_reg_209(.CP(n_63150), .D(n_42490), .CD(n_62552), .Q(to_acu0
		[209]));
	notech_mux2 i_46842(.S(n_56642), .A(n_44368), .B(to_acu0[209]), .Z(n_42490
		));
	notech_nao3 i_28580372(.A(cpl[0]), .B(cpl[1]), .C(n_1912), .Z(n_1537));
	notech_reg to_acu0_reg_210(.CP(n_63150), .D(n_42497), .CD(n_62552), .Q(to_acu0
		[210]));
	notech_mux2 i_46850(.S(n_56642), .A(n_43533), .B(to_acu0[210]), .Z(n_42497
		));
	notech_reg opz0_reg_0(.CP(n_63150), .D(n_42505), .CD(n_62552), .Q(opz0[0
		]));
	notech_mux2 i_46858(.S(n_56612), .A(n_42562), .B(opz0[0]), .Z(n_42505)
		);
	notech_reg opz0_reg_1(.CP(n_63152), .D(n_42512), .CD(n_62554), .Q(opz0[1
		]));
	notech_mux2 i_46866(.S(n_56612), .A(n_42563), .B(opz0[1]), .Z(n_42512)
		);
	notech_reg_set opz0_reg_2(.CP(n_63152), .D(n_42519), .SD(n_62554), .Q(opz0
		[2]));
	notech_mux2 i_46874(.S(n_56642), .A(n_2931), .B(opz0[2]), .Z(n_42519));
	notech_and2 i_9580633(.A(n_44744), .B(n_60859), .Z(n_1533));
	notech_reg reps0_reg_0(.CP(n_63152), .D(n_42526), .CD(n_62554), .Q(reps0
		[0]));
	notech_mux2 i_46882(.S(n_56642), .A(n_42559), .B(reps0[0]), .Z(n_42526)
		);
	notech_nao3 i_4080636(.A(n_2395), .B(n_44744), .C(n_60248), .Z(n_5767)
		);
	notech_reg reps0_reg_1(.CP(n_63152), .D(n_42533), .CD(n_62554), .Q(reps0
		[1]));
	notech_mux2 i_46890(.S(n_56642), .A(n_42560), .B(reps0[1]), .Z(n_42533)
		);
	notech_reg reps0_reg_2(.CP(n_63152), .D(n_42541), .CD(n_62554), .Q(reps0
		[2]));
	notech_mux2 i_46898(.S(n_56642), .A(n_42561), .B(reps0[2]), .Z(n_42541)
		);
	notech_inv i_52104(.A(n_5712), .Z(n_42548));
	notech_inv i_52105(.A(n_2997), .Z(n_42549));
	notech_inv i_52106(.A(n_1598100903), .Z(n_42550));
	notech_inv i_52107(.A(n_1878), .Z(n_42551));
	notech_inv i_52108(.A(n_2957), .Z(n_42553));
	notech_inv i_52109(.A(n_5765), .Z(n_42554));
	notech_inv i_52110(.A(n_160356214), .Z(n_42555));
	notech_inv i_52111(.A(n_1892), .Z(n_42556));
	notech_inv i_52113(.A(n_2941), .Z(n_42559));
	notech_inv i_52114(.A(n_2939), .Z(n_42560));
	notech_inv i_52115(.A(n_2937), .Z(n_42561));
	notech_inv i_52116(.A(n_2935), .Z(n_42562));
	notech_inv i_52117(.A(n_2933), .Z(n_42563));
	notech_inv i_52118(.A(n_2929), .Z(n_42565));
	notech_inv i_52119(.A(n_2927), .Z(n_42566));
	notech_inv i_52120(.A(n_2925), .Z(n_42567));
	notech_inv i_52121(.A(n_2923), .Z(n_42568));
	notech_inv i_52122(.A(n_2921), .Z(n_42569));
	notech_inv i_52123(.A(n_2919), .Z(n_42571));
	notech_inv i_52124(.A(n_2917), .Z(n_42572));
	notech_inv i_52125(.A(n_2915), .Z(n_42573));
	notech_inv i_52126(.A(n_2904), .Z(n_42574));
	notech_inv i_52127(.A(n_2902), .Z(n_42575));
	notech_inv i_52128(.A(n_2900), .Z(n_42577));
	notech_inv i_52129(.A(n_2898), .Z(n_42578));
	notech_inv i_52130(.A(n_2896), .Z(n_42579));
	notech_inv i_52131(.A(n_2894), .Z(n_42580));
	notech_inv i_52132(.A(n_2890), .Z(n_42581));
	notech_inv i_52133(.A(n_2888), .Z(n_42583));
	notech_inv i_52134(.A(n_2881), .Z(n_42584));
	notech_inv i_52135(.A(n_2871), .Z(n_42585));
	notech_inv i_52136(.A(n_2842), .Z(n_42586));
	notech_inv i_52137(.A(n_2840), .Z(n_42587));
	notech_inv i_52138(.A(n_2838), .Z(n_42589));
	notech_inv i_52139(.A(n_2836), .Z(n_42590));
	notech_inv i_52140(.A(n_2834), .Z(n_42591));
	notech_inv i_52141(.A(n_2832), .Z(n_42592));
	notech_inv i_52142(.A(n_2830), .Z(n_42593));
	notech_inv i_52143(.A(n_2828), .Z(n_42595));
	notech_inv i_52144(.A(n_2826), .Z(n_42596));
	notech_inv i_52145(.A(n_2824), .Z(n_42597));
	notech_inv i_52146(.A(n_2822), .Z(n_42598));
	notech_inv i_52147(.A(n_2820), .Z(n_42599));
	notech_inv i_52148(.A(n_2818), .Z(n_42601));
	notech_inv i_52149(.A(n_1240100547), .Z(n_42602));
	notech_inv i_52150(.A(n_2816), .Z(n_42603));
	notech_inv i_52151(.A(n_1621100926), .Z(n_42604));
	notech_inv i_52152(.A(n_2814), .Z(n_42605));
	notech_inv i_52153(.A(n_2812), .Z(n_42607));
	notech_inv i_52154(.A(n_2810), .Z(n_42608));
	notech_inv i_52155(.A(n_2808), .Z(n_42609));
	notech_inv i_52156(.A(n_2806), .Z(n_42610));
	notech_inv i_52157(.A(n_2401), .Z(n_42611));
	notech_inv i_52158(.A(n_1632100937), .Z(n_42613));
	notech_inv i_52159(.A(n_2804), .Z(n_42614));
	notech_inv i_52160(.A(n_2802), .Z(n_42615));
	notech_inv i_52161(.A(n_1634100939), .Z(n_42616));
	notech_inv i_52162(.A(n_1915), .Z(start));
	notech_inv i_52163(.A(n_2800), .Z(n_42619));
	notech_inv i_52164(.A(n_2798), .Z(n_42620));
	notech_inv i_52165(.A(n_2796), .Z(n_42621));
	notech_inv i_52166(.A(term_f), .Z(n_42622));
	notech_inv i_52167(.A(n_2794), .Z(n_42623));
	notech_inv i_52168(.A(n_2792), .Z(n_42625));
	notech_inv i_52169(.A(n_2790), .Z(n_42626));
	notech_inv i_52170(.A(n_2788), .Z(n_42627));
	notech_inv i_52171(.A(n_2786), .Z(n_42628));
	notech_inv i_52172(.A(n_2784), .Z(n_42629));
	notech_inv i_52173(.A(n_2782), .Z(n_42631));
	notech_inv i_52174(.A(n_2780), .Z(n_42632));
	notech_inv i_52175(.A(n_2778), .Z(n_42633));
	notech_inv i_52176(.A(n_2776), .Z(n_42634));
	notech_inv i_52177(.A(n_2774), .Z(n_42635));
	notech_inv i_52178(.A(n_2772), .Z(n_42637));
	notech_inv i_52179(.A(\fpu_indrm[2] ), .Z(n_42638));
	notech_inv i_52180(.A(n_2770), .Z(n_42639));
	notech_inv i_52181(.A(n_2768), .Z(n_42640));
	notech_inv i_52182(.A(\fpu_indrm[3] ), .Z(n_42641));
	notech_inv i_52183(.A(n_2766), .Z(n_42643));
	notech_inv i_52184(.A(n_2764), .Z(n_42644));
	notech_inv i_52185(.A(\fpu_indrm[4] ), .Z(n_42645));
	notech_inv i_52186(.A(n_2762), .Z(n_42646));
	notech_inv i_52187(.A(n_2760), .Z(n_42647));
	notech_inv i_52188(.A(n_2758), .Z(n_42648));
	notech_inv i_52189(.A(n_2756), .Z(n_42649));
	notech_inv i_52190(.A(n_2754), .Z(n_42650));
	notech_inv i_52191(.A(n_2752), .Z(n_42651));
	notech_inv i_52192(.A(n_2750), .Z(n_42652));
	notech_inv i_52193(.A(n_2748), .Z(n_42653));
	notech_inv i_52194(.A(n_2746), .Z(n_42654));
	notech_inv i_52195(.A(n_2744), .Z(n_42655));
	notech_inv i_52196(.A(n_2742), .Z(n_42656));
	notech_inv i_52197(.A(n_2740), .Z(n_42657));
	notech_inv i_52198(.A(n_2738), .Z(n_42659));
	notech_inv i_52199(.A(n_2736), .Z(n_42660));
	notech_inv i_52200(.A(n_2734), .Z(n_42661));
	notech_inv i_52201(.A(n_2732), .Z(n_42662));
	notech_inv i_52202(.A(n_2730), .Z(n_42663));
	notech_inv i_52203(.A(n_2728), .Z(n_42665));
	notech_inv i_52204(.A(n_2726), .Z(n_42666));
	notech_inv i_52205(.A(n_2724), .Z(n_42667));
	notech_inv i_52206(.A(n_2722), .Z(n_42668));
	notech_inv i_52207(.A(n_2720), .Z(n_42669));
	notech_inv i_52208(.A(\imm2[0] ), .Z(n_42671));
	notech_inv i_52209(.A(n_2718), .Z(n_42672));
	notech_inv i_52210(.A(\imm2[1] ), .Z(n_42673));
	notech_inv i_52211(.A(n_2716), .Z(n_42674));
	notech_inv i_52212(.A(\imm2[2] ), .Z(n_42675));
	notech_inv i_52213(.A(n_2714), .Z(n_42676));
	notech_inv i_52214(.A(\imm2[3] ), .Z(n_42677));
	notech_inv i_52215(.A(n_2712), .Z(n_42678));
	notech_inv i_52216(.A(\imm2[4] ), .Z(n_42679));
	notech_inv i_52217(.A(n_2710), .Z(n_42680));
	notech_inv i_52218(.A(\imm2[5] ), .Z(n_42681));
	notech_inv i_52219(.A(\imm2[6] ), .Z(n_42682));
	notech_inv i_52220(.A(n_2696), .Z(n_42683));
	notech_inv i_52221(.A(\imm2[7] ), .Z(n_42684));
	notech_inv i_52222(.A(\imm2[8] ), .Z(n_42685));
	notech_inv i_52223(.A(\imm2[9] ), .Z(n_42686));
	notech_inv i_52224(.A(\imm2[10] ), .Z(n_42687));
	notech_inv i_52225(.A(\imm2[11] ), .Z(n_42688));
	notech_inv i_52226(.A(\imm2[12] ), .Z(n_42689));
	notech_inv i_52227(.A(\imm2[13] ), .Z(n_42690));
	notech_inv i_52228(.A(\imm2[14] ), .Z(n_42691));
	notech_inv i_52229(.A(\imm2[15] ), .Z(n_42692));
	notech_inv i_52230(.A(\imm2[16] ), .Z(n_42693));
	notech_inv i_52231(.A(\imm2[17] ), .Z(n_42694));
	notech_inv i_52232(.A(\imm2[18] ), .Z(n_42695));
	notech_inv i_52233(.A(\imm2[19] ), .Z(n_42696));
	notech_inv i_52234(.A(\imm2[20] ), .Z(n_42697));
	notech_inv i_52235(.A(\imm2[21] ), .Z(n_42698));
	notech_inv i_52236(.A(\imm2[22] ), .Z(n_42699));
	notech_inv i_52237(.A(\imm2[23] ), .Z(n_42700));
	notech_inv i_52238(.A(\imm2[24] ), .Z(n_42701));
	notech_inv i_52239(.A(\imm2[25] ), .Z(n_42702));
	notech_inv i_52240(.A(\imm2[26] ), .Z(n_42703));
	notech_inv i_52241(.A(\imm2[27] ), .Z(n_42704));
	notech_inv i_52242(.A(\imm2[28] ), .Z(n_42705));
	notech_inv i_52243(.A(\imm2[29] ), .Z(n_42706));
	notech_inv i_52244(.A(\imm2[30] ), .Z(n_42707));
	notech_inv i_52245(.A(\imm2[31] ), .Z(n_42708));
	notech_inv i_52246(.A(\imm2[32] ), .Z(n_42709));
	notech_inv i_52247(.A(\imm2[33] ), .Z(n_42710));
	notech_inv i_52248(.A(\imm2[34] ), .Z(n_42711));
	notech_inv i_52249(.A(\imm2[35] ), .Z(n_42712));
	notech_inv i_52250(.A(\imm2[36] ), .Z(n_42713));
	notech_inv i_52251(.A(\imm2[37] ), .Z(n_42714));
	notech_inv i_52252(.A(\imm2[38] ), .Z(n_42715));
	notech_inv i_52253(.A(\imm2[39] ), .Z(n_42716));
	notech_inv i_52254(.A(\imm2[40] ), .Z(n_42717));
	notech_inv i_52255(.A(\imm2[41] ), .Z(n_42718));
	notech_inv i_52256(.A(\imm2[42] ), .Z(n_42719));
	notech_inv i_52257(.A(\imm2[43] ), .Z(n_42720));
	notech_inv i_52258(.A(n_2850), .Z(n_42721));
	notech_inv i_52259(.A(\imm2[44] ), .Z(n_42722));
	notech_inv i_52260(.A(\imm2[45] ), .Z(n_42723));
	notech_inv i_52261(.A(n_2391), .Z(n_42724));
	notech_inv i_52262(.A(\imm2[46] ), .Z(n_42725));
	notech_inv i_52263(.A(\imm2[47] ), .Z(n_42726));
	notech_inv i_52264(.A(n_3861), .Z(n_42727));
	notech_inv i_52265(.A(\imm1[0] ), .Z(n_42729));
	notech_inv i_52266(.A(n_3860), .Z(n_42730));
	notech_inv i_52267(.A(\imm1[1] ), .Z(n_42731));
	notech_inv i_52268(.A(n_3859), .Z(n_42732));
	notech_inv i_52269(.A(\imm1[2] ), .Z(n_42733));
	notech_inv i_52270(.A(n_3858), .Z(n_42735));
	notech_inv i_52271(.A(\imm1[3] ), .Z(n_42736));
	notech_inv i_52272(.A(n_3857), .Z(n_42737));
	notech_inv i_52273(.A(\imm1[4] ), .Z(n_42738));
	notech_inv i_52274(.A(n_3856), .Z(n_42739));
	notech_inv i_52275(.A(\imm1[5] ), .Z(n_42741));
	notech_inv i_52276(.A(n_3855), .Z(n_42742));
	notech_inv i_52277(.A(\imm1[6] ), .Z(n_42743));
	notech_inv i_52278(.A(n_3854), .Z(n_42744));
	notech_inv i_52279(.A(\imm1[7] ), .Z(n_42745));
	notech_inv i_52280(.A(n_3853), .Z(n_42746));
	notech_inv i_52281(.A(\imm1[8] ), .Z(n_42747));
	notech_inv i_52282(.A(n_3852), .Z(n_42748));
	notech_inv i_52283(.A(\imm1[9] ), .Z(n_42749));
	notech_inv i_52284(.A(n_3851), .Z(n_42750));
	notech_inv i_52285(.A(\imm1[10] ), .Z(n_42751));
	notech_inv i_52286(.A(n_3850), .Z(n_42752));
	notech_inv i_52287(.A(\imm1[11] ), .Z(n_42753));
	notech_inv i_52288(.A(n_3849), .Z(n_42754));
	notech_inv i_52289(.A(\imm1[12] ), .Z(n_42756));
	notech_inv i_52290(.A(n_3848), .Z(n_42757));
	notech_inv i_52291(.A(\imm1[13] ), .Z(n_42759));
	notech_inv i_52292(.A(n_3847), .Z(n_42760));
	notech_inv i_52293(.A(\imm1[14] ), .Z(n_42761));
	notech_inv i_52294(.A(n_3846), .Z(n_42762));
	notech_inv i_52295(.A(\imm1[15] ), .Z(n_42763));
	notech_inv i_52296(.A(n_3845), .Z(n_42764));
	notech_inv i_52297(.A(\imm1[16] ), .Z(n_42765));
	notech_inv i_52298(.A(n_3844), .Z(n_42766));
	notech_inv i_52299(.A(\imm1[17] ), .Z(n_42767));
	notech_inv i_52300(.A(n_3843), .Z(n_42768));
	notech_inv i_52301(.A(\imm1[18] ), .Z(n_42769));
	notech_inv i_52302(.A(n_3842), .Z(n_42770));
	notech_inv i_52303(.A(\imm1[19] ), .Z(n_42771));
	notech_inv i_52304(.A(n_3841), .Z(n_42773));
	notech_inv i_52305(.A(\imm1[20] ), .Z(n_42774));
	notech_inv i_52306(.A(n_3840), .Z(n_42775));
	notech_inv i_52307(.A(\imm1[21] ), .Z(n_42776));
	notech_inv i_52308(.A(n_3839), .Z(n_42777));
	notech_inv i_52309(.A(\imm1[22] ), .Z(n_42779));
	notech_inv i_52310(.A(n_3838), .Z(n_42780));
	notech_inv i_52311(.A(\imm1[23] ), .Z(n_42781));
	notech_inv i_52312(.A(n_3837), .Z(n_42782));
	notech_inv i_52313(.A(\imm1[24] ), .Z(n_42783));
	notech_inv i_52314(.A(n_3836), .Z(n_42785));
	notech_inv i_52315(.A(\imm1[25] ), .Z(n_42786));
	notech_inv i_52316(.A(n_45809), .Z(n_42787));
	notech_inv i_52317(.A(\imm1[26] ), .Z(n_42788));
	notech_inv i_52318(.A(n_3835), .Z(n_42789));
	notech_inv i_52319(.A(\imm1[27] ), .Z(n_42791));
	notech_inv i_52320(.A(n_3834), .Z(n_42792));
	notech_inv i_52321(.A(\imm1[28] ), .Z(n_42793));
	notech_inv i_52322(.A(n_3833), .Z(n_42794));
	notech_inv i_52323(.A(\imm1[29] ), .Z(n_42795));
	notech_inv i_52324(.A(n_3832), .Z(n_42797));
	notech_inv i_52325(.A(\imm1[30] ), .Z(n_42798));
	notech_inv i_52326(.A(n_3831), .Z(n_42799));
	notech_inv i_52327(.A(\imm1[31] ), .Z(n_42800));
	notech_inv i_52328(.A(n_3830), .Z(n_42801));
	notech_inv i_52329(.A(\imm1[32] ), .Z(n_42803));
	notech_inv i_52330(.A(n_3829), .Z(n_42804));
	notech_inv i_52331(.A(\imm1[33] ), .Z(n_42805));
	notech_inv i_52332(.A(n_3828), .Z(n_42806));
	notech_inv i_52333(.A(\imm1[34] ), .Z(n_42807));
	notech_inv i_52334(.A(n_3827), .Z(n_42809));
	notech_inv i_52335(.A(\imm1[35] ), .Z(n_42810));
	notech_inv i_52336(.A(n_3826), .Z(n_42811));
	notech_inv i_52337(.A(\imm1[36] ), .Z(n_42812));
	notech_inv i_52338(.A(n_3825), .Z(n_42813));
	notech_inv i_52339(.A(\imm1[37] ), .Z(n_42815));
	notech_inv i_52340(.A(n_3824), .Z(n_42816));
	notech_inv i_52341(.A(\imm1[38] ), .Z(n_42817));
	notech_inv i_52342(.A(n_3823), .Z(n_42818));
	notech_inv i_52343(.A(\imm1[39] ), .Z(n_42819));
	notech_inv i_52344(.A(n_3822), .Z(n_42821));
	notech_inv i_52345(.A(\imm1[40] ), .Z(n_42822));
	notech_inv i_52346(.A(n_3821), .Z(n_42823));
	notech_inv i_52347(.A(\imm1[41] ), .Z(n_42824));
	notech_inv i_52348(.A(n_3820), .Z(n_42825));
	notech_inv i_52349(.A(\imm1[42] ), .Z(n_42827));
	notech_inv i_52350(.A(n_3819), .Z(n_42828));
	notech_inv i_52351(.A(\imm1[43] ), .Z(n_42829));
	notech_inv i_52352(.A(n_3818), .Z(n_42830));
	notech_inv i_52353(.A(\imm1[44] ), .Z(n_42831));
	notech_inv i_52354(.A(n_3817), .Z(n_42833));
	notech_inv i_52355(.A(\imm1[45] ), .Z(n_42834));
	notech_inv i_52356(.A(n_3816), .Z(n_42835));
	notech_inv i_52357(.A(\imm1[46] ), .Z(n_42836));
	notech_inv i_52358(.A(n_3815), .Z(n_42837));
	notech_inv i_52359(.A(\imm1[47] ), .Z(n_42839));
	notech_inv i_52360(.A(n_3814), .Z(n_42840));
	notech_inv i_52361(.A(inst_deco2[0]), .Z(n_42841));
	notech_inv i_52362(.A(n_3813), .Z(n_42842));
	notech_inv i_52363(.A(inst_deco2[1]), .Z(n_42843));
	notech_inv i_52364(.A(inst_deco2[2]), .Z(n_42845));
	notech_inv i_52365(.A(n_3812), .Z(n_42846));
	notech_inv i_52366(.A(inst_deco2[3]), .Z(n_42847));
	notech_inv i_52367(.A(inst_deco2[4]), .Z(n_42848));
	notech_inv i_52368(.A(n_3811), .Z(n_42849));
	notech_inv i_52369(.A(inst_deco2[5]), .Z(n_42851));
	notech_inv i_52370(.A(n_3810), .Z(n_42852));
	notech_inv i_52371(.A(inst_deco2[6]), .Z(n_42853));
	notech_inv i_52372(.A(n_3809), .Z(n_42854));
	notech_inv i_52373(.A(inst_deco2[7]), .Z(n_42855));
	notech_inv i_52374(.A(n_3808), .Z(n_42857));
	notech_inv i_52375(.A(inst_deco2[8]), .Z(n_42858));
	notech_inv i_52376(.A(inst_deco2[9]), .Z(n_42859));
	notech_inv i_52377(.A(n_3807), .Z(n_42860));
	notech_inv i_52378(.A(inst_deco2[10]), .Z(n_42861));
	notech_inv i_52379(.A(inst_deco2[11]), .Z(n_42863));
	notech_inv i_52380(.A(n_3806), .Z(n_42864));
	notech_inv i_52381(.A(inst_deco2[12]), .Z(n_42865));
	notech_inv i_52382(.A(inst_deco2[13]), .Z(n_42866));
	notech_inv i_52383(.A(n_3805), .Z(n_42867));
	notech_inv i_52384(.A(inst_deco2[14]), .Z(n_42869));
	notech_inv i_52385(.A(inst_deco2[15]), .Z(n_42870));
	notech_inv i_52386(.A(n_3804), .Z(n_42871));
	notech_inv i_52387(.A(inst_deco2[16]), .Z(n_42872));
	notech_inv i_52388(.A(inst_deco2[17]), .Z(n_42873));
	notech_inv i_52389(.A(n_3803), .Z(n_42875));
	notech_inv i_52390(.A(inst_deco2[18]), .Z(n_42876));
	notech_inv i_52391(.A(inst_deco2[19]), .Z(n_42877));
	notech_inv i_52392(.A(n_3802), .Z(n_42878));
	notech_inv i_52393(.A(inst_deco2[20]), .Z(n_42879));
	notech_inv i_52394(.A(inst_deco2[21]), .Z(n_42881));
	notech_inv i_52395(.A(n_3801), .Z(n_42882));
	notech_inv i_52396(.A(inst_deco2[22]), .Z(n_42883));
	notech_inv i_52397(.A(inst_deco2[23]), .Z(n_42884));
	notech_inv i_52398(.A(n_3800), .Z(n_42885));
	notech_inv i_52399(.A(inst_deco2[24]), .Z(n_42887));
	notech_inv i_52400(.A(inst_deco2[25]), .Z(n_42888));
	notech_inv i_52401(.A(n_3799), .Z(n_42889));
	notech_inv i_52402(.A(inst_deco2[26]), .Z(n_42890));
	notech_inv i_52403(.A(inst_deco2[27]), .Z(n_42891));
	notech_inv i_52404(.A(n_3798), .Z(n_42893));
	notech_inv i_52405(.A(inst_deco2[28]), .Z(n_42894));
	notech_inv i_52406(.A(inst_deco2[29]), .Z(n_42895));
	notech_inv i_52407(.A(n_3797), .Z(n_42896));
	notech_inv i_52408(.A(inst_deco2[30]), .Z(n_42897));
	notech_inv i_52409(.A(inst_deco2[31]), .Z(n_42899));
	notech_inv i_52410(.A(n_3796), .Z(n_42900));
	notech_inv i_52411(.A(inst_deco2[32]), .Z(n_42901));
	notech_inv i_52412(.A(inst_deco2[33]), .Z(n_42902));
	notech_inv i_52413(.A(n_3794), .Z(n_42903));
	notech_inv i_52414(.A(inst_deco2[34]), .Z(n_42905));
	notech_inv i_52415(.A(inst_deco2[35]), .Z(n_42906));
	notech_inv i_52416(.A(n_3792), .Z(n_42907));
	notech_inv i_52417(.A(inst_deco2[36]), .Z(n_42908));
	notech_inv i_52418(.A(inst_deco2[37]), .Z(n_42909));
	notech_inv i_52419(.A(n_3790), .Z(n_42911));
	notech_inv i_52420(.A(inst_deco2[38]), .Z(n_42912));
	notech_inv i_52421(.A(inst_deco2[39]), .Z(n_42913));
	notech_inv i_52422(.A(n_3788), .Z(n_42914));
	notech_inv i_52423(.A(inst_deco2[40]), .Z(n_42915));
	notech_inv i_52424(.A(n_3786), .Z(n_42917));
	notech_inv i_52425(.A(inst_deco2[41]), .Z(n_42918));
	notech_inv i_52426(.A(n_3784), .Z(n_42919));
	notech_inv i_52427(.A(inst_deco2[42]), .Z(n_42920));
	notech_inv i_52428(.A(n_3782), .Z(n_42921));
	notech_inv i_52429(.A(inst_deco2[43]), .Z(n_42923));
	notech_inv i_52430(.A(n_3780), .Z(n_42924));
	notech_inv i_52431(.A(inst_deco2[44]), .Z(n_42925));
	notech_inv i_52432(.A(n_3778), .Z(n_42926));
	notech_inv i_52433(.A(inst_deco2[45]), .Z(n_42927));
	notech_inv i_52434(.A(inst_deco2[46]), .Z(n_42929));
	notech_inv i_52435(.A(n_3776), .Z(n_42930));
	notech_inv i_52436(.A(inst_deco2[47]), .Z(n_42931));
	notech_inv i_52437(.A(inst_deco2[48]), .Z(n_42932));
	notech_inv i_52438(.A(n_3774), .Z(n_42933));
	notech_inv i_52439(.A(inst_deco2[49]), .Z(n_42935));
	notech_inv i_52440(.A(inst_deco2[50]), .Z(n_42936));
	notech_inv i_52441(.A(n_3772), .Z(n_42937));
	notech_inv i_52442(.A(inst_deco2[51]), .Z(n_42938));
	notech_inv i_52443(.A(inst_deco2[52]), .Z(n_42939));
	notech_inv i_52444(.A(n_3770), .Z(n_42941));
	notech_inv i_52445(.A(inst_deco2[53]), .Z(n_42942));
	notech_inv i_52446(.A(inst_deco2[54]), .Z(n_42943));
	notech_inv i_52447(.A(n_3768), .Z(n_42944));
	notech_inv i_52448(.A(inst_deco2[55]), .Z(n_42945));
	notech_inv i_52449(.A(inst_deco2[56]), .Z(n_42947));
	notech_inv i_52450(.A(n_3766), .Z(n_42948));
	notech_inv i_52451(.A(inst_deco2[57]), .Z(n_42949));
	notech_inv i_52452(.A(inst_deco2[58]), .Z(n_42950));
	notech_inv i_52453(.A(n_3764), .Z(n_42951));
	notech_inv i_52454(.A(inst_deco2[59]), .Z(n_42953));
	notech_inv i_52455(.A(inst_deco2[60]), .Z(n_42954));
	notech_inv i_52456(.A(n_3762), .Z(n_42955));
	notech_inv i_52457(.A(inst_deco2[61]), .Z(n_42956));
	notech_inv i_52458(.A(inst_deco2[62]), .Z(n_42957));
	notech_inv i_52459(.A(n_3760), .Z(n_42959));
	notech_inv i_52460(.A(inst_deco2[63]), .Z(n_42960));
	notech_inv i_52461(.A(inst_deco2[64]), .Z(n_42961));
	notech_inv i_52462(.A(n_3758), .Z(n_42962));
	notech_inv i_52463(.A(inst_deco2[65]), .Z(n_42963));
	notech_inv i_52464(.A(inst_deco2[66]), .Z(n_42965));
	notech_inv i_52465(.A(n_3756), .Z(n_42966));
	notech_inv i_52466(.A(inst_deco2[67]), .Z(n_42967));
	notech_inv i_52467(.A(inst_deco2[68]), .Z(n_42968));
	notech_inv i_52468(.A(n_3754), .Z(n_42969));
	notech_inv i_52469(.A(inst_deco2[69]), .Z(n_42971));
	notech_inv i_52470(.A(inst_deco2[70]), .Z(n_42972));
	notech_inv i_52471(.A(n_3752), .Z(n_42973));
	notech_inv i_52472(.A(inst_deco2[71]), .Z(n_42974));
	notech_inv i_52473(.A(inst_deco2[72]), .Z(n_42975));
	notech_inv i_52474(.A(n_3750), .Z(n_42977));
	notech_inv i_52475(.A(inst_deco2[73]), .Z(n_42978));
	notech_inv i_52476(.A(inst_deco2[74]), .Z(n_42979));
	notech_inv i_52477(.A(n_3748), .Z(n_42980));
	notech_inv i_52478(.A(inst_deco2[75]), .Z(n_42981));
	notech_inv i_52479(.A(inst_deco2[76]), .Z(n_42983));
	notech_inv i_52480(.A(n_3746), .Z(n_42984));
	notech_inv i_52481(.A(inst_deco2[77]), .Z(n_42985));
	notech_inv i_52482(.A(inst_deco2[78]), .Z(n_42986));
	notech_inv i_52483(.A(n_3744), .Z(n_42987));
	notech_inv i_52484(.A(inst_deco2[79]), .Z(n_42989));
	notech_inv i_52485(.A(inst_deco2[80]), .Z(n_42990));
	notech_inv i_52486(.A(n_3742), .Z(n_42991));
	notech_inv i_52487(.A(inst_deco2[81]), .Z(n_42992));
	notech_inv i_52488(.A(inst_deco2[82]), .Z(n_42993));
	notech_inv i_52489(.A(n_3740), .Z(n_42995));
	notech_inv i_52490(.A(inst_deco2[83]), .Z(n_42996));
	notech_inv i_52491(.A(inst_deco2[84]), .Z(n_42997));
	notech_inv i_52492(.A(n_3738), .Z(n_42998));
	notech_inv i_52493(.A(inst_deco2[85]), .Z(n_42999));
	notech_inv i_52494(.A(inst_deco2[86]), .Z(n_43001));
	notech_inv i_52495(.A(n_3736), .Z(n_43002));
	notech_inv i_52496(.A(inst_deco2[87]), .Z(n_43003));
	notech_inv i_52497(.A(inst_deco2[88]), .Z(n_43004));
	notech_inv i_52498(.A(n_3734), .Z(n_43005));
	notech_inv i_52499(.A(inst_deco2[89]), .Z(n_43007));
	notech_inv i_52500(.A(inst_deco2[90]), .Z(n_43008));
	notech_inv i_52501(.A(n_3732), .Z(n_43009));
	notech_inv i_52502(.A(inst_deco2[91]), .Z(n_43010));
	notech_inv i_52503(.A(inst_deco2[92]), .Z(n_43011));
	notech_inv i_52504(.A(n_3730), .Z(n_43013));
	notech_inv i_52505(.A(inst_deco2[93]), .Z(n_43014));
	notech_inv i_52506(.A(inst_deco2[94]), .Z(n_43015));
	notech_inv i_52507(.A(n_3728), .Z(n_43016));
	notech_inv i_52508(.A(inst_deco2[95]), .Z(n_43017));
	notech_inv i_52509(.A(inst_deco2[96]), .Z(n_43019));
	notech_inv i_52510(.A(n_3726), .Z(n_43020));
	notech_inv i_52511(.A(inst_deco2[97]), .Z(n_43021));
	notech_inv i_52512(.A(inst_deco2[98]), .Z(n_43022));
	notech_inv i_52513(.A(n_3724), .Z(n_43023));
	notech_inv i_52514(.A(inst_deco2[99]), .Z(n_43025));
	notech_inv i_52515(.A(inst_deco2[100]), .Z(n_43026));
	notech_inv i_52516(.A(n_3722), .Z(n_43027));
	notech_inv i_52517(.A(inst_deco2[101]), .Z(n_43028));
	notech_inv i_52518(.A(inst_deco2[102]), .Z(n_43029));
	notech_inv i_52519(.A(n_3720), .Z(n_43031));
	notech_inv i_52520(.A(n_42498), .Z(n_43032));
	notech_inv i_52521(.A(inst_deco2[103]), .Z(n_43033));
	notech_inv i_52522(.A(inst_deco2[104]), .Z(n_43034));
	notech_inv i_52523(.A(n_3718), .Z(n_43035));
	notech_inv i_52524(.A(inst_deco2[105]), .Z(n_43037));
	notech_inv i_52525(.A(inst_deco2[106]), .Z(n_43038));
	notech_inv i_52526(.A(n_3716), .Z(n_43039));
	notech_inv i_52527(.A(inst_deco2[107]), .Z(n_43040));
	notech_inv i_52528(.A(inst_deco2[108]), .Z(n_43041));
	notech_inv i_52529(.A(n_3714), .Z(n_43043));
	notech_inv i_52530(.A(inst_deco2[109]), .Z(n_43044));
	notech_inv i_52531(.A(inst_deco2[110]), .Z(n_43045));
	notech_inv i_52532(.A(n_3712), .Z(n_43046));
	notech_inv i_52533(.A(inst_deco2[111]), .Z(n_43047));
	notech_inv i_52534(.A(inst_deco2[112]), .Z(n_43049));
	notech_inv i_52535(.A(n_3710), .Z(n_43050));
	notech_inv i_52536(.A(inst_deco2[113]), .Z(n_43051));
	notech_inv i_52537(.A(inst_deco2[114]), .Z(n_43052));
	notech_inv i_52538(.A(n_3708), .Z(n_43053));
	notech_inv i_52539(.A(inst_deco2[115]), .Z(n_43055));
	notech_inv i_52540(.A(inst_deco2[116]), .Z(n_43056));
	notech_inv i_52541(.A(n_3706), .Z(n_43057));
	notech_inv i_52542(.A(inst_deco2[117]), .Z(n_43058));
	notech_inv i_52543(.A(inst_deco2[118]), .Z(n_43059));
	notech_inv i_52544(.A(n_3704), .Z(n_43061));
	notech_inv i_52545(.A(inst_deco2[119]), .Z(n_43062));
	notech_inv i_52546(.A(inst_deco2[120]), .Z(n_43063));
	notech_inv i_52547(.A(n_3702), .Z(n_43064));
	notech_inv i_52548(.A(inst_deco2[121]), .Z(n_43065));
	notech_inv i_52549(.A(inst_deco2[122]), .Z(n_43067));
	notech_inv i_52550(.A(n_3700), .Z(n_43068));
	notech_inv i_52551(.A(inst_deco2[123]), .Z(n_43069));
	notech_inv i_52552(.A(inst_deco2[124]), .Z(n_43070));
	notech_inv i_52553(.A(n_3698), .Z(n_43071));
	notech_inv i_52554(.A(inst_deco2[125]), .Z(n_43073));
	notech_inv i_52555(.A(inst_deco2[126]), .Z(n_43074));
	notech_inv i_52556(.A(n_3696), .Z(n_43075));
	notech_inv i_52557(.A(inst_deco2[127]), .Z(n_43076));
	notech_inv i_52558(.A(n_49895), .Z(n_43077));
	notech_inv i_52559(.A(inst_deco1[0]), .Z(n_43079));
	notech_inv i_52560(.A(n_3694), .Z(n_43080));
	notech_inv i_52561(.A(inst_deco1[1]), .Z(n_43081));
	notech_inv i_52562(.A(n_3692), .Z(n_43082));
	notech_inv i_52563(.A(inst_deco1[2]), .Z(n_43083));
	notech_inv i_52564(.A(n_3690), .Z(n_43085));
	notech_inv i_52565(.A(inst_deco1[3]), .Z(n_43086));
	notech_inv i_52566(.A(n_3688), .Z(n_43087));
	notech_inv i_52567(.A(inst_deco1[4]), .Z(n_43088));
	notech_inv i_52568(.A(n_3686), .Z(n_43089));
	notech_inv i_52569(.A(n_49925), .Z(n_43091));
	notech_inv i_52570(.A(inst_deco1[5]), .Z(n_43092));
	notech_inv i_52571(.A(n_3684), .Z(n_43093));
	notech_inv i_52572(.A(inst_deco1[6]), .Z(n_43094));
	notech_inv i_52573(.A(n_49937), .Z(n_43095));
	notech_inv i_52574(.A(inst_deco1[7]), .Z(n_43097));
	notech_inv i_52575(.A(n_3682), .Z(n_43098));
	notech_inv i_52576(.A(n_49943), .Z(n_43099));
	notech_inv i_52577(.A(inst_deco1[8]), .Z(n_43100));
	notech_inv i_52578(.A(n_3680), .Z(n_43101));
	notech_inv i_52579(.A(inst_deco1[9]), .Z(n_43103));
	notech_inv i_52580(.A(n_3678), .Z(n_43104));
	notech_inv i_52581(.A(inst_deco1[10]), .Z(n_43105));
	notech_inv i_52582(.A(n_3676), .Z(n_43106));
	notech_inv i_52583(.A(inst_deco1[11]), .Z(n_43107));
	notech_inv i_52584(.A(n_3674), .Z(n_43109));
	notech_inv i_52585(.A(inst_deco1[12]), .Z(n_43110));
	notech_inv i_52586(.A(n_3672), .Z(n_43111));
	notech_inv i_52587(.A(inst_deco1[13]), .Z(n_43112));
	notech_inv i_52588(.A(n_3670), .Z(n_43113));
	notech_inv i_52589(.A(inst_deco1[14]), .Z(n_43115));
	notech_inv i_52590(.A(n_3669), .Z(n_43116));
	notech_inv i_52591(.A(inst_deco1[15]), .Z(n_43117));
	notech_inv i_52592(.A(n_3668), .Z(n_43118));
	notech_inv i_52593(.A(inst_deco1[16]), .Z(n_43119));
	notech_inv i_52594(.A(n_3667), .Z(n_43121));
	notech_inv i_52595(.A(n_3666), .Z(n_43122));
	notech_inv i_52596(.A(inst_deco1[18]), .Z(n_43123));
	notech_inv i_52597(.A(n_3665), .Z(n_43124));
	notech_inv i_52598(.A(inst_deco1[19]), .Z(n_43125));
	notech_inv i_52599(.A(n_3664), .Z(n_43127));
	notech_inv i_52600(.A(inst_deco1[20]), .Z(n_43128));
	notech_inv i_52601(.A(n_3663), .Z(n_43129));
	notech_inv i_52602(.A(n_3662), .Z(n_43130));
	notech_inv i_52603(.A(inst_deco1[22]), .Z(n_43131));
	notech_inv i_52604(.A(n_3661), .Z(n_43133));
	notech_inv i_52605(.A(inst_deco1[23]), .Z(n_43134));
	notech_inv i_52606(.A(n_3660), .Z(n_43135));
	notech_inv i_52607(.A(inst_deco1[24]), .Z(n_43136));
	notech_inv i_52608(.A(n_3659), .Z(n_43137));
	notech_inv i_52609(.A(inst_deco1[25]), .Z(n_43139));
	notech_inv i_52610(.A(n_3658), .Z(n_43140));
	notech_inv i_52611(.A(inst_deco1[26]), .Z(n_43141));
	notech_inv i_52612(.A(n_3657), .Z(n_43142));
	notech_inv i_52613(.A(inst_deco1[27]), .Z(n_43143));
	notech_inv i_52614(.A(n_3656), .Z(n_43145));
	notech_inv i_52615(.A(inst_deco1[28]), .Z(n_43146));
	notech_inv i_52616(.A(n_3655), .Z(n_43147));
	notech_inv i_52617(.A(inst_deco1[29]), .Z(n_43148));
	notech_inv i_52618(.A(n_3654), .Z(n_43149));
	notech_inv i_52619(.A(inst_deco1[30]), .Z(n_43151));
	notech_inv i_52620(.A(n_3653), .Z(n_43152));
	notech_inv i_52621(.A(inst_deco1[31]), .Z(n_43153));
	notech_inv i_52622(.A(n_3652), .Z(n_43154));
	notech_inv i_52623(.A(inst_deco1[32]), .Z(n_43155));
	notech_inv i_52624(.A(n_3651), .Z(n_43157));
	notech_inv i_52625(.A(inst_deco1[33]), .Z(n_43158));
	notech_inv i_52626(.A(n_3650), .Z(n_43159));
	notech_inv i_52627(.A(inst_deco1[34]), .Z(n_43160));
	notech_inv i_52628(.A(n_3649), .Z(n_43161));
	notech_inv i_52629(.A(inst_deco1[35]), .Z(n_43163));
	notech_inv i_52630(.A(n_3648), .Z(n_43164));
	notech_inv i_52631(.A(inst_deco1[36]), .Z(n_43165));
	notech_inv i_52632(.A(n_3647), .Z(n_43166));
	notech_inv i_52633(.A(inst_deco1[37]), .Z(n_43167));
	notech_inv i_52634(.A(n_3646), .Z(n_43169));
	notech_inv i_52635(.A(inst_deco1[38]), .Z(n_43170));
	notech_inv i_52636(.A(n_3645), .Z(n_43171));
	notech_inv i_52637(.A(inst_deco1[39]), .Z(n_43172));
	notech_inv i_52638(.A(n_3644), .Z(n_43173));
	notech_inv i_52639(.A(inst_deco1[40]), .Z(n_43175));
	notech_inv i_52640(.A(n_50141), .Z(n_43176));
	notech_inv i_52641(.A(inst_deco1[41]), .Z(n_43177));
	notech_inv i_52642(.A(n_3643), .Z(n_43178));
	notech_inv i_52643(.A(n_50147), .Z(n_43179));
	notech_inv i_52644(.A(inst_deco1[42]), .Z(n_43181));
	notech_inv i_52645(.A(n_50153), .Z(n_43182));
	notech_inv i_52646(.A(inst_deco1[43]), .Z(n_43183));
	notech_inv i_52647(.A(n_3642), .Z(n_43184));
	notech_inv i_52648(.A(n_50159), .Z(n_43185));
	notech_inv i_52649(.A(inst_deco1[44]), .Z(n_43187));
	notech_inv i_52650(.A(n_50165), .Z(n_43188));
	notech_inv i_52651(.A(inst_deco1[45]), .Z(n_43189));
	notech_inv i_52652(.A(n_3641), .Z(n_43190));
	notech_inv i_52653(.A(inst_deco1[46]), .Z(n_43191));
	notech_inv i_52654(.A(n_3640), .Z(n_43193));
	notech_inv i_52655(.A(inst_deco1[47]), .Z(n_43194));
	notech_inv i_52656(.A(n_3639), .Z(n_43195));
	notech_inv i_52657(.A(inst_deco1[48]), .Z(n_43196));
	notech_inv i_52658(.A(n_3638), .Z(n_43197));
	notech_inv i_52659(.A(inst_deco1[49]), .Z(n_43199));
	notech_inv i_52660(.A(n_3637), .Z(n_43200));
	notech_inv i_52661(.A(inst_deco1[50]), .Z(n_43201));
	notech_inv i_52662(.A(n_3636), .Z(n_43202));
	notech_inv i_52663(.A(inst_deco1[51]), .Z(n_43203));
	notech_inv i_52664(.A(n_3635), .Z(n_43205));
	notech_inv i_52665(.A(inst_deco1[52]), .Z(n_43206));
	notech_inv i_52666(.A(n_3634), .Z(n_43207));
	notech_inv i_52667(.A(inst_deco1[53]), .Z(n_43208));
	notech_inv i_52668(.A(n_3633), .Z(n_43209));
	notech_inv i_52669(.A(inst_deco1[54]), .Z(n_43211));
	notech_inv i_52670(.A(n_3632), .Z(n_43212));
	notech_inv i_52671(.A(inst_deco1[55]), .Z(n_43213));
	notech_inv i_52672(.A(n_3631), .Z(n_43214));
	notech_inv i_52673(.A(inst_deco1[56]), .Z(n_43215));
	notech_inv i_52674(.A(n_3630), .Z(n_43217));
	notech_inv i_52675(.A(inst_deco1[57]), .Z(n_43218));
	notech_inv i_52676(.A(n_3629), .Z(n_43219));
	notech_inv i_52677(.A(inst_deco1[58]), .Z(n_43220));
	notech_inv i_52678(.A(n_3628), .Z(n_43221));
	notech_inv i_52679(.A(inst_deco1[59]), .Z(n_43223));
	notech_inv i_52680(.A(n_3627), .Z(n_43224));
	notech_inv i_52681(.A(inst_deco1[60]), .Z(n_43225));
	notech_inv i_52682(.A(n_3626), .Z(n_43226));
	notech_inv i_52683(.A(inst_deco1[61]), .Z(n_43227));
	notech_inv i_52684(.A(n_3625), .Z(n_43229));
	notech_inv i_52685(.A(inst_deco1[62]), .Z(n_43230));
	notech_inv i_52686(.A(n_3624), .Z(n_43231));
	notech_inv i_52687(.A(inst_deco1[63]), .Z(n_43232));
	notech_inv i_52688(.A(n_3623), .Z(n_43233));
	notech_inv i_52689(.A(inst_deco1[64]), .Z(n_43235));
	notech_inv i_52690(.A(n_3622), .Z(n_43236));
	notech_inv i_52691(.A(inst_deco1[65]), .Z(n_43237));
	notech_inv i_52692(.A(n_3621), .Z(n_43238));
	notech_inv i_52693(.A(inst_deco1[66]), .Z(n_43239));
	notech_inv i_52694(.A(n_3620), .Z(n_43241));
	notech_inv i_52695(.A(inst_deco1[67]), .Z(n_43242));
	notech_inv i_52696(.A(n_3619), .Z(n_43243));
	notech_inv i_52697(.A(inst_deco1[68]), .Z(n_43244));
	notech_inv i_52698(.A(n_3618), .Z(n_43245));
	notech_inv i_52699(.A(inst_deco1[69]), .Z(n_43247));
	notech_inv i_52700(.A(n_3617), .Z(n_43248));
	notech_inv i_52701(.A(inst_deco1[70]), .Z(n_43249));
	notech_inv i_52702(.A(n_3616), .Z(n_43250));
	notech_inv i_52703(.A(inst_deco1[71]), .Z(n_43251));
	notech_inv i_52704(.A(n_3615), .Z(n_43253));
	notech_inv i_52705(.A(inst_deco1[72]), .Z(n_43254));
	notech_inv i_52706(.A(n_3614), .Z(n_43255));
	notech_inv i_52707(.A(inst_deco1[73]), .Z(n_43256));
	notech_inv i_52708(.A(n_3613), .Z(n_43257));
	notech_inv i_52709(.A(inst_deco1[74]), .Z(n_43259));
	notech_inv i_52710(.A(n_3612), .Z(n_43260));
	notech_inv i_52711(.A(inst_deco1[75]), .Z(n_43261));
	notech_inv i_52712(.A(n_3611), .Z(n_43262));
	notech_inv i_52713(.A(inst_deco1[76]), .Z(n_43263));
	notech_inv i_52714(.A(n_3610), .Z(n_43265));
	notech_inv i_52715(.A(inst_deco1[77]), .Z(n_43266));
	notech_inv i_52716(.A(n_3609), .Z(n_43267));
	notech_inv i_52717(.A(inst_deco1[78]), .Z(n_43268));
	notech_inv i_52718(.A(n_3608), .Z(n_43269));
	notech_inv i_52719(.A(inst_deco1[79]), .Z(n_43271));
	notech_inv i_52720(.A(n_3607), .Z(n_43272));
	notech_inv i_52721(.A(n_3606), .Z(n_43273));
	notech_inv i_52722(.A(n_3605), .Z(n_43274));
	notech_inv i_52723(.A(n_3603), .Z(n_43275));
	notech_inv i_52724(.A(n_3601), .Z(n_43277));
	notech_inv i_52725(.A(n_3599), .Z(n_43278));
	notech_inv i_52726(.A(n_3597), .Z(n_43279));
	notech_inv i_52727(.A(n_3595), .Z(n_43280));
	notech_inv i_52728(.A(n_3593), .Z(n_43281));
	notech_inv i_52729(.A(inst_deco1[88]), .Z(n_43283));
	notech_inv i_52730(.A(n_3591), .Z(n_43284));
	notech_inv i_52731(.A(inst_deco1[89]), .Z(n_43285));
	notech_inv i_52732(.A(n_3589), .Z(n_43286));
	notech_inv i_52733(.A(inst_deco1[90]), .Z(n_43287));
	notech_inv i_52734(.A(n_3587), .Z(n_43289));
	notech_inv i_52735(.A(inst_deco1[91]), .Z(n_43290));
	notech_inv i_52736(.A(n_3585), .Z(n_43291));
	notech_inv i_52737(.A(inst_deco1[92]), .Z(n_43292));
	notech_inv i_52738(.A(n_3583), .Z(n_43293));
	notech_inv i_52739(.A(inst_deco1[93]), .Z(n_43295));
	notech_inv i_52740(.A(n_3581), .Z(n_43296));
	notech_inv i_52741(.A(inst_deco1[94]), .Z(n_43297));
	notech_inv i_52742(.A(n_3579), .Z(n_43298));
	notech_inv i_52743(.A(inst_deco1[95]), .Z(n_43299));
	notech_inv i_52744(.A(n_3577), .Z(n_43301));
	notech_inv i_52745(.A(inst_deco1[96]), .Z(n_43302));
	notech_inv i_52746(.A(n_3576), .Z(n_43303));
	notech_inv i_52747(.A(inst_deco1[97]), .Z(n_43304));
	notech_inv i_52748(.A(n_3575), .Z(n_43305));
	notech_inv i_52749(.A(inst_deco1[98]), .Z(n_43307));
	notech_inv i_52750(.A(n_3573), .Z(n_43308));
	notech_inv i_52751(.A(inst_deco1[99]), .Z(n_43309));
	notech_inv i_52752(.A(n_3572), .Z(n_43310));
	notech_inv i_52753(.A(inst_deco1[100]), .Z(n_43311));
	notech_inv i_52754(.A(n_3571), .Z(n_43313));
	notech_inv i_52755(.A(inst_deco1[101]), .Z(n_43314));
	notech_inv i_52756(.A(n_3570), .Z(n_43315));
	notech_inv i_52757(.A(inst_deco1[102]), .Z(n_43316));
	notech_inv i_52758(.A(n_3569), .Z(n_43317));
	notech_inv i_52759(.A(inst_deco1[103]), .Z(n_43319));
	notech_inv i_52760(.A(n_3568), .Z(n_43320));
	notech_inv i_52761(.A(inst_deco1[104]), .Z(n_43321));
	notech_inv i_52762(.A(n_3567), .Z(n_43322));
	notech_inv i_52763(.A(inst_deco1[105]), .Z(n_43323));
	notech_inv i_52764(.A(n_3566), .Z(n_43325));
	notech_inv i_52765(.A(n_3565), .Z(n_43326));
	notech_inv i_52766(.A(inst_deco1[107]), .Z(n_43327));
	notech_inv i_52767(.A(n_3564), .Z(n_43328));
	notech_inv i_52768(.A(inst_deco1[108]), .Z(n_43329));
	notech_inv i_52769(.A(n_3563), .Z(n_43331));
	notech_inv i_52770(.A(inst_deco1[109]), .Z(n_43332));
	notech_inv i_52771(.A(n_3562), .Z(n_43333));
	notech_inv i_52772(.A(inst_deco1[110]), .Z(n_43334));
	notech_inv i_52773(.A(n_3561), .Z(n_43335));
	notech_inv i_52774(.A(inst_deco1[111]), .Z(n_43337));
	notech_inv i_52775(.A(n_3560), .Z(n_43338));
	notech_inv i_52776(.A(inst_deco1[112]), .Z(n_43339));
	notech_inv i_52777(.A(n_3559), .Z(n_43340));
	notech_inv i_52778(.A(n_3558), .Z(n_43341));
	notech_inv i_52779(.A(inst_deco1[114]), .Z(n_43343));
	notech_inv i_52780(.A(n_3557), .Z(n_43344));
	notech_inv i_52781(.A(inst_deco1[115]), .Z(n_43345));
	notech_inv i_52782(.A(n_3556), .Z(n_43346));
	notech_inv i_52783(.A(inst_deco1[116]), .Z(n_43347));
	notech_inv i_52784(.A(n_3555), .Z(n_43349));
	notech_inv i_52785(.A(inst_deco1[117]), .Z(n_43350));
	notech_inv i_52786(.A(n_3554), .Z(n_43351));
	notech_inv i_52787(.A(inst_deco1[118]), .Z(n_43352));
	notech_inv i_52788(.A(n_3553), .Z(n_43353));
	notech_inv i_52789(.A(inst_deco1[119]), .Z(n_43355));
	notech_inv i_52790(.A(n_3552), .Z(n_43356));
	notech_inv i_52791(.A(inst_deco1[120]), .Z(n_43357));
	notech_inv i_52792(.A(n_3551), .Z(n_43358));
	notech_inv i_52793(.A(inst_deco1[121]), .Z(n_43359));
	notech_inv i_52794(.A(n_3550), .Z(n_43361));
	notech_inv i_52795(.A(inst_deco1[122]), .Z(n_43362));
	notech_inv i_52796(.A(n_3549), .Z(n_43363));
	notech_inv i_52797(.A(inst_deco1[123]), .Z(n_43364));
	notech_inv i_52798(.A(n_3548), .Z(n_43365));
	notech_inv i_52799(.A(inst_deco1[124]), .Z(n_43367));
	notech_inv i_52800(.A(n_3547), .Z(n_43368));
	notech_inv i_52801(.A(inst_deco1[125]), .Z(n_43369));
	notech_inv i_52802(.A(n_3546), .Z(n_43370));
	notech_inv i_52803(.A(inst_deco1[126]), .Z(n_43371));
	notech_inv i_52804(.A(n_3545), .Z(n_43373));
	notech_inv i_52805(.A(inst_deco1[127]), .Z(n_43374));
	notech_inv i_52806(.A(n_3544), .Z(n_43375));
	notech_inv i_52807(.A(n_3543), .Z(n_43376));
	notech_inv i_52808(.A(trig_itf), .Z(n_43377));
	notech_inv i_52809(.A(intf), .Z(n_43379));
	notech_inv i_52810(.A(n_3542), .Z(n_43380));
	notech_inv i_52811(.A(n_3541), .Z(n_43381));
	notech_inv i_52812(.A(n_3540), .Z(n_43382));
	notech_inv i_52813(.A(n_3539), .Z(n_43383));
	notech_inv i_52814(.A(n_3538), .Z(n_43385));
	notech_inv i_52815(.A(n_3537), .Z(n_43386));
	notech_inv i_52816(.A(n_3536), .Z(n_43387));
	notech_inv i_52817(.A(n_3535), .Z(n_43388));
	notech_inv i_52818(.A(n_3534), .Z(n_43389));
	notech_inv i_52819(.A(n_3533), .Z(n_43391));
	notech_inv i_52820(.A(n_3532), .Z(n_43392));
	notech_inv i_52821(.A(n_3531), .Z(n_43393));
	notech_inv i_52822(.A(n_3530), .Z(n_43394));
	notech_inv i_52823(.A(n_3529), .Z(n_43395));
	notech_inv i_52824(.A(n_3528), .Z(n_43397));
	notech_inv i_52825(.A(n_3527), .Z(n_43398));
	notech_inv i_52826(.A(ififo_rvect1[0]), .Z(n_43399));
	notech_inv i_52827(.A(n_3526), .Z(n_43400));
	notech_inv i_52828(.A(ififo_rvect1[1]), .Z(n_43401));
	notech_inv i_52829(.A(ififo_rvect1[2]), .Z(n_43403));
	notech_inv i_52830(.A(n_3525), .Z(n_43404));
	notech_inv i_52831(.A(ififo_rvect1[3]), .Z(n_43405));
	notech_inv i_52832(.A(ififo_rvect1[4]), .Z(n_43406));
	notech_inv i_52833(.A(n_3524), .Z(n_43407));
	notech_inv i_52834(.A(ififo_rvect1[5]), .Z(n_43409));
	notech_inv i_52835(.A(ififo_rvect1[6]), .Z(n_43410));
	notech_inv i_52836(.A(n_3523), .Z(n_43411));
	notech_inv i_52837(.A(ififo_rvect1[7]), .Z(n_43412));
	notech_inv i_52838(.A(n_3522), .Z(n_43413));
	notech_inv i_52839(.A(n_3521), .Z(n_43415));
	notech_inv i_52840(.A(n_3520), .Z(n_43416));
	notech_inv i_52841(.A(n_3519), .Z(n_43417));
	notech_inv i_52842(.A(n_3518), .Z(n_43418));
	notech_inv i_52843(.A(n_3517), .Z(n_43419));
	notech_inv i_52844(.A(n_3516), .Z(n_43421));
	notech_inv i_52845(.A(n_3515), .Z(n_43422));
	notech_inv i_52846(.A(n_3514), .Z(n_43423));
	notech_inv i_52847(.A(n_3513), .Z(n_43424));
	notech_inv i_52848(.A(n_3512), .Z(n_43425));
	notech_inv i_52849(.A(n_3511), .Z(n_43427));
	notech_inv i_52850(.A(i_ptr[2]), .Z(n_43428));
	notech_inv i_52851(.A(n_3510), .Z(n_43429));
	notech_inv i_52852(.A(n_3509), .Z(n_43430));
	notech_inv i_52853(.A(idx_deco[0]), .Z(n_43431));
	notech_inv i_52854(.A(n_3508), .Z(n_43433));
	notech_inv i_52855(.A(idx_deco[1]), .Z(n_43434));
	notech_inv i_52856(.A(n_3507), .Z(n_43435));
	notech_inv i_52857(.A(n_3506), .Z(n_43436));
	notech_inv i_52858(.A(fsm[1]), .Z(n_43437));
	notech_inv i_52859(.A(n_3505), .Z(n_43439));
	notech_inv i_52860(.A(n_3504), .Z(n_43440));
	notech_inv i_52861(.A(fsm[4]), .Z(n_43441));
	notech_inv i_52862(.A(n_3503), .Z(n_43442));
	notech_inv i_52863(.A(n_3502), .Z(n_43443));
	notech_inv i_52864(.A(repz), .Z(n_43445));
	notech_inv i_52865(.A(rep), .Z(n_43446));
	notech_inv i_52866(.A(n_3501), .Z(n_43447));
	notech_inv i_52867(.A(opz2[0]), .Z(n_43448));
	notech_inv i_52868(.A(opz2[1]), .Z(n_43449));
	notech_inv i_52869(.A(n_3500), .Z(n_43451));
	notech_inv i_52870(.A(n_3499), .Z(n_43452));
	notech_inv i_52871(.A(reps2[0]), .Z(n_43453));
	notech_inv i_52872(.A(reps2[1]), .Z(n_43454));
	notech_inv i_52873(.A(n_3498), .Z(n_43455));
	notech_inv i_52874(.A(reps2[2]), .Z(n_43457));
	notech_inv i_52875(.A(n_3497), .Z(n_43458));
	notech_inv i_52876(.A(reps1[0]), .Z(n_43459));
	notech_inv i_52877(.A(n_3496), .Z(n_43460));
	notech_inv i_52878(.A(reps1[1]), .Z(n_43461));
	notech_inv i_52879(.A(n_3495), .Z(n_43463));
	notech_inv i_52880(.A(reps1[2]), .Z(n_43464));
	notech_inv i_52881(.A(n_41609), .Z(n_43465));
	notech_inv i_52882(.A(overgs), .Z(n_43466));
	notech_inv i_52883(.A(n_3494), .Z(n_43467));
	notech_inv i_52884(.A(\over_seg2[5] ), .Z(n_43469));
	notech_inv i_52885(.A(n_3493), .Z(n_43470));
	notech_inv i_52886(.A(\over_seg1[5] ), .Z(n_43471));
	notech_inv i_52887(.A(n_3492), .Z(n_43472));
	notech_inv i_52888(.A(to_acu2[0]), .Z(n_43473));
	notech_inv i_52889(.A(to_acu2[1]), .Z(n_43475));
	notech_inv i_52890(.A(n_3491), .Z(n_43476));
	notech_inv i_52891(.A(to_acu2[2]), .Z(n_43477));
	notech_inv i_52892(.A(to_acu2[3]), .Z(n_43478));
	notech_inv i_52893(.A(n_3490), .Z(n_43479));
	notech_inv i_52894(.A(to_acu2[4]), .Z(n_43481));
	notech_inv i_52895(.A(to_acu2[5]), .Z(n_43482));
	notech_inv i_52896(.A(n_3489), .Z(n_43483));
	notech_inv i_52897(.A(to_acu2[6]), .Z(n_43484));
	notech_inv i_52898(.A(to_acu2[7]), .Z(n_43485));
	notech_inv i_52899(.A(n_3488), .Z(n_43487));
	notech_inv i_52900(.A(to_acu2[8]), .Z(n_43488));
	notech_inv i_52901(.A(to_acu2[9]), .Z(n_43489));
	notech_inv i_52902(.A(n_3487), .Z(n_43490));
	notech_inv i_52903(.A(to_acu2[10]), .Z(n_43491));
	notech_inv i_52904(.A(n_3486), .Z(n_43493));
	notech_inv i_52905(.A(to_acu2[11]), .Z(n_43494));
	notech_inv i_52906(.A(to_acu2[12]), .Z(n_43495));
	notech_inv i_52907(.A(n_3485), .Z(n_43496));
	notech_inv i_52908(.A(to_acu2[13]), .Z(n_43497));
	notech_inv i_52909(.A(to_acu2[14]), .Z(n_43499));
	notech_inv i_52910(.A(n_3484), .Z(n_43500));
	notech_inv i_52911(.A(to_acu2[15]), .Z(n_43501));
	notech_inv i_52912(.A(to_acu2[16]), .Z(n_43502));
	notech_inv i_52913(.A(n_3483), .Z(n_43503));
	notech_inv i_52914(.A(to_acu2[17]), .Z(n_43505));
	notech_inv i_52915(.A(to_acu2[18]), .Z(n_43506));
	notech_inv i_52916(.A(n_3482), .Z(n_43507));
	notech_inv i_52917(.A(to_acu2[19]), .Z(n_43508));
	notech_inv i_52918(.A(n_3481), .Z(n_43509));
	notech_inv i_52919(.A(to_acu2[20]), .Z(n_43511));
	notech_inv i_52920(.A(n_3480), .Z(n_43512));
	notech_inv i_52921(.A(to_acu2[21]), .Z(n_43513));
	notech_inv i_52922(.A(n_3479), .Z(n_43514));
	notech_inv i_52923(.A(to_acu2[22]), .Z(n_43515));
	notech_inv i_52924(.A(n_3478), .Z(n_43517));
	notech_inv i_52925(.A(to_acu2[23]), .Z(n_43518));
	notech_inv i_52926(.A(n_3477), .Z(n_43519));
	notech_inv i_52927(.A(to_acu2[24]), .Z(n_43520));
	notech_inv i_52928(.A(n_3476), .Z(n_43521));
	notech_inv i_52929(.A(to_acu2[25]), .Z(n_43523));
	notech_inv i_52930(.A(n_3475), .Z(n_43524));
	notech_inv i_52931(.A(to_acu2[26]), .Z(n_43525));
	notech_inv i_52932(.A(to_acu2[27]), .Z(n_43526));
	notech_inv i_52933(.A(to_acu2[28]), .Z(n_43527));
	notech_inv i_52934(.A(to_acu2[29]), .Z(n_43529));
	notech_inv i_52935(.A(n_3467), .Z(n_43530));
	notech_inv i_52936(.A(to_acu2[30]), .Z(n_43531));
	notech_inv i_52937(.A(to_acu2[31]), .Z(n_43532));
	notech_inv i_52938(.A(n_3466), .Z(n_43533));
	notech_inv i_52939(.A(to_acu2[32]), .Z(n_43535));
	notech_inv i_52940(.A(to_acu2[33]), .Z(n_43536));
	notech_inv i_52941(.A(to_acu2[34]), .Z(n_43537));
	notech_inv i_52942(.A(to_acu2[35]), .Z(n_43538));
	notech_inv i_52943(.A(to_acu2[36]), .Z(n_43539));
	notech_inv i_52944(.A(to_acu2[37]), .Z(n_43541));
	notech_inv i_52945(.A(to_acu2[38]), .Z(n_43542));
	notech_inv i_52946(.A(to_acu2[40]), .Z(n_43543));
	notech_inv i_52947(.A(to_acu2[41]), .Z(n_43544));
	notech_inv i_52948(.A(to_acu2[42]), .Z(n_43545));
	notech_inv i_52949(.A(to_acu2[43]), .Z(n_43547));
	notech_inv i_52950(.A(to_acu2[44]), .Z(n_43548));
	notech_inv i_52951(.A(to_acu2[45]), .Z(n_43549));
	notech_inv i_52952(.A(to_acu2[46]), .Z(n_43550));
	notech_inv i_52953(.A(to_acu2[47]), .Z(n_43551));
	notech_inv i_52954(.A(to_acu2[48]), .Z(n_43553));
	notech_inv i_52955(.A(to_acu2[49]), .Z(n_43554));
	notech_inv i_52956(.A(to_acu2[50]), .Z(n_43555));
	notech_inv i_52957(.A(to_acu2[51]), .Z(n_43556));
	notech_inv i_52958(.A(to_acu2[52]), .Z(n_43557));
	notech_inv i_52959(.A(to_acu2[53]), .Z(n_43559));
	notech_inv i_52960(.A(to_acu2[54]), .Z(n_43560));
	notech_inv i_52961(.A(to_acu2[55]), .Z(n_43561));
	notech_inv i_52962(.A(to_acu2[56]), .Z(n_43562));
	notech_inv i_52963(.A(to_acu2[57]), .Z(n_43563));
	notech_inv i_52964(.A(to_acu2[58]), .Z(n_43565));
	notech_inv i_52965(.A(to_acu2[59]), .Z(n_43566));
	notech_inv i_52966(.A(to_acu2[60]), .Z(n_43567));
	notech_inv i_52967(.A(to_acu2[61]), .Z(n_43568));
	notech_inv i_52968(.A(to_acu2[62]), .Z(n_43569));
	notech_inv i_52969(.A(to_acu2[63]), .Z(n_43571));
	notech_inv i_52970(.A(to_acu2[64]), .Z(n_43572));
	notech_inv i_52971(.A(to_acu2[65]), .Z(n_43573));
	notech_inv i_52972(.A(to_acu2[66]), .Z(n_43574));
	notech_inv i_52973(.A(to_acu2[67]), .Z(n_43575));
	notech_inv i_52974(.A(to_acu2[68]), .Z(n_43577));
	notech_inv i_52975(.A(to_acu2[69]), .Z(n_43578));
	notech_inv i_52976(.A(to_acu2[70]), .Z(n_43579));
	notech_inv i_52977(.A(to_acu2[71]), .Z(n_43580));
	notech_inv i_52978(.A(to_acu2[72]), .Z(n_43581));
	notech_inv i_52979(.A(to_acu2[73]), .Z(n_43583));
	notech_inv i_52980(.A(to_acu2[74]), .Z(n_43584));
	notech_inv i_52981(.A(to_acu2[75]), .Z(n_43585));
	notech_inv i_52982(.A(to_acu2[76]), .Z(n_43586));
	notech_inv i_52983(.A(to_acu2[77]), .Z(n_43587));
	notech_inv i_52984(.A(to_acu2[78]), .Z(n_43589));
	notech_inv i_52985(.A(to_acu2[79]), .Z(n_43590));
	notech_inv i_52986(.A(to_acu2[80]), .Z(n_43591));
	notech_inv i_52987(.A(to_acu2[81]), .Z(n_43592));
	notech_inv i_52988(.A(to_acu2[82]), .Z(n_43593));
	notech_inv i_52989(.A(to_acu2[83]), .Z(n_43595));
	notech_inv i_52990(.A(n_47596), .Z(n_43596));
	notech_inv i_52991(.A(to_acu2[84]), .Z(n_43597));
	notech_inv i_52992(.A(to_acu2[85]), .Z(n_43598));
	notech_inv i_52993(.A(to_acu2[86]), .Z(n_43599));
	notech_inv i_52994(.A(to_acu2[87]), .Z(n_43601));
	notech_inv i_52995(.A(to_acu2[88]), .Z(n_43602));
	notech_inv i_52996(.A(to_acu2[89]), .Z(n_43603));
	notech_inv i_52997(.A(to_acu2[90]), .Z(n_43604));
	notech_inv i_52998(.A(to_acu2[91]), .Z(n_43605));
	notech_inv i_52999(.A(to_acu2[92]), .Z(n_43607));
	notech_inv i_53000(.A(to_acu2[93]), .Z(n_43608));
	notech_inv i_53001(.A(to_acu2[94]), .Z(n_43609));
	notech_inv i_53002(.A(to_acu2[95]), .Z(n_43610));
	notech_inv i_53003(.A(to_acu2[96]), .Z(n_43611));
	notech_inv i_53004(.A(to_acu2[97]), .Z(n_43613));
	notech_inv i_53005(.A(to_acu2[98]), .Z(n_43614));
	notech_inv i_53006(.A(to_acu2[99]), .Z(n_43615));
	notech_inv i_53007(.A(to_acu2[100]), .Z(n_43616));
	notech_inv i_53008(.A(to_acu2[101]), .Z(n_43617));
	notech_inv i_53009(.A(to_acu2[102]), .Z(n_43619));
	notech_inv i_53010(.A(to_acu2[103]), .Z(n_43620));
	notech_inv i_53011(.A(to_acu2[104]), .Z(n_43621));
	notech_inv i_53012(.A(to_acu2[105]), .Z(n_43622));
	notech_inv i_53013(.A(to_acu2[106]), .Z(n_43623));
	notech_inv i_53014(.A(to_acu2[107]), .Z(n_43625));
	notech_inv i_53015(.A(to_acu2[108]), .Z(n_43626));
	notech_inv i_53016(.A(n_3379), .Z(n_43627));
	notech_inv i_53017(.A(to_acu2[109]), .Z(n_43628));
	notech_inv i_53018(.A(n_3378), .Z(n_43629));
	notech_inv i_53019(.A(to_acu2[110]), .Z(n_43631));
	notech_inv i_53020(.A(n_3377), .Z(n_43632));
	notech_inv i_53021(.A(to_acu2[111]), .Z(n_43633));
	notech_inv i_53022(.A(n_3376), .Z(n_43634));
	notech_inv i_53023(.A(to_acu2[112]), .Z(n_43635));
	notech_inv i_53024(.A(n_3375), .Z(n_43637));
	notech_inv i_53025(.A(to_acu2[113]), .Z(n_43638));
	notech_inv i_53026(.A(n_3374), .Z(n_43639));
	notech_inv i_53027(.A(to_acu2[114]), .Z(n_43640));
	notech_inv i_53028(.A(n_3373), .Z(n_43641));
	notech_inv i_53029(.A(to_acu2[115]), .Z(n_43643));
	notech_inv i_53030(.A(n_3372), .Z(n_43644));
	notech_inv i_53031(.A(to_acu2[116]), .Z(n_43645));
	notech_inv i_53032(.A(n_3371), .Z(n_43646));
	notech_inv i_53033(.A(to_acu2[117]), .Z(n_43647));
	notech_inv i_53034(.A(n_3370), .Z(n_43649));
	notech_inv i_53035(.A(to_acu2[118]), .Z(n_43650));
	notech_inv i_53036(.A(n_3369), .Z(n_43651));
	notech_inv i_53037(.A(to_acu2[119]), .Z(n_43652));
	notech_inv i_53038(.A(n_3368), .Z(n_43653));
	notech_inv i_53039(.A(to_acu2[120]), .Z(n_43655));
	notech_inv i_53040(.A(n_3367), .Z(n_43656));
	notech_inv i_53041(.A(to_acu2[121]), .Z(n_43657));
	notech_inv i_53042(.A(n_3366), .Z(n_43658));
	notech_inv i_53043(.A(to_acu2[122]), .Z(n_43659));
	notech_inv i_53044(.A(n_3365), .Z(n_43661));
	notech_inv i_53045(.A(to_acu2[123]), .Z(n_43662));
	notech_inv i_53046(.A(n_3364), .Z(n_43663));
	notech_inv i_53047(.A(to_acu2[124]), .Z(n_43664));
	notech_inv i_53048(.A(n_3363), .Z(n_43665));
	notech_inv i_53049(.A(to_acu2[125]), .Z(n_43667));
	notech_inv i_53050(.A(n_3362), .Z(n_43668));
	notech_inv i_53051(.A(to_acu2[126]), .Z(n_43669));
	notech_inv i_53052(.A(n_3361), .Z(n_43670));
	notech_inv i_53053(.A(to_acu2[127]), .Z(n_43671));
	notech_inv i_53054(.A(n_3360), .Z(n_43673));
	notech_inv i_53055(.A(to_acu2[128]), .Z(n_43674));
	notech_inv i_53056(.A(n_3359), .Z(n_43675));
	notech_inv i_53057(.A(to_acu2[129]), .Z(n_43676));
	notech_inv i_53058(.A(n_3358), .Z(n_43677));
	notech_inv i_53059(.A(to_acu2[130]), .Z(n_43679));
	notech_inv i_53060(.A(n_3357), .Z(n_43680));
	notech_inv i_53061(.A(to_acu2[131]), .Z(n_43681));
	notech_inv i_53062(.A(n_3356), .Z(n_43682));
	notech_inv i_53063(.A(to_acu2[132]), .Z(n_43683));
	notech_inv i_53064(.A(n_3355), .Z(n_43685));
	notech_inv i_53065(.A(to_acu2[133]), .Z(n_43686));
	notech_inv i_53066(.A(n_3354), .Z(n_43687));
	notech_inv i_53067(.A(to_acu2[134]), .Z(n_43688));
	notech_inv i_53068(.A(n_3353), .Z(n_43689));
	notech_inv i_53069(.A(to_acu2[135]), .Z(n_43691));
	notech_inv i_53070(.A(n_3352), .Z(n_43692));
	notech_inv i_53071(.A(to_acu2[136]), .Z(n_43693));
	notech_inv i_53072(.A(n_3351), .Z(n_43694));
	notech_inv i_53073(.A(to_acu2[137]), .Z(n_43695));
	notech_inv i_53074(.A(n_3350), .Z(n_43697));
	notech_inv i_53075(.A(to_acu2[138]), .Z(n_43698));
	notech_inv i_53076(.A(n_3349), .Z(n_43699));
	notech_inv i_53077(.A(to_acu2[139]), .Z(n_43700));
	notech_inv i_53078(.A(n_3348), .Z(n_43701));
	notech_inv i_53079(.A(to_acu2[140]), .Z(n_43703));
	notech_inv i_53080(.A(n_3347), .Z(n_43704));
	notech_inv i_53081(.A(to_acu2[141]), .Z(n_43705));
	notech_inv i_53082(.A(n_3346), .Z(n_43706));
	notech_inv i_53083(.A(to_acu2[142]), .Z(n_43707));
	notech_inv i_53084(.A(n_3345), .Z(n_43709));
	notech_inv i_53085(.A(to_acu2[143]), .Z(n_43710));
	notech_inv i_53086(.A(n_3344), .Z(n_43711));
	notech_inv i_53087(.A(to_acu2[144]), .Z(n_43712));
	notech_inv i_53088(.A(n_3343), .Z(n_43713));
	notech_inv i_53089(.A(to_acu2[145]), .Z(n_43715));
	notech_inv i_53090(.A(n_3342), .Z(n_43716));
	notech_inv i_53091(.A(to_acu2[146]), .Z(n_43717));
	notech_inv i_53092(.A(n_3341), .Z(n_43718));
	notech_inv i_53093(.A(to_acu2[147]), .Z(n_43719));
	notech_inv i_53094(.A(n_3340), .Z(n_43721));
	notech_inv i_53095(.A(to_acu2[148]), .Z(n_43722));
	notech_inv i_53096(.A(n_3339), .Z(n_43723));
	notech_inv i_53097(.A(to_acu2[149]), .Z(n_43724));
	notech_inv i_53098(.A(n_3338), .Z(n_43725));
	notech_inv i_53099(.A(to_acu2[150]), .Z(n_43727));
	notech_inv i_53100(.A(n_3336), .Z(n_43728));
	notech_inv i_53101(.A(to_acu2[151]), .Z(n_43729));
	notech_inv i_53102(.A(n_3334), .Z(n_43730));
	notech_inv i_53103(.A(to_acu2[152]), .Z(n_43731));
	notech_inv i_53104(.A(n_3332), .Z(n_43733));
	notech_inv i_53105(.A(to_acu2[153]), .Z(n_43734));
	notech_inv i_53106(.A(n_3330), .Z(n_43735));
	notech_inv i_53107(.A(to_acu2[154]), .Z(n_43736));
	notech_inv i_53108(.A(n_3328), .Z(n_43737));
	notech_inv i_53109(.A(to_acu2[155]), .Z(n_43739));
	notech_inv i_53110(.A(n_3326), .Z(n_43740));
	notech_inv i_53111(.A(to_acu2[156]), .Z(n_43741));
	notech_inv i_53112(.A(n_3324), .Z(n_43742));
	notech_inv i_53113(.A(to_acu2[157]), .Z(n_43743));
	notech_inv i_53114(.A(n_3322), .Z(n_43745));
	notech_inv i_53115(.A(to_acu2[158]), .Z(n_43746));
	notech_inv i_53116(.A(n_3320), .Z(n_43747));
	notech_inv i_53117(.A(to_acu2[159]), .Z(n_43748));
	notech_inv i_53118(.A(n_3318), .Z(n_43749));
	notech_inv i_53119(.A(to_acu2[160]), .Z(n_43751));
	notech_inv i_53120(.A(n_3316), .Z(n_43752));
	notech_inv i_53121(.A(to_acu2[161]), .Z(n_43753));
	notech_inv i_53122(.A(n_3315), .Z(n_43754));
	notech_inv i_53123(.A(to_acu2[162]), .Z(n_43755));
	notech_inv i_53124(.A(n_3314), .Z(n_43757));
	notech_inv i_53125(.A(to_acu2[163]), .Z(n_43758));
	notech_inv i_53126(.A(n_3312), .Z(n_43759));
	notech_inv i_53127(.A(to_acu2[164]), .Z(n_43760));
	notech_inv i_53128(.A(n_3310), .Z(n_43761));
	notech_inv i_53129(.A(to_acu2[165]), .Z(n_43763));
	notech_inv i_53130(.A(n_3308), .Z(n_43764));
	notech_inv i_53131(.A(to_acu2[166]), .Z(n_43765));
	notech_inv i_53132(.A(n_3306), .Z(n_43766));
	notech_inv i_53133(.A(to_acu2[167]), .Z(n_43767));
	notech_inv i_53134(.A(n_3304), .Z(n_43769));
	notech_inv i_53135(.A(to_acu2[168]), .Z(n_43770));
	notech_inv i_53136(.A(to_acu2[169]), .Z(n_43771));
	notech_inv i_53137(.A(to_acu2[170]), .Z(n_43772));
	notech_inv i_53138(.A(to_acu2[171]), .Z(n_43773));
	notech_inv i_53139(.A(to_acu2[172]), .Z(n_43775));
	notech_inv i_53140(.A(to_acu2[173]), .Z(n_43776));
	notech_inv i_53141(.A(to_acu2[174]), .Z(n_43777));
	notech_inv i_53142(.A(to_acu2[175]), .Z(n_43778));
	notech_inv i_53143(.A(to_acu2[176]), .Z(n_43779));
	notech_inv i_53144(.A(to_acu2[177]), .Z(n_43781));
	notech_inv i_53145(.A(to_acu2[178]), .Z(n_43782));
	notech_inv i_53146(.A(to_acu2[179]), .Z(n_43783));
	notech_inv i_53147(.A(to_acu2[180]), .Z(n_43784));
	notech_inv i_53148(.A(to_acu2[181]), .Z(n_43785));
	notech_inv i_53149(.A(n_1608), .Z(n_43787));
	notech_inv i_53150(.A(to_acu2[182]), .Z(n_43788));
	notech_inv i_53151(.A(to_acu2[183]), .Z(n_43789));
	notech_inv i_53152(.A(to_acu2[184]), .Z(n_43790));
	notech_inv i_53153(.A(to_acu2[185]), .Z(n_43791));
	notech_inv i_53154(.A(to_acu2[186]), .Z(n_43793));
	notech_inv i_53155(.A(to_acu2[187]), .Z(n_43794));
	notech_inv i_53156(.A(to_acu2[188]), .Z(n_43795));
	notech_inv i_53157(.A(to_acu2[189]), .Z(n_43796));
	notech_inv i_53158(.A(n_2846), .Z(n_43797));
	notech_inv i_53159(.A(to_acu2[190]), .Z(n_43799));
	notech_inv i_53160(.A(to_acu2[191]), .Z(n_43800));
	notech_inv i_53161(.A(to_acu2[192]), .Z(n_43801));
	notech_inv i_53162(.A(to_acu2[193]), .Z(n_43802));
	notech_inv i_53163(.A(to_acu2[194]), .Z(n_43803));
	notech_inv i_53164(.A(to_acu2[195]), .Z(n_43805));
	notech_inv i_53165(.A(to_acu2[196]), .Z(n_43806));
	notech_inv i_53166(.A(to_acu2[197]), .Z(n_43807));
	notech_inv i_53167(.A(to_acu2[198]), .Z(n_43808));
	notech_inv i_53168(.A(to_acu2[199]), .Z(n_43809));
	notech_inv i_53169(.A(to_acu2[200]), .Z(n_43811));
	notech_inv i_53170(.A(to_acu2[201]), .Z(n_43812));
	notech_inv i_53171(.A(to_acu2[202]), .Z(n_43813));
	notech_inv i_53172(.A(n_3270), .Z(n_43814));
	notech_inv i_53173(.A(to_acu2[203]), .Z(n_43815));
	notech_inv i_53174(.A(to_acu2[204]), .Z(n_43817));
	notech_inv i_53175(.A(to_acu2[205]), .Z(n_43818));
	notech_inv i_53176(.A(to_acu2[206]), .Z(n_43819));
	notech_inv i_53177(.A(n_3272), .Z(n_43820));
	notech_inv i_53178(.A(to_acu2[207]), .Z(n_43821));
	notech_inv i_53179(.A(to_acu2[208]), .Z(n_43823));
	notech_inv i_53180(.A(to_acu2[209]), .Z(n_43824));
	notech_inv i_53181(.A(to_acu2[210]), .Z(n_43825));
	notech_inv i_53182(.A(to_acu1[0]), .Z(n_43826));
	notech_inv i_53183(.A(n_3266), .Z(n_43827));
	notech_inv i_53184(.A(to_acu1[1]), .Z(n_43829));
	notech_inv i_53185(.A(to_acu1[2]), .Z(n_43830));
	notech_inv i_53186(.A(to_acu1[3]), .Z(n_43831));
	notech_inv i_53187(.A(n_3260), .Z(n_43832));
	notech_inv i_53188(.A(to_acu1[4]), .Z(n_43833));
	notech_inv i_53189(.A(to_acu1[5]), .Z(n_43835));
	notech_inv i_53190(.A(to_acu1[6]), .Z(n_43836));
	notech_inv i_53191(.A(to_acu1[7]), .Z(n_43837));
	notech_inv i_53192(.A(n_3254), .Z(n_43838));
	notech_inv i_53193(.A(to_acu1[8]), .Z(n_43839));
	notech_inv i_53194(.A(n_3253), .Z(n_43841));
	notech_inv i_53195(.A(to_acu1[9]), .Z(n_43842));
	notech_inv i_53196(.A(n_48498), .Z(n_43843));
	notech_inv i_53197(.A(to_acu1[10]), .Z(n_43844));
	notech_inv i_53198(.A(n_3252), .Z(n_43845));
	notech_inv i_53199(.A(to_acu1[11]), .Z(n_43847));
	notech_inv i_53200(.A(to_acu1[12]), .Z(n_43848));
	notech_inv i_53201(.A(n_3251), .Z(n_43849));
	notech_inv i_53202(.A(to_acu1[13]), .Z(n_43850));
	notech_inv i_53203(.A(n_3250), .Z(n_43851));
	notech_inv i_53204(.A(to_acu1[14]), .Z(n_43853));
	notech_inv i_53205(.A(to_acu1[15]), .Z(n_43854));
	notech_inv i_53206(.A(n_3249), .Z(n_43855));
	notech_inv i_53207(.A(to_acu1[16]), .Z(n_43856));
	notech_inv i_53208(.A(n_3248), .Z(n_43857));
	notech_inv i_53209(.A(to_acu1[17]), .Z(n_43859));
	notech_inv i_53210(.A(to_acu1[18]), .Z(n_43860));
	notech_inv i_53211(.A(n_3247), .Z(n_43861));
	notech_inv i_53212(.A(n_48552), .Z(n_43862));
	notech_inv i_53213(.A(to_acu1[19]), .Z(n_43863));
	notech_inv i_53214(.A(n_48558), .Z(n_43865));
	notech_inv i_53215(.A(to_acu1[20]), .Z(n_43866));
	notech_inv i_53216(.A(n_48564), .Z(n_43867));
	notech_inv i_53217(.A(to_acu1[21]), .Z(n_43868));
	notech_inv i_53218(.A(n_48570), .Z(n_43869));
	notech_inv i_53219(.A(to_acu1[22]), .Z(n_43871));
	notech_inv i_53220(.A(n_48576), .Z(n_43872));
	notech_inv i_53221(.A(to_acu1[23]), .Z(n_43873));
	notech_inv i_53222(.A(n_48582), .Z(n_43874));
	notech_inv i_53223(.A(to_acu1[24]), .Z(n_43875));
	notech_inv i_53224(.A(n_48588), .Z(n_43877));
	notech_inv i_53225(.A(to_acu1[25]), .Z(n_43878));
	notech_inv i_53226(.A(n_3243), .Z(n_43879));
	notech_inv i_53227(.A(n_48594), .Z(n_43880));
	notech_inv i_53228(.A(to_acu1[26]), .Z(n_43881));
	notech_inv i_53229(.A(n_48600), .Z(n_43883));
	notech_inv i_53230(.A(to_acu1[27]), .Z(n_43884));
	notech_inv i_53231(.A(n_48606), .Z(n_43885));
	notech_inv i_53232(.A(to_acu1[28]), .Z(n_43886));
	notech_inv i_53233(.A(n_3242), .Z(n_43887));
	notech_inv i_53234(.A(n_48612), .Z(n_43889));
	notech_inv i_53235(.A(to_acu1[29]), .Z(n_43890));
	notech_inv i_53236(.A(n_48618), .Z(n_43891));
	notech_inv i_53237(.A(to_acu1[30]), .Z(n_43892));
	notech_inv i_53238(.A(n_3241), .Z(n_43893));
	notech_inv i_53239(.A(to_acu1[31]), .Z(n_43895));
	notech_inv i_53240(.A(to_acu1[32]), .Z(n_43896));
	notech_inv i_53241(.A(n_3240), .Z(n_43897));
	notech_inv i_53242(.A(to_acu1[33]), .Z(n_43898));
	notech_inv i_53243(.A(n_3239), .Z(n_43899));
	notech_inv i_53244(.A(to_acu1[34]), .Z(n_43901));
	notech_inv i_53245(.A(to_acu1[35]), .Z(n_43902));
	notech_inv i_53246(.A(n_3238), .Z(n_43903));
	notech_inv i_53247(.A(to_acu1[36]), .Z(n_43904));
	notech_inv i_53248(.A(n_3237), .Z(n_43905));
	notech_inv i_53249(.A(to_acu1[37]), .Z(n_43907));
	notech_inv i_53250(.A(to_acu1[38]), .Z(n_43908));
	notech_inv i_53251(.A(to_acu1[40]), .Z(n_43909));
	notech_inv i_53252(.A(n_2590), .Z(n_43910));
	notech_inv i_53253(.A(n_48684), .Z(n_43911));
	notech_inv i_53254(.A(to_acu1[41]), .Z(n_43913));
	notech_inv i_53255(.A(to_acu1[42]), .Z(n_43914));
	notech_inv i_53256(.A(to_acu1[43]), .Z(n_43915));
	notech_inv i_53257(.A(to_acu1[44]), .Z(n_43916));
	notech_inv i_53258(.A(n_48708), .Z(n_43917));
	notech_inv i_53259(.A(to_acu1[45]), .Z(n_43919));
	notech_inv i_53260(.A(to_acu1[46]), .Z(n_43920));
	notech_inv i_53261(.A(to_acu1[47]), .Z(n_43921));
	notech_inv i_53262(.A(to_acu1[48]), .Z(n_43922));
	notech_inv i_53263(.A(to_acu1[49]), .Z(n_43923));
	notech_inv i_53264(.A(to_acu1[50]), .Z(n_43925));
	notech_inv i_53265(.A(to_acu1[51]), .Z(n_43926));
	notech_inv i_53266(.A(to_acu1[52]), .Z(n_43927));
	notech_inv i_53267(.A(to_acu1[53]), .Z(n_43928));
	notech_inv i_53268(.A(to_acu1[54]), .Z(n_43929));
	notech_inv i_53269(.A(to_acu1[55]), .Z(n_43931));
	notech_inv i_53270(.A(to_acu1[56]), .Z(n_43932));
	notech_inv i_53271(.A(to_acu1[57]), .Z(n_43933));
	notech_inv i_53272(.A(to_acu1[58]), .Z(n_43934));
	notech_inv i_53273(.A(to_acu1[59]), .Z(n_43935));
	notech_inv i_53274(.A(to_acu1[60]), .Z(n_43937));
	notech_inv i_53275(.A(to_acu1[61]), .Z(n_43938));
	notech_inv i_53276(.A(to_acu1[62]), .Z(n_43939));
	notech_inv i_53277(.A(to_acu1[63]), .Z(n_43940));
	notech_inv i_53278(.A(to_acu1[64]), .Z(n_43941));
	notech_inv i_53279(.A(to_acu1[65]), .Z(n_43943));
	notech_inv i_53280(.A(to_acu1[66]), .Z(n_43944));
	notech_inv i_53281(.A(to_acu1[67]), .Z(n_43945));
	notech_inv i_53282(.A(to_acu1[68]), .Z(n_43946));
	notech_inv i_53283(.A(to_acu1[69]), .Z(n_43947));
	notech_inv i_53284(.A(to_acu1[70]), .Z(n_43949));
	notech_inv i_53285(.A(to_acu1[71]), .Z(n_43950));
	notech_inv i_53286(.A(to_acu1[72]), .Z(n_43951));
	notech_inv i_53287(.A(to_acu1[73]), .Z(n_43952));
	notech_inv i_53288(.A(to_acu1[74]), .Z(n_43953));
	notech_inv i_53289(.A(to_acu1[75]), .Z(n_43955));
	notech_inv i_53290(.A(to_acu1[76]), .Z(n_43956));
	notech_inv i_53291(.A(to_acu1[77]), .Z(n_43957));
	notech_inv i_53292(.A(to_acu1[78]), .Z(n_43958));
	notech_inv i_53293(.A(to_acu1[79]), .Z(n_43959));
	notech_inv i_53294(.A(to_acu1[80]), .Z(n_43961));
	notech_inv i_53295(.A(to_acu1[81]), .Z(n_43962));
	notech_inv i_53296(.A(to_acu1[82]), .Z(n_43963));
	notech_inv i_53297(.A(to_acu1[83]), .Z(n_43964));
	notech_inv i_53298(.A(to_acu1[84]), .Z(n_43965));
	notech_inv i_53299(.A(to_acu1[85]), .Z(n_43967));
	notech_inv i_53300(.A(to_acu1[86]), .Z(n_43968));
	notech_inv i_53301(.A(to_acu1[87]), .Z(n_43969));
	notech_inv i_53302(.A(to_acu1[88]), .Z(n_43970));
	notech_inv i_53303(.A(to_acu1[89]), .Z(n_43971));
	notech_inv i_53304(.A(to_acu1[90]), .Z(n_43973));
	notech_inv i_53305(.A(to_acu1[91]), .Z(n_43974));
	notech_inv i_53306(.A(to_acu1[92]), .Z(n_43975));
	notech_inv i_53307(.A(to_acu1[93]), .Z(n_43976));
	notech_inv i_53308(.A(to_acu1[94]), .Z(n_43977));
	notech_inv i_53309(.A(to_acu1[95]), .Z(n_43979));
	notech_inv i_53310(.A(to_acu1[96]), .Z(n_43980));
	notech_inv i_53311(.A(to_acu1[97]), .Z(n_43981));
	notech_inv i_53312(.A(to_acu1[98]), .Z(n_43982));
	notech_inv i_53313(.A(n_49032), .Z(n_43983));
	notech_inv i_53314(.A(to_acu1[99]), .Z(n_43985));
	notech_inv i_53315(.A(n_49038), .Z(n_43986));
	notech_inv i_53316(.A(to_acu1[100]), .Z(n_43987));
	notech_inv i_53317(.A(to_acu1[101]), .Z(n_43988));
	notech_inv i_53318(.A(n_49050), .Z(n_43989));
	notech_inv i_53319(.A(to_acu1[102]), .Z(n_43991));
	notech_inv i_53320(.A(n_49056), .Z(n_43992));
	notech_inv i_53321(.A(to_acu1[103]), .Z(n_43993));
	notech_inv i_53322(.A(to_acu1[104]), .Z(n_43994));
	notech_inv i_53323(.A(n_49068), .Z(n_43995));
	notech_inv i_53324(.A(to_acu1[105]), .Z(n_43997));
	notech_inv i_53325(.A(to_acu1[106]), .Z(n_43998));
	notech_inv i_53326(.A(n_49080), .Z(n_43999));
	notech_inv i_53327(.A(to_acu1[107]), .Z(n_44000));
	notech_inv i_53328(.A(n_49086), .Z(n_44001));
	notech_inv i_53329(.A(to_acu1[108]), .Z(n_44003));
	notech_inv i_53330(.A(n_49092), .Z(n_44004));
	notech_inv i_53331(.A(to_acu1[109]), .Z(n_44005));
	notech_inv i_53332(.A(n_49098), .Z(n_44006));
	notech_inv i_53333(.A(to_acu1[110]), .Z(n_44007));
	notech_inv i_53334(.A(n_49104), .Z(n_44009));
	notech_inv i_53335(.A(to_acu1[111]), .Z(n_44010));
	notech_inv i_53336(.A(n_49110), .Z(n_44011));
	notech_inv i_53337(.A(to_acu1[112]), .Z(n_44012));
	notech_inv i_53338(.A(to_acu1[113]), .Z(n_44013));
	notech_inv i_53339(.A(n_49122), .Z(n_44015));
	notech_inv i_53340(.A(to_acu1[114]), .Z(n_44016));
	notech_inv i_53341(.A(n_49128), .Z(n_44017));
	notech_inv i_53342(.A(to_acu1[115]), .Z(n_44018));
	notech_inv i_53343(.A(n_49134), .Z(n_44019));
	notech_inv i_53344(.A(to_acu1[116]), .Z(n_44021));
	notech_inv i_53345(.A(n_49140), .Z(n_44022));
	notech_inv i_53346(.A(to_acu1[117]), .Z(n_44023));
	notech_inv i_53347(.A(n_49146), .Z(n_44024));
	notech_inv i_53348(.A(to_acu1[118]), .Z(n_44025));
	notech_inv i_53349(.A(n_49152), .Z(n_44027));
	notech_inv i_53350(.A(to_acu1[119]), .Z(n_44028));
	notech_inv i_53351(.A(n_49158), .Z(n_44029));
	notech_inv i_53352(.A(to_acu1[120]), .Z(n_44030));
	notech_inv i_53353(.A(n_49164), .Z(n_44031));
	notech_inv i_53354(.A(to_acu1[121]), .Z(n_44033));
	notech_inv i_53355(.A(n_49170), .Z(n_44034));
	notech_inv i_53356(.A(to_acu1[122]), .Z(n_44035));
	notech_inv i_53357(.A(to_acu1[123]), .Z(n_44036));
	notech_inv i_53358(.A(n_49182), .Z(n_44037));
	notech_inv i_53359(.A(to_acu1[124]), .Z(n_44038));
	notech_inv i_53360(.A(to_acu1[125]), .Z(n_44039));
	notech_inv i_53361(.A(to_acu1[126]), .Z(n_44040));
	notech_inv i_53362(.A(to_acu1[127]), .Z(n_44042));
	notech_inv i_53363(.A(to_acu1[128]), .Z(n_44043));
	notech_inv i_53364(.A(to_acu1[129]), .Z(n_44045));
	notech_inv i_53365(.A(to_acu1[130]), .Z(n_44046));
	notech_inv i_53366(.A(to_acu1[131]), .Z(n_44047));
	notech_inv i_53367(.A(to_acu1[132]), .Z(n_44048));
	notech_inv i_53368(.A(to_acu1[133]), .Z(n_44049));
	notech_inv i_53369(.A(to_acu1[134]), .Z(n_44050));
	notech_inv i_53370(.A(to_acu1[135]), .Z(n_44051));
	notech_inv i_53371(.A(to_acu1[136]), .Z(n_44052));
	notech_inv i_53372(.A(to_acu1[137]), .Z(n_44053));
	notech_inv i_53373(.A(to_acu1[138]), .Z(n_44054));
	notech_inv i_53374(.A(to_acu1[139]), .Z(n_44055));
	notech_inv i_53375(.A(to_acu1[140]), .Z(n_44056));
	notech_inv i_53376(.A(to_acu1[141]), .Z(n_44057));
	notech_inv i_53377(.A(to_acu1[142]), .Z(n_44059));
	notech_inv i_53378(.A(to_acu1[143]), .Z(n_44060));
	notech_inv i_53379(.A(to_acu1[144]), .Z(n_44061));
	notech_inv i_53380(.A(to_acu1[145]), .Z(n_44062));
	notech_inv i_53381(.A(to_acu1[146]), .Z(n_44063));
	notech_inv i_53382(.A(to_acu1[147]), .Z(n_44065));
	notech_inv i_53383(.A(to_acu1[148]), .Z(n_44066));
	notech_inv i_53384(.A(to_acu1[149]), .Z(n_44067));
	notech_inv i_53385(.A(to_acu1[150]), .Z(n_44068));
	notech_inv i_53386(.A(to_acu1[151]), .Z(n_44069));
	notech_inv i_53387(.A(to_acu1[152]), .Z(n_44071));
	notech_inv i_53388(.A(to_acu1[153]), .Z(n_44072));
	notech_inv i_53389(.A(to_acu1[154]), .Z(n_44073));
	notech_inv i_53390(.A(to_acu1[155]), .Z(n_44074));
	notech_inv i_53391(.A(to_acu1[156]), .Z(n_44075));
	notech_inv i_53392(.A(to_acu1[157]), .Z(n_44077));
	notech_inv i_53393(.A(to_acu1[158]), .Z(n_44078));
	notech_inv i_53394(.A(to_acu1[159]), .Z(n_44079));
	notech_inv i_53395(.A(to_acu1[160]), .Z(n_44080));
	notech_inv i_53396(.A(to_acu1[161]), .Z(n_44081));
	notech_inv i_53397(.A(to_acu1[162]), .Z(n_44083));
	notech_inv i_53398(.A(to_acu1[163]), .Z(n_44084));
	notech_inv i_53399(.A(to_acu1[164]), .Z(n_44085));
	notech_inv i_53400(.A(to_acu1[165]), .Z(n_44086));
	notech_inv i_53401(.A(to_acu1[166]), .Z(n_44087));
	notech_inv i_53402(.A(to_acu1[167]), .Z(n_44089));
	notech_inv i_53403(.A(to_acu1[168]), .Z(n_44090));
	notech_inv i_53404(.A(to_acu1[169]), .Z(n_44091));
	notech_inv i_53405(.A(to_acu1[170]), .Z(n_44092));
	notech_inv i_53406(.A(to_acu1[171]), .Z(n_44093));
	notech_inv i_53407(.A(to_acu1[172]), .Z(n_44095));
	notech_inv i_53408(.A(to_acu1[173]), .Z(n_44096));
	notech_inv i_53409(.A(to_acu1[174]), .Z(n_44097));
	notech_inv i_53410(.A(to_acu1[175]), .Z(n_44098));
	notech_inv i_53411(.A(to_acu1[176]), .Z(n_44099));
	notech_inv i_53412(.A(to_acu1[177]), .Z(n_44101));
	notech_inv i_53413(.A(to_acu1[178]), .Z(n_44102));
	notech_inv i_53414(.A(to_acu1[179]), .Z(n_44103));
	notech_inv i_53415(.A(to_acu1[180]), .Z(n_44104));
	notech_inv i_53416(.A(n_3117), .Z(n_44105));
	notech_inv i_53417(.A(to_acu1[181]), .Z(n_44107));
	notech_inv i_53418(.A(to_acu1[182]), .Z(n_44108));
	notech_inv i_53419(.A(to_acu1[183]), .Z(n_44109));
	notech_inv i_53420(.A(to_acu1[184]), .Z(n_44110));
	notech_inv i_53421(.A(to_acu1[185]), .Z(n_44111));
	notech_inv i_53422(.A(to_acu1[186]), .Z(n_44113));
	notech_inv i_53423(.A(to_acu1[187]), .Z(n_44114));
	notech_inv i_53424(.A(to_acu1[188]), .Z(n_44115));
	notech_inv i_53425(.A(to_acu1[189]), .Z(n_44116));
	notech_inv i_53426(.A(n_49578), .Z(n_44117));
	notech_inv i_53427(.A(to_acu1[190]), .Z(n_44119));
	notech_inv i_53428(.A(n_49584), .Z(n_44120));
	notech_inv i_53429(.A(to_acu1[191]), .Z(n_44121));
	notech_inv i_53430(.A(n_49590), .Z(n_44122));
	notech_inv i_53431(.A(to_acu1[192]), .Z(n_44123));
	notech_inv i_53432(.A(to_acu1[193]), .Z(n_44125));
	notech_inv i_53433(.A(to_acu1[194]), .Z(n_44126));
	notech_inv i_53434(.A(to_acu1[195]), .Z(n_44127));
	notech_inv i_53435(.A(to_acu1[196]), .Z(n_44128));
	notech_inv i_53436(.A(to_acu1[197]), .Z(n_44129));
	notech_inv i_53437(.A(to_acu1[198]), .Z(n_44131));
	notech_inv i_53438(.A(to_acu1[199]), .Z(n_44132));
	notech_inv i_53439(.A(to_acu1[200]), .Z(n_44133));
	notech_inv i_53440(.A(to_acu1[201]), .Z(n_44134));
	notech_inv i_53441(.A(to_acu1[202]), .Z(n_44135));
	notech_inv i_53442(.A(to_acu1[203]), .Z(n_44137));
	notech_inv i_53443(.A(to_acu1[204]), .Z(n_44138));
	notech_inv i_53444(.A(to_acu1[205]), .Z(n_44139));
	notech_inv i_53445(.A(to_acu1[206]), .Z(n_44140));
	notech_inv i_53446(.A(n_49680), .Z(n_44141));
	notech_inv i_53447(.A(to_acu1[207]), .Z(n_44143));
	notech_inv i_53448(.A(to_acu1[208]), .Z(n_44144));
	notech_inv i_53449(.A(n_49692), .Z(n_44145));
	notech_inv i_53450(.A(to_acu1[209]), .Z(n_44146));
	notech_inv i_53451(.A(to_acu1[210]), .Z(n_44147));
	notech_inv i_53452(.A(n_41736), .Z(n_44149));
	notech_inv i_53453(.A(lenpc2[0]), .Z(n_44150));
	notech_inv i_53454(.A(lenpc2[1]), .Z(n_44151));
	notech_inv i_53455(.A(lenpc2[2]), .Z(n_44152));
	notech_inv i_53456(.A(lenpc2[3]), .Z(n_44153));
	notech_inv i_53457(.A(lenpc2[4]), .Z(n_44155));
	notech_inv i_53458(.A(lenpc2[5]), .Z(n_44156));
	notech_inv i_53459(.A(n_3079), .Z(n_44157));
	notech_inv i_53460(.A(n_3077), .Z(n_44158));
	notech_inv i_53461(.A(n_3072), .Z(n_44159));
	notech_inv i_53462(.A(n_2423), .Z(n_44161));
	notech_inv i_53463(.A(n_3064), .Z(n_44162));
	notech_inv i_53464(.A(n_3058), .Z(n_44163));
	notech_inv i_53465(.A(n_2942), .Z(n_44164));
	notech_inv i_53466(.A(n_3009), .Z(n_44165));
	notech_inv i_53467(.A(n_3012), .Z(n_44167));
	notech_inv i_53468(.A(n_2998), .Z(n_44168));
	notech_inv i_53469(.A(n_2996), .Z(n_44169));
	notech_inv i_53470(.A(n_2995), .Z(n_44170));
	notech_inv i_53471(.A(lenpc1[0]), .Z(n_44171));
	notech_inv i_53472(.A(n_44064), .Z(n_44173));
	notech_inv i_53473(.A(lenpc1[1]), .Z(n_44174));
	notech_inv i_53474(.A(n_44070), .Z(n_44175));
	notech_inv i_53475(.A(lenpc1[2]), .Z(n_44176));
	notech_inv i_53476(.A(n_44076), .Z(n_44177));
	notech_inv i_53477(.A(lenpc1[3]), .Z(n_44179));
	notech_inv i_53478(.A(n_44082), .Z(n_44180));
	notech_inv i_53479(.A(lenpc1[4]), .Z(n_44181));
	notech_inv i_53480(.A(n_44088), .Z(n_44182));
	notech_inv i_53481(.A(lenpc1[5]), .Z(n_44183));
	notech_inv i_53482(.A(n_2985), .Z(n_44185));
	notech_inv i_53483(.A(n_2983), .Z(n_44186));
	notech_inv i_53484(.A(n_2979), .Z(n_44187));
	notech_inv i_53485(.A(n_2978), .Z(n_44188));
	notech_inv i_53486(.A(n_46130), .Z(n_44189));
	notech_inv i_53487(.A(n_46136), .Z(n_44191));
	notech_inv i_53488(.A(n_46142), .Z(n_44192));
	notech_inv i_53489(.A(n_46148), .Z(n_44193));
	notech_inv i_53490(.A(n_46154), .Z(n_44194));
	notech_inv i_53491(.A(n_46160), .Z(n_44195));
	notech_inv i_53492(.A(opz1[0]), .Z(n_44197));
	notech_inv i_53493(.A(opz1[1]), .Z(n_44198));
	notech_inv i_53494(.A(n_2849), .Z(n_44199));
	notech_inv i_53495(.A(n_2379), .Z(n_44200));
	notech_inv i_53496(.A(n_42814), .Z(n_44201));
	notech_inv i_53497(.A(n_42820), .Z(n_44203));
	notech_inv i_53498(.A(n_42826), .Z(n_44204));
	notech_inv i_53499(.A(n_42832), .Z(n_44205));
	notech_inv i_53500(.A(n_42838), .Z(n_44206));
	notech_inv i_53501(.A(n_42844), .Z(n_44207));
	notech_inv i_53502(.A(n_42850), .Z(n_44209));
	notech_inv i_53503(.A(n_42856), .Z(n_44210));
	notech_inv i_53504(.A(n_42862), .Z(n_44211));
	notech_inv i_53505(.A(n_42868), .Z(n_44212));
	notech_inv i_53506(.A(n_42874), .Z(n_44213));
	notech_inv i_53507(.A(n_42880), .Z(n_44215));
	notech_inv i_53508(.A(n_42892), .Z(n_44216));
	notech_inv i_53509(.A(n_42946), .Z(n_44217));
	notech_inv i_53510(.A(n_42952), .Z(n_44218));
	notech_inv i_53511(.A(n_42958), .Z(n_44219));
	notech_inv i_53512(.A(n_42964), .Z(n_44221));
	notech_inv i_53513(.A(n_42982), .Z(n_44222));
	notech_inv i_53514(.A(n_42988), .Z(n_44223));
	notech_inv i_53515(.A(n_42994), .Z(n_44224));
	notech_inv i_53516(.A(n_43000), .Z(n_44225));
	notech_inv i_53517(.A(n_43024), .Z(n_44227));
	notech_inv i_53518(.A(n_43030), .Z(n_44228));
	notech_inv i_53519(.A(n_43036), .Z(n_44229));
	notech_inv i_53520(.A(n_43042), .Z(n_44230));
	notech_inv i_53521(.A(n_43048), .Z(n_44231));
	notech_inv i_53522(.A(n_43054), .Z(n_44233));
	notech_inv i_53523(.A(n_43060), .Z(n_44234));
	notech_inv i_53524(.A(n_43090), .Z(n_44235));
	notech_inv i_53525(.A(n_43120), .Z(n_44236));
	notech_inv i_53526(.A(n_43126), .Z(n_44237));
	notech_inv i_53527(.A(n_43144), .Z(n_44239));
	notech_inv i_53528(.A(n_43156), .Z(n_44240));
	notech_inv i_53529(.A(n_43162), .Z(n_44241));
	notech_inv i_53530(.A(n_43174), .Z(n_44242));
	notech_inv i_53531(.A(n_43180), .Z(n_44243));
	notech_inv i_53532(.A(n_43186), .Z(n_44245));
	notech_inv i_53533(.A(n_43192), .Z(n_44246));
	notech_inv i_53534(.A(n_43198), .Z(n_44247));
	notech_inv i_53535(.A(n_43204), .Z(n_44248));
	notech_inv i_53536(.A(n_43210), .Z(n_44249));
	notech_inv i_53537(.A(n_43216), .Z(n_44250));
	notech_inv i_53538(.A(n_43222), .Z(n_44251));
	notech_inv i_53539(.A(n_43228), .Z(n_44252));
	notech_inv i_53540(.A(n_43234), .Z(n_44253));
	notech_inv i_53541(.A(n_43240), .Z(n_44254));
	notech_inv i_53542(.A(n_43246), .Z(n_44255));
	notech_inv i_53543(.A(n_43252), .Z(n_44256));
	notech_inv i_53544(.A(n_43258), .Z(n_44257));
	notech_inv i_53545(.A(n_43264), .Z(n_44258));
	notech_inv i_53546(.A(n_43270), .Z(n_44259));
	notech_inv i_53547(.A(n_43282), .Z(n_44260));
	notech_inv i_53548(.A(n_43288), .Z(n_44261));
	notech_inv i_53549(.A(n_43294), .Z(n_44262));
	notech_inv i_53550(.A(n_43300), .Z(n_44263));
	notech_inv i_53551(.A(n_43306), .Z(n_44264));
	notech_inv i_53552(.A(n_43312), .Z(n_44265));
	notech_inv i_53553(.A(n_43318), .Z(n_44266));
	notech_inv i_53554(.A(n_43354), .Z(n_44267));
	notech_inv i_53555(.A(n_43360), .Z(n_44268));
	notech_inv i_53556(.A(n_43366), .Z(n_44269));
	notech_inv i_53557(.A(n_43408), .Z(n_44270));
	notech_inv i_53558(.A(n_43420), .Z(n_44271));
	notech_inv i_53559(.A(n_43432), .Z(n_44272));
	notech_inv i_53560(.A(n_43516), .Z(n_44273));
	notech_inv i_53561(.A(n_43522), .Z(n_44274));
	notech_inv i_53562(.A(n_43528), .Z(n_44275));
	notech_inv i_53563(.A(n_43534), .Z(n_44276));
	notech_inv i_53564(.A(n_43540), .Z(n_44277));
	notech_inv i_53565(.A(n_43546), .Z(n_44279));
	notech_inv i_53566(.A(n_43552), .Z(n_44280));
	notech_inv i_53567(.A(n_43558), .Z(n_44281));
	notech_inv i_53568(.A(n_43564), .Z(n_44282));
	notech_inv i_53569(.A(n_43570), .Z(n_44283));
	notech_inv i_53570(.A(n_43582), .Z(n_44285));
	notech_inv i_53571(.A(n_43588), .Z(n_44286));
	notech_inv i_53572(.A(n_43594), .Z(n_44287));
	notech_inv i_53573(.A(n_43600), .Z(n_44288));
	notech_inv i_53574(.A(n_43606), .Z(n_44289));
	notech_inv i_53575(.A(n_43612), .Z(n_44290));
	notech_inv i_53576(.A(n_43618), .Z(n_44291));
	notech_inv i_53577(.A(n_43624), .Z(n_44293));
	notech_inv i_53578(.A(n_43630), .Z(n_44294));
	notech_inv i_53579(.A(n_43636), .Z(n_44295));
	notech_inv i_53580(.A(n_43642), .Z(n_44296));
	notech_inv i_53581(.A(n_43648), .Z(n_44297));
	notech_inv i_53582(.A(n_43654), .Z(n_44299));
	notech_inv i_53583(.A(n_43660), .Z(n_44300));
	notech_inv i_53584(.A(n_43666), .Z(n_44301));
	notech_inv i_53585(.A(n_43672), .Z(n_44302));
	notech_inv i_53586(.A(n_43678), .Z(n_44303));
	notech_inv i_53587(.A(n_43684), .Z(n_44305));
	notech_inv i_53588(.A(n_43690), .Z(n_44306));
	notech_inv i_53589(.A(n_43696), .Z(n_44307));
	notech_inv i_53590(.A(n_43702), .Z(n_44308));
	notech_inv i_53591(.A(n_43708), .Z(n_44309));
	notech_inv i_53592(.A(n_43714), .Z(n_44311));
	notech_inv i_53593(.A(n_43720), .Z(n_44312));
	notech_inv i_53594(.A(n_43726), .Z(n_44313));
	notech_inv i_53595(.A(n_43732), .Z(n_44314));
	notech_inv i_53596(.A(n_43738), .Z(n_44315));
	notech_inv i_53597(.A(n_43744), .Z(n_44317));
	notech_inv i_53598(.A(n_43750), .Z(n_44318));
	notech_inv i_53599(.A(n_43756), .Z(n_44319));
	notech_inv i_53600(.A(n_43762), .Z(n_44320));
	notech_inv i_53601(.A(n_43768), .Z(n_44321));
	notech_inv i_53602(.A(n_43774), .Z(n_44323));
	notech_inv i_53603(.A(n_43780), .Z(n_44324));
	notech_inv i_53604(.A(n_43786), .Z(n_44325));
	notech_inv i_53605(.A(n_43792), .Z(n_44326));
	notech_inv i_53606(.A(n_43798), .Z(n_44327));
	notech_inv i_53607(.A(n_43804), .Z(n_44329));
	notech_inv i_53608(.A(n_43810), .Z(n_44330));
	notech_inv i_53609(.A(n_43816), .Z(n_44331));
	notech_inv i_53610(.A(n_43822), .Z(n_44332));
	notech_inv i_53611(.A(n_43828), .Z(n_44333));
	notech_inv i_53612(.A(n_43834), .Z(n_44335));
	notech_inv i_53613(.A(n_43840), .Z(n_44336));
	notech_inv i_53614(.A(n_43846), .Z(n_44337));
	notech_inv i_53615(.A(n_43852), .Z(n_44338));
	notech_inv i_53616(.A(n_43858), .Z(n_44339));
	notech_inv i_53617(.A(n_43864), .Z(n_44340));
	notech_inv i_53618(.A(n_43870), .Z(n_44341));
	notech_inv i_53619(.A(n_43876), .Z(n_44342));
	notech_inv i_53620(.A(n_43882), .Z(n_44343));
	notech_inv i_53621(.A(n_43888), .Z(n_44344));
	notech_inv i_53622(.A(n_43894), .Z(n_44345));
	notech_inv i_53623(.A(n_43900), .Z(n_44346));
	notech_inv i_53624(.A(n_43906), .Z(n_44347));
	notech_inv i_53625(.A(n_43912), .Z(n_44348));
	notech_inv i_53626(.A(n_43918), .Z(n_44349));
	notech_inv i_53627(.A(n_43924), .Z(n_44350));
	notech_inv i_53628(.A(n_43930), .Z(n_44351));
	notech_inv i_53629(.A(n_43936), .Z(n_44352));
	notech_inv i_53630(.A(n_43942), .Z(n_44353));
	notech_inv i_53631(.A(n_43948), .Z(n_44354));
	notech_inv i_53632(.A(n_43954), .Z(n_44355));
	notech_inv i_53633(.A(n_43960), .Z(n_44356));
	notech_inv i_53634(.A(n_43966), .Z(n_44357));
	notech_inv i_53635(.A(n_43972), .Z(n_44358));
	notech_inv i_53636(.A(n_43978), .Z(n_44359));
	notech_inv i_53637(.A(n_43984), .Z(n_44361));
	notech_inv i_53638(.A(n_43990), .Z(n_44362));
	notech_inv i_53639(.A(n_43996), .Z(n_44363));
	notech_inv i_53640(.A(n_44002), .Z(n_44364));
	notech_inv i_53641(.A(n_44008), .Z(n_44365));
	notech_inv i_53642(.A(n_44014), .Z(n_44366));
	notech_inv i_53643(.A(n_44020), .Z(n_44367));
	notech_inv i_53644(.A(n_44026), .Z(n_44368));
	notech_inv i_53645(.A(n_1804), .Z(n_44369));
	notech_inv i_53646(.A(displc[0]), .Z(n_44370));
	notech_inv i_53647(.A(imm_sz[0]), .Z(n_44371));
	notech_inv i_53648(.A(imm_sz[2]), .Z(n_44372));
	notech_inv i_53649(.A(pfx_sz[1]), .Z(n_44373));
	notech_inv i_53650(.A(udeco[0]), .Z(n_44374));
	notech_inv i_53651(.A(udeco[1]), .Z(n_44376));
	notech_inv i_53652(.A(udeco[2]), .Z(n_44377));
	notech_inv i_53653(.A(udeco[3]), .Z(n_44378));
	notech_inv i_53654(.A(udeco[4]), .Z(n_44379));
	notech_inv i_53655(.A(udeco[5]), .Z(n_44380));
	notech_inv i_53656(.A(udeco[6]), .Z(n_44382));
	notech_inv i_53657(.A(udeco[7]), .Z(n_44383));
	notech_inv i_53658(.A(udeco[8]), .Z(n_44384));
	notech_inv i_53659(.A(udeco[9]), .Z(n_44385));
	notech_inv i_53660(.A(udeco[10]), .Z(n_44386));
	notech_inv i_53661(.A(udeco[11]), .Z(n_44388));
	notech_inv i_53662(.A(udeco[12]), .Z(n_44389));
	notech_inv i_53663(.A(udeco[13]), .Z(n_44390));
	notech_inv i_53664(.A(udeco[14]), .Z(n_44391));
	notech_inv i_53665(.A(udeco[15]), .Z(n_44392));
	notech_inv i_53666(.A(udeco[16]), .Z(n_44394));
	notech_inv i_53667(.A(udeco[17]), .Z(n_44395));
	notech_inv i_53668(.A(udeco[18]), .Z(n_44396));
	notech_inv i_53669(.A(udeco[19]), .Z(n_44397));
	notech_inv i_53670(.A(udeco[20]), .Z(n_44398));
	notech_inv i_53671(.A(udeco[21]), .Z(n_44400));
	notech_inv i_53672(.A(udeco[22]), .Z(n_44401));
	notech_inv i_53673(.A(udeco[23]), .Z(n_44402));
	notech_inv i_53674(.A(udeco[24]), .Z(n_44403));
	notech_inv i_53675(.A(udeco[25]), .Z(n_44404));
	notech_inv i_53676(.A(udeco[26]), .Z(n_44406));
	notech_inv i_53677(.A(udeco[27]), .Z(n_44407));
	notech_inv i_53678(.A(udeco[28]), .Z(n_44408));
	notech_inv i_53679(.A(udeco[29]), .Z(n_44409));
	notech_inv i_53680(.A(udeco[30]), .Z(n_44410));
	notech_inv i_53681(.A(udeco[31]), .Z(n_44412));
	notech_inv i_53682(.A(udeco[32]), .Z(n_44413));
	notech_inv i_53683(.A(udeco[33]), .Z(n_44414));
	notech_inv i_53684(.A(udeco[34]), .Z(n_44415));
	notech_inv i_53685(.A(udeco[35]), .Z(n_44416));
	notech_inv i_53686(.A(udeco[36]), .Z(n_44418));
	notech_inv i_53687(.A(udeco[37]), .Z(n_44419));
	notech_inv i_53688(.A(udeco[38]), .Z(n_44420));
	notech_inv i_53689(.A(udeco[39]), .Z(n_44421));
	notech_inv i_53690(.A(udeco[40]), .Z(n_44422));
	notech_inv i_53691(.A(udeco[41]), .Z(n_44424));
	notech_inv i_53692(.A(udeco[42]), .Z(n_44425));
	notech_inv i_53693(.A(udeco[43]), .Z(n_44426));
	notech_inv i_53694(.A(udeco[44]), .Z(n_44427));
	notech_inv i_53695(.A(udeco[45]), .Z(n_44428));
	notech_inv i_53696(.A(udeco[46]), .Z(n_44429));
	notech_inv i_53697(.A(udeco[47]), .Z(n_44430));
	notech_inv i_53698(.A(udeco[48]), .Z(n_44431));
	notech_inv i_53699(.A(udeco[49]), .Z(n_44432));
	notech_inv i_53700(.A(udeco[50]), .Z(n_44433));
	notech_inv i_53701(.A(udeco[51]), .Z(n_44434));
	notech_inv i_53702(.A(udeco[52]), .Z(n_44436));
	notech_inv i_53703(.A(udeco[53]), .Z(n_44437));
	notech_inv i_53704(.A(udeco[54]), .Z(n_44438));
	notech_inv i_53705(.A(udeco[55]), .Z(n_44439));
	notech_inv i_53706(.A(udeco[56]), .Z(n_44440));
	notech_inv i_53707(.A(udeco[57]), .Z(n_44442));
	notech_inv i_53708(.A(udeco[58]), .Z(n_44443));
	notech_inv i_53709(.A(udeco[59]), .Z(n_44444));
	notech_inv i_53710(.A(udeco[60]), .Z(n_44445));
	notech_inv i_53711(.A(udeco[61]), .Z(n_44446));
	notech_inv i_53712(.A(udeco[62]), .Z(n_44448));
	notech_inv i_53713(.A(udeco[63]), .Z(n_44449));
	notech_inv i_53714(.A(udeco[64]), .Z(n_44450));
	notech_inv i_53715(.A(udeco[65]), .Z(n_44451));
	notech_inv i_53716(.A(udeco[66]), .Z(n_44452));
	notech_inv i_53717(.A(udeco[67]), .Z(n_44453));
	notech_inv i_53718(.A(udeco[68]), .Z(n_44454));
	notech_inv i_53719(.A(udeco[69]), .Z(n_44455));
	notech_inv i_53720(.A(udeco[70]), .Z(n_44456));
	notech_inv i_53721(.A(udeco[71]), .Z(n_44457));
	notech_inv i_53722(.A(udeco[72]), .Z(n_44458));
	notech_inv i_53723(.A(udeco[73]), .Z(n_44459));
	notech_inv i_53724(.A(udeco[74]), .Z(n_44460));
	notech_inv i_53725(.A(udeco[75]), .Z(n_44461));
	notech_inv i_53726(.A(udeco[76]), .Z(n_44462));
	notech_inv i_53727(.A(udeco[77]), .Z(n_44463));
	notech_inv i_53728(.A(udeco[78]), .Z(n_44464));
	notech_inv i_53729(.A(udeco[79]), .Z(n_44466));
	notech_inv i_53730(.A(udeco[80]), .Z(n_44467));
	notech_inv i_53731(.A(udeco[81]), .Z(n_44468));
	notech_inv i_53732(.A(udeco[82]), .Z(n_44469));
	notech_inv i_53733(.A(udeco[83]), .Z(n_44470));
	notech_inv i_53734(.A(udeco[84]), .Z(n_44472));
	notech_inv i_53735(.A(udeco[85]), .Z(n_44473));
	notech_inv i_53736(.A(udeco[86]), .Z(n_44474));
	notech_inv i_53737(.A(udeco[87]), .Z(n_44475));
	notech_inv i_53738(.A(udeco[88]), .Z(n_44476));
	notech_inv i_53739(.A(udeco[89]), .Z(n_44478));
	notech_inv i_53740(.A(udeco[90]), .Z(n_44479));
	notech_inv i_53741(.A(udeco[91]), .Z(n_44480));
	notech_inv i_53742(.A(udeco[92]), .Z(n_44481));
	notech_inv i_53743(.A(udeco[93]), .Z(n_44482));
	notech_inv i_53744(.A(udeco[94]), .Z(n_44484));
	notech_inv i_53745(.A(udeco[95]), .Z(n_44485));
	notech_inv i_53746(.A(udeco[96]), .Z(n_44486));
	notech_inv i_53747(.A(udeco[97]), .Z(n_44487));
	notech_inv i_53748(.A(udeco[98]), .Z(n_44488));
	notech_inv i_53749(.A(udeco[99]), .Z(n_44490));
	notech_inv i_53750(.A(udeco[100]), .Z(n_44491));
	notech_inv i_53751(.A(udeco[101]), .Z(n_44492));
	notech_inv i_53752(.A(udeco[102]), .Z(n_44493));
	notech_inv i_53753(.A(udeco[103]), .Z(n_44494));
	notech_inv i_53754(.A(udeco[104]), .Z(n_44496));
	notech_inv i_53755(.A(udeco[105]), .Z(n_44497));
	notech_inv i_53756(.A(udeco[106]), .Z(n_44498));
	notech_inv i_53757(.A(udeco[107]), .Z(n_44499));
	notech_inv i_53758(.A(udeco[108]), .Z(n_44500));
	notech_inv i_53759(.A(udeco[109]), .Z(n_44501));
	notech_inv i_53760(.A(udeco[110]), .Z(n_44502));
	notech_inv i_53761(.A(udeco[111]), .Z(n_44503));
	notech_inv i_53762(.A(udeco[112]), .Z(n_44504));
	notech_inv i_53763(.A(udeco[113]), .Z(n_44505));
	notech_inv i_53764(.A(udeco[114]), .Z(n_44506));
	notech_inv i_53765(.A(udeco[115]), .Z(n_44508));
	notech_inv i_53766(.A(udeco[116]), .Z(n_44509));
	notech_inv i_53767(.A(udeco[117]), .Z(n_44510));
	notech_inv i_53768(.A(udeco[118]), .Z(n_44511));
	notech_inv i_53769(.A(udeco[119]), .Z(n_44512));
	notech_inv i_53770(.A(udeco[120]), .Z(n_44514));
	notech_inv i_53771(.A(udeco[121]), .Z(n_44515));
	notech_inv i_53772(.A(udeco[122]), .Z(n_44516));
	notech_inv i_53773(.A(udeco[123]), .Z(n_44517));
	notech_inv i_53774(.A(udeco[124]), .Z(n_44518));
	notech_inv i_53775(.A(udeco[125]), .Z(n_44520));
	notech_inv i_53776(.A(udeco[126]), .Z(n_44521));
	notech_inv i_53777(.A(udeco[127]), .Z(n_44522));
	notech_inv i_53778(.A(opz[0]), .Z(n_44523));
	notech_inv i_53779(.A(opz[1]), .Z(n_44524));
	notech_inv i_53780(.A(in128[16]), .Z(n_44525));
	notech_inv i_53781(.A(in128[17]), .Z(n_44526));
	notech_inv i_53782(.A(in128[18]), .Z(n_44527));
	notech_inv i_53783(.A(in128[19]), .Z(n_44528));
	notech_inv i_53784(.A(in128[20]), .Z(n_44529));
	notech_inv i_53785(.A(in128[21]), .Z(n_44530));
	notech_inv i_53786(.A(in128[22]), .Z(n_44532));
	notech_inv i_53787(.A(in128[23]), .Z(n_44533));
	notech_inv i_53788(.A(in128[24]), .Z(n_44534));
	notech_inv i_53789(.A(in128[25]), .Z(n_44535));
	notech_inv i_53790(.A(in128[26]), .Z(n_44536));
	notech_inv i_53791(.A(in128[27]), .Z(n_44538));
	notech_inv i_53792(.A(in128[28]), .Z(n_44539));
	notech_inv i_53793(.A(in128[29]), .Z(n_44540));
	notech_inv i_53794(.A(in128[30]), .Z(n_44541));
	notech_inv i_53795(.A(in128[31]), .Z(n_44542));
	notech_inv i_53796(.A(in128[32]), .Z(n_44544));
	notech_inv i_53797(.A(in128[33]), .Z(n_44545));
	notech_inv i_53798(.A(in128[34]), .Z(n_44546));
	notech_inv i_53799(.A(in128[35]), .Z(n_44547));
	notech_inv i_53800(.A(in128[36]), .Z(n_44548));
	notech_inv i_53801(.A(in128[37]), .Z(n_44550));
	notech_inv i_53802(.A(in128[38]), .Z(n_44551));
	notech_inv i_53803(.A(in128[39]), .Z(n_44552));
	notech_inv i_53804(.A(in128[40]), .Z(n_44553));
	notech_inv i_53805(.A(in128[41]), .Z(n_44554));
	notech_inv i_53806(.A(in128[42]), .Z(n_44556));
	notech_inv i_53807(.A(in128[43]), .Z(n_44557));
	notech_inv i_53808(.A(in128[44]), .Z(n_44558));
	notech_inv i_53809(.A(in128[45]), .Z(n_44559));
	notech_inv i_53810(.A(in128[46]), .Z(n_44560));
	notech_inv i_53811(.A(in128[47]), .Z(n_44562));
	notech_inv i_53812(.A(in128[48]), .Z(n_44563));
	notech_inv i_53813(.A(in128[49]), .Z(n_44564));
	notech_inv i_53814(.A(in128[50]), .Z(n_44565));
	notech_inv i_53815(.A(in128[51]), .Z(n_44566));
	notech_inv i_53816(.A(in128[52]), .Z(n_44568));
	notech_inv i_53817(.A(in128[53]), .Z(n_44569));
	notech_inv i_53818(.A(in128[54]), .Z(n_44570));
	notech_inv i_53819(.A(in128[55]), .Z(n_44571));
	notech_inv i_53820(.A(in128[56]), .Z(n_44572));
	notech_inv i_53821(.A(in128[57]), .Z(n_44574));
	notech_inv i_53822(.A(in128[58]), .Z(n_44575));
	notech_inv i_53823(.A(in128[59]), .Z(n_44576));
	notech_inv i_53824(.A(in128[60]), .Z(n_44577));
	notech_inv i_53825(.A(in128[61]), .Z(n_44578));
	notech_inv i_53826(.A(in128[62]), .Z(n_44580));
	notech_inv i_53827(.A(in128[63]), .Z(n_44581));
	notech_inv i_53828(.A(in128[64]), .Z(n_44582));
	notech_inv i_53829(.A(in128[65]), .Z(n_44583));
	notech_inv i_53830(.A(in128[66]), .Z(n_44584));
	notech_inv i_53831(.A(in128[67]), .Z(n_44586));
	notech_inv i_53832(.A(in128[68]), .Z(n_44587));
	notech_inv i_53833(.A(in128[69]), .Z(n_44588));
	notech_inv i_53834(.A(in128[70]), .Z(n_44589));
	notech_inv i_53835(.A(in128[71]), .Z(n_44590));
	notech_inv i_53836(.A(in128[72]), .Z(n_44592));
	notech_inv i_53837(.A(in128[73]), .Z(n_44593));
	notech_inv i_53838(.A(in128[74]), .Z(n_44594));
	notech_inv i_53839(.A(in128[75]), .Z(n_44595));
	notech_inv i_53840(.A(in128[76]), .Z(n_44596));
	notech_inv i_53841(.A(in128[77]), .Z(n_44598));
	notech_inv i_53842(.A(in128[78]), .Z(n_44599));
	notech_inv i_53843(.A(in128[79]), .Z(n_44600));
	notech_inv i_53844(.A(in128[80]), .Z(n_44601));
	notech_inv i_53845(.A(in128[81]), .Z(n_44602));
	notech_inv i_53846(.A(in128[82]), .Z(n_44604));
	notech_inv i_53847(.A(in128[83]), .Z(n_44605));
	notech_inv i_53848(.A(in128[84]), .Z(n_44606));
	notech_inv i_53849(.A(in128[85]), .Z(n_44607));
	notech_inv i_53850(.A(in128[86]), .Z(n_44608));
	notech_inv i_53851(.A(in128[87]), .Z(n_44610));
	notech_inv i_53852(.A(in128[88]), .Z(n_44611));
	notech_inv i_53853(.A(in128[89]), .Z(n_44612));
	notech_inv i_53854(.A(in128[90]), .Z(n_44613));
	notech_inv i_53855(.A(in128[91]), .Z(n_44614));
	notech_inv i_53856(.A(in128[92]), .Z(n_44616));
	notech_inv i_53857(.A(in128[93]), .Z(n_44617));
	notech_inv i_53858(.A(in128[94]), .Z(n_44618));
	notech_inv i_53859(.A(in128[95]), .Z(n_44619));
	notech_inv i_53860(.A(in128[96]), .Z(n_44620));
	notech_inv i_53861(.A(in128[97]), .Z(n_44622));
	notech_inv i_53862(.A(in128[98]), .Z(n_44623));
	notech_inv i_53863(.A(in128[99]), .Z(n_44624));
	notech_inv i_53864(.A(in128[100]), .Z(n_44625));
	notech_inv i_53865(.A(in128[101]), .Z(n_44626));
	notech_inv i_53866(.A(in128[102]), .Z(n_44628));
	notech_inv i_53867(.A(in128[103]), .Z(n_44629));
	notech_inv i_53868(.A(in128[104]), .Z(n_44630));
	notech_inv i_53869(.A(in128[105]), .Z(n_44631));
	notech_inv i_53870(.A(in128[106]), .Z(n_44632));
	notech_inv i_53871(.A(in128[107]), .Z(n_44634));
	notech_inv i_53872(.A(in128[108]), .Z(n_44635));
	notech_inv i_53873(.A(in128[109]), .Z(n_44636));
	notech_inv i_53874(.A(in128[110]), .Z(n_44637));
	notech_inv i_53875(.A(in128[111]), .Z(n_44638));
	notech_inv i_53876(.A(in128[112]), .Z(n_44640));
	notech_inv i_53877(.A(in128[113]), .Z(n_44641));
	notech_inv i_53878(.A(in128[114]), .Z(n_44642));
	notech_inv i_53879(.A(in128[115]), .Z(n_44643));
	notech_inv i_53880(.A(in128[116]), .Z(n_44644));
	notech_inv i_53881(.A(in128[117]), .Z(n_44646));
	notech_inv i_53882(.A(in128[118]), .Z(n_44647));
	notech_inv i_53883(.A(in128[119]), .Z(n_44648));
	notech_inv i_53884(.A(in128[120]), .Z(n_44649));
	notech_inv i_53885(.A(in128[121]), .Z(n_44650));
	notech_inv i_53886(.A(in128[122]), .Z(n_44652));
	notech_inv i_53887(.A(in128[123]), .Z(n_44653));
	notech_inv i_53888(.A(in128[124]), .Z(n_44654));
	notech_inv i_53889(.A(in128[125]), .Z(n_44655));
	notech_inv i_53890(.A(in128[126]), .Z(n_44656));
	notech_inv i_53891(.A(in128[127]), .Z(n_44658));
	notech_inv i_53892(.A(in128[0]), .Z(n_44659));
	notech_inv i_53893(.A(\to_acu2_0[77] ), .Z(n_44660));
	notech_inv i_53894(.A(\to_acu2_0[67] ), .Z(n_44661));
	notech_inv i_53895(.A(\to_acu2_0[65] ), .Z(n_44662));
	notech_inv i_53896(.A(\to_acu2_0[64] ), .Z(n_44663));
	notech_inv i_53897(.A(\to_acu2_0[32] ), .Z(n_44664));
	notech_inv i_53898(.A(\to_acu2_0[31] ), .Z(n_44665));
	notech_inv i_53899(.A(\to_acu2_0[66] ), .Z(n_44666));
	notech_inv i_53900(.A(\to_acu2_0[63] ), .Z(n_44667));
	notech_inv i_53901(.A(\to_acu2_0[60] ), .Z(n_44668));
	notech_inv i_53902(.A(\to_acu2_0[49] ), .Z(n_44669));
	notech_inv i_53903(.A(\to_acu2_0[33] ), .Z(n_44670));
	notech_inv i_53904(.A(\to_acu2_0[71] ), .Z(n_44671));
	notech_inv i_53905(.A(\to_acu2_0[70] ), .Z(n_44672));
	notech_inv i_53906(.A(\to_acu2_0[75] ), .Z(n_44673));
	notech_inv i_53907(.A(in128[7]), .Z(n_44674));
	notech_inv i_53908(.A(in128[6]), .Z(n_44675));
	notech_inv i_53909(.A(in128[5]), .Z(n_44676));
	notech_inv i_53910(.A(in128[4]), .Z(n_44677));
	notech_inv i_53911(.A(in128[3]), .Z(n_44678));
	notech_inv i_53912(.A(\to_acu2_0[80] ), .Z(n_44679));
	notech_inv i_53913(.A(\to_acu2_0[56] ), .Z(n_44680));
	notech_inv i_53914(.A(\to_acu2_0[50] ), .Z(n_44681));
	notech_inv i_53915(.A(\to_acu2_0[76] ), .Z(n_44682));
	notech_inv i_53916(.A(\to_acu2_0[72] ), .Z(n_44683));
	notech_inv i_53917(.A(\to_acu2_0[73] ), .Z(n_44684));
	notech_inv i_53918(.A(\to_acu2_0[74] ), .Z(n_44685));
	notech_inv i_53919(.A(\to_acu2_0[58] ), .Z(n_44686));
	notech_inv i_53920(.A(\to_acu2_0[57] ), .Z(n_44687));
	notech_inv i_53921(.A(\to_acu2_0[52] ), .Z(n_44688));
	notech_inv i_53922(.A(\to_acu2_0[51] ), .Z(n_44689));
	notech_inv i_53923(.A(\to_acu2_0[53] ), .Z(n_44690));
	notech_inv i_53924(.A(\to_acu2_0[55] ), .Z(n_44691));
	notech_inv i_53925(.A(\to_acu2_0[59] ), .Z(n_44692));
	notech_inv i_53926(.A(\to_acu2_0[48] ), .Z(n_44693));
	notech_inv i_53927(.A(\to_acu2_0[35] ), .Z(n_44694));
	notech_inv i_53928(.A(\to_acu2_0[34] ), .Z(n_44695));
	notech_inv i_53929(.A(\to_acu2_0[37] ), .Z(n_44696));
	notech_inv i_53930(.A(\to_acu2_0[36] ), .Z(n_44697));
	notech_inv i_53931(.A(\to_acu2_0[40] ), .Z(n_44698));
	notech_inv i_53932(.A(\to_acu2_0[38] ), .Z(n_44699));
	notech_inv i_53933(.A(\to_acu2_0[43] ), .Z(n_44700));
	notech_inv i_53934(.A(\to_acu2_0[42] ), .Z(n_44701));
	notech_inv i_53935(.A(\to_acu2_0[44] ), .Z(n_44702));
	notech_inv i_53936(.A(\to_acu2_0[46] ), .Z(n_44703));
	notech_inv i_53937(.A(\to_acu2_0[47] ), .Z(n_44704));
	notech_inv i_53938(.A(\to_acu2_0[79] ), .Z(n_44705));
	notech_inv i_53939(.A(\to_acu2_0[61] ), .Z(n_44706));
	notech_inv i_53940(.A(\to_acu2_0[78] ), .Z(n_44707));
	notech_inv i_53941(.A(in128[13]), .Z(n_44708));
	notech_inv i_53942(.A(in128[12]), .Z(n_44709));
	notech_inv i_53943(.A(in128[11]), .Z(n_44710));
	notech_inv i_53944(.A(\to_acu2_0[15] ), .Z(n_44711));
	notech_inv i_53945(.A(\to_acu2_0[14] ), .Z(n_44712));
	notech_inv i_53946(.A(\to_acu2_0[13] ), .Z(n_44713));
	notech_inv i_53947(.A(\to_acu2_0[18] ), .Z(n_44714));
	notech_inv i_53948(.A(\to_acu2_0[17] ), .Z(n_44715));
	notech_inv i_53949(.A(\to_acu2_0[12] ), .Z(n_44716));
	notech_inv i_53950(.A(\to_acu2_0[68] ), .Z(n_44717));
	notech_inv i_53951(.A(\to_acu2_0[16] ), .Z(n_44718));
	notech_inv i_53952(.A(in128[15]), .Z(n_44719));
	notech_inv i_53953(.A(n_59489), .Z(n_44720));
	notech_inv i_53954(.A(in128[14]), .Z(n_44721));
	notech_inv i_53955(.A(in128[8]), .Z(n_44722));
	notech_inv i_53956(.A(in128[9]), .Z(n_44723));
	notech_inv i_53957(.A(\to_acu2_0[62] ), .Z(n_44724));
	notech_inv i_53958(.A(\to_acu2_0[69] ), .Z(n_44725));
	notech_inv i_53959(.A(\to_acu2_0[8] ), .Z(n_44726));
	notech_inv i_53960(.A(\to_acu2_0[11] ), .Z(n_44727));
	notech_inv i_53961(.A(\to_acu2_0[9] ), .Z(n_44728));
	notech_inv i_53962(.A(fpu), .Z(n_44729));
	notech_inv i_53963(.A(sib_dec), .Z(n_44730));
	notech_inv i_53964(.A(mod_dec), .Z(n_44731));
	notech_inv i_53965(.A(\to_acu2_0[54] ), .Z(n_44732));
	notech_inv i_53966(.A(\to_acu2_0[6] ), .Z(n_44733));
	notech_inv i_53967(.A(\to_acu2_0[5] ), .Z(n_44734));
	notech_inv i_53968(.A(\to_acu2_0[1] ), .Z(n_44735));
	notech_inv i_53969(.A(in128[1]), .Z(n_44736));
	notech_inv i_53970(.A(in128[2]), .Z(n_44737));
	notech_inv i_53971(.A(pc_req), .Z(n_44738));
	notech_inv i_53972(.A(\nbus_12406[0] ), .Z(n_44739));
	notech_inv i_53973(.A(\to_acu2_0[22] ), .Z(n_44740));
	notech_inv i_53974(.A(\to_acu2_0[23] ), .Z(n_44741));
	notech_inv i_53975(.A(\to_acu2_0[21] ), .Z(n_44742));
	notech_inv i_53976(.A(\to_acu2_0[26] ), .Z(n_44743));
	notech_inv i_53977(.A(pg_fault), .Z(n_44744));
	notech_inv i_53978(.A(twobyte), .Z(n_44745));
	notech_inv i_53979(.A(\to_acu2_0[27] ), .Z(n_44746));
	notech_inv i_53980(.A(\to_acu2_0[3] ), .Z(n_44747));
	notech_inv i_53981(.A(\to_acu2_0[2] ), .Z(n_44748));
	notech_inv i_53982(.A(\to_acu2_0[41] ), .Z(n_44749));
	notech_inv i_53983(.A(\to_acu2_0[45] ), .Z(n_44750));
	notech_inv i_53984(.A(\to_acu2_0[4] ), .Z(n_44751));
	notech_inv i_53985(.A(\to_acu2_0[10] ), .Z(n_44752));
	notech_inv i_53986(.A(\to_acu2_0[19] ), .Z(n_44753));
	notech_inv i_53987(.A(\to_acu2_0[20] ), .Z(n_44754));
	notech_inv i_53988(.A(\to_acu2_0[25] ), .Z(n_44755));
	notech_inv i_53989(.A(\to_acu2_0[24] ), .Z(n_44756));
	notech_inv i_53990(.A(\to_acu2_0[28] ), .Z(n_44757));
	notech_inv i_53991(.A(\to_acu2_0[0] ), .Z(n_44758));
	notech_inv i_53992(.A(\to_acu2_0[7] ), .Z(n_44759));
	notech_inv i_53993(.A(adz), .Z(n_44760));
	notech_inv i_53994(.A(\nbus_12406[1] ), .Z(n_44761));
	notech_inv i_53995(.A(\nbus_12406[2] ), .Z(n_44762));
	notech_inv i_53996(.A(\nbus_12406[3] ), .Z(n_44763));
	notech_inv i_53997(.A(\nbus_12406[4] ), .Z(n_44764));
	notech_inv i_53998(.A(\nbus_12406[5] ), .Z(n_44765));
	notech_inv i_53999(.A(\to_acu2_0[29] ), .Z(n_44766));
	notech_inv i_54000(.A(\to_acu2_0[30] ), .Z(n_44767));
	notech_inv i_54001(.A(int_main), .Z(n_44768));
	deco8 i_deco_1(.in8({in128[7], in128[6], in128[5], in128[4], in128[3], in128
		[2], in128[1], in128[0]}), .indic({\to_acu2_0[80] , \to_acu2_0[79] 
		, \to_acu2_0[78] , \to_acu2_0[77] , \to_acu2_0[76] , \to_acu2_0[75] 
		, \to_acu2_0[74] , \to_acu2_0[73] , \to_acu2_0[72] , \to_acu2_0[71] 
		, \to_acu2_0[70] , \to_acu2_0[69] , \to_acu2_0[68] , \to_acu2_0[67] 
		, \to_acu2_0[66] , \to_acu2_0[65] , \to_acu2_0[64] , \to_acu2_0[63] 
		, \to_acu2_0[62] , \to_acu2_0[61] , \to_acu2_0[60] , \to_acu2_0[59] 
		, \to_acu2_0[58] , \to_acu2_0[57] , \to_acu2_0[56] , \to_acu2_0[55] 
		, \to_acu2_0[54] , \to_acu2_0[53] , \to_acu2_0[52] , \to_acu2_0[51] 
		, \to_acu2_0[50] , \to_acu2_0[49] , \to_acu2_0[48] , \to_acu2_0[47] 
		, \to_acu2_0[46] , \to_acu2_0[45] , \to_acu2_0[44] , \to_acu2_0[43] 
		, \to_acu2_0[42] , \to_acu2_0[41] , \to_acu2_0[40] , 
		UNCONNECTED_000, \to_acu2_0[38] , \to_acu2_0[37] , \to_acu2_0[36] 
		, \to_acu2_0[35] , \to_acu2_0[34] , \to_acu2_0[33] , \to_acu2_0[32] 
		, \to_acu2_0[31] , \to_acu2_0[30] , \to_acu2_0[29] , \to_acu2_0[28] 
		, \to_acu2_0[27] , \to_acu2_0[26] , \to_acu2_0[25] , \to_acu2_0[24] 
		, \to_acu2_0[23] , \to_acu2_0[22] , \to_acu2_0[21] , \to_acu2_0[20] 
		, \to_acu2_0[19] , \to_acu2_0[18] , \to_acu2_0[17] , \to_acu2_0[16] 
		, \to_acu2_0[15] , \to_acu2_0[14] , \to_acu2_0[13] , \to_acu2_0[12] 
		, \to_acu2_0[11] , \to_acu2_0[10] , \to_acu2_0[9] , \to_acu2_0[8] 
		}));
	udecox i_udeco(.op({in128[7], in128[6], in128[5], in128[4], in128[3], in128
		[2], in128[1], in128[0]}), .modrm({in128[15], in128[14], in128[
		13], in128[12], in128[11], n_59489, in128[9], in128[8]}), .twobyte
		(twobyte), .cpl(cpl), .adz(adz), .opz(opz), .udeco(udeco), .fpu(fpu
		), .emul(cr0[2]), .ipg_fault(ipg_fault));
	deco_rm i_deco_3(.in8({in128[15], in128[14], in128[13], in128[12], 
		UNCONNECTED_001, n_59488, in128[9], in128[8]}), .indic({\to_acu2_0[7] 
		, \to_acu2_0[6] , \to_acu2_0[5] , \to_acu2_0[4] , \to_acu2_0[3] 
		, \to_acu2_0[2] , \to_acu2_0[1] , \to_acu2_0[0] }));
	AWDP_partition_5 i_65646(.O0({\nbus_12406[5] , \nbus_12406[4] , \nbus_12406[3] 
		, \nbus_12406[2] , \nbus_12406[1] , \nbus_12406[0] }), .pfx_sz(pfx_sz
		), .twobyte(twobyte), .fpu(fpu), .sib_dec(sib_dec), .displc(displc
		), .mod_dec(mod_dec), .imm_sz(imm_sz));
endmodule
module AWDP_ADD_101(O0, opa, opd);
    output [8:0] O0;
    input [7:0] opa;
    input [7:0] opd;
    // Line 601
    wire [8:0] O0;
    // Line 601
    wire [8:0] N54;

    // Line 601
    assign O0 = N54;
    // Line 601
    assign N54 = opa + opd;
endmodule

module AWDP_ADD_103(O0, opa, opd);
    output [16:0] O0;
    input [15:0] opa;
    input [15:0] opd;
    // Line 600
    wire [16:0] O0;
    // Line 600
    wire [16:0] N63;

    // Line 600
    assign O0 = N63;
    // Line 600
    assign N63 = opa + opd;
endmodule

module AWDP_ADD_107(O0, opd, I0);

	output [31:0] O0;
	input [31:0] opd;
	input [31:0] I0;

	wire \opd[2] ;
	wire \opd[3] ;
	wire \opd[4] ;
	wire \opd[5] ;
	wire \opd[6] ;
	wire \opd[7] ;
	wire \opd[8] ;
	wire \opd[9] ;
	wire \opd[10] ;
	wire \opd[11] ;
	wire \opd[12] ;
	wire \opd[13] ;
	wire \opd[14] ;
	wire \opd[15] ;
	wire \opd[16] ;
	wire \opd[17] ;
	wire \opd[18] ;
	wire \opd[19] ;
	wire \opd[20] ;
	wire \opd[21] ;
	wire \opd[22] ;
	wire \opd[23] ;
	wire \opd[24] ;
	wire \opd[25] ;
	wire \opd[26] ;
	wire \opd[27] ;
	wire \opd[28] ;
	wire \opd[29] ;
	wire \opd[30] ;
	wire \opd[31] ;


	assign O0[0] = opd[0];
	assign O0[1] = opd[1];
	assign \opd[2]  = opd[2];
	assign \opd[3]  = opd[3];
	assign \opd[4]  = opd[4];
	assign \opd[5]  = opd[5];
	assign \opd[6]  = opd[6];
	assign \opd[7]  = opd[7];
	assign \opd[8]  = opd[8];
	assign \opd[9]  = opd[9];
	assign \opd[10]  = opd[10];
	assign \opd[11]  = opd[11];
	assign \opd[12]  = opd[12];
	assign \opd[13]  = opd[13];
	assign \opd[14]  = opd[14];
	assign \opd[15]  = opd[15];
	assign \opd[16]  = opd[16];
	assign \opd[17]  = opd[17];
	assign \opd[18]  = opd[18];
	assign \opd[19]  = opd[19];
	assign \opd[20]  = opd[20];
	assign \opd[21]  = opd[21];
	assign \opd[22]  = opd[22];
	assign \opd[23]  = opd[23];
	assign \opd[24]  = opd[24];
	assign \opd[25]  = opd[25];
	assign \opd[26]  = opd[26];
	assign \opd[27]  = opd[27];
	assign \opd[28]  = opd[28];
	assign \opd[29]  = opd[29];
	assign \opd[30]  = opd[30];
	assign \opd[31]  = opd[31];

	notech_ha2 i_29(.A(\opd[31] ), .B(n_354), .Z(O0[31]));
	notech_ha2 i_28(.A(\opd[30] ), .B(n_352), .Z(O0[30]), .CO(n_354));
	notech_ha2 i_27(.A(\opd[29] ), .B(n_341), .Z(O0[29]), .CO(n_352));
	notech_fa2 i_26(.A(I0[28]), .B(n_339), .CI(\opd[28] ), .Z(O0[28]), .CO(n_341
		));
	notech_fa2 i_25(.A(I0[27]), .B(n_337), .CI(\opd[27] ), .Z(O0[27]), .CO(n_339
		));
	notech_fa2 i_24(.A(I0[26]), .B(n_335), .CI(\opd[26] ), .Z(O0[26]), .CO(n_337
		));
	notech_fa2 i_23(.A(I0[25]), .B(n_333), .CI(\opd[25] ), .Z(O0[25]), .CO(n_335
		));
	notech_fa2 i_22(.A(I0[24]), .B(n_331), .CI(\opd[24] ), .Z(O0[24]), .CO(n_333
		));
	notech_fa2 i_21(.A(I0[23]), .B(n_329), .CI(\opd[23] ), .Z(O0[23]), .CO(n_331
		));
	notech_fa2 i_20(.A(I0[22]), .B(n_327), .CI(\opd[22] ), .Z(O0[22]), .CO(n_329
		));
	notech_fa2 i_19(.A(I0[21]), .B(n_325), .CI(\opd[21] ), .Z(O0[21]), .CO(n_327
		));
	notech_fa2 i_18(.A(I0[20]), .B(n_323), .CI(\opd[20] ), .Z(O0[20]), .CO(n_325
		));
	notech_fa2 i_17(.A(I0[19]), .B(n_321), .CI(\opd[19] ), .Z(O0[19]), .CO(n_323
		));
	notech_fa2 i_16(.A(I0[18]), .B(n_319), .CI(\opd[18] ), .Z(O0[18]), .CO(n_321
		));
	notech_fa2 i_15(.A(I0[17]), .B(n_317), .CI(\opd[17] ), .Z(O0[17]), .CO(n_319
		));
	notech_fa2 i_14(.A(I0[16]), .B(n_315), .CI(\opd[16] ), .Z(O0[16]), .CO(n_317
		));
	notech_fa2 i_13(.A(I0[15]), .B(n_313), .CI(\opd[15] ), .Z(O0[15]), .CO(n_315
		));
	notech_fa2 i_12(.A(I0[14]), .B(n_311), .CI(\opd[14] ), .Z(O0[14]), .CO(n_313
		));
	notech_fa2 i_11(.A(I0[13]), .B(n_309), .CI(\opd[13] ), .Z(O0[13]), .CO(n_311
		));
	notech_fa2 i_10(.A(I0[12]), .B(n_307), .CI(\opd[12] ), .Z(O0[12]), .CO(n_309
		));
	notech_fa2 i_9(.A(I0[11]), .B(n_305), .CI(\opd[11] ), .Z(O0[11]), .CO(n_307
		));
	notech_fa2 i_8(.A(I0[10]), .B(n_303), .CI(\opd[10] ), .Z(O0[10]), .CO(n_305
		));
	notech_fa2 i_7(.A(I0[9]), .B(n_301), .CI(\opd[9] ), .Z(O0[9]), .CO(n_303
		));
	notech_fa2 i_6(.A(I0[8]), .B(n_299), .CI(\opd[8] ), .Z(O0[8]), .CO(n_301
		));
	notech_fa2 i_5(.A(I0[7]), .B(n_297), .CI(\opd[7] ), .Z(O0[7]), .CO(n_299
		));
	notech_fa2 i_4(.A(I0[6]), .B(n_295), .CI(\opd[6] ), .Z(O0[6]), .CO(n_297
		));
	notech_fa2 i_3(.A(I0[5]), .B(n_293), .CI(\opd[5] ), .Z(O0[5]), .CO(n_295
		));
	notech_fa2 i_2(.A(I0[4]), .B(n_291), .CI(\opd[4] ), .Z(O0[4]), .CO(n_293
		));
	notech_fa2 i_1(.A(I0[3]), .B(n_350), .CI(\opd[3] ), .Z(O0[3]), .CO(n_291
		));
	notech_ha2 i_0(.A(I0[2]), .B(\opd[2] ), .Z(O0[2]), .CO(n_350));
endmodule
module AWDP_ADD_11(O0, opc, I0);
    output [31:0] O0;
    input [31:0] opc;
    input [31:0] I0;
    // Line 1006
    wire [31:0] O0;
    // Line 1006
    wire [31:0] N87;

    // Line 1006
    assign O0 = N87;
    // Line 1006
    assign N87 = opc + I0;
endmodule

module AWDP_ADD_110(O0, regs_4, calc_sz);
    output [31:0] O0;
    input [31:0] regs_4;
    input [2:0] calc_sz;
    // Line 470
    wire [31:0] N98;
    // Line 348
    wire [31:0] O0;

    // Line 470
    assign N98 = calc_sz + regs_4;
    // Line 348
    assign O0 = N98;
endmodule

module AWDP_ADD_117(O0, idtr, I0);

	output [31:0] O0;
	input [31:0] idtr;
	input [18:0] I0;

	wire \idtr[3] ;
	wire \idtr[4] ;
	wire \idtr[5] ;
	wire \idtr[6] ;
	wire \idtr[7] ;
	wire \idtr[8] ;
	wire \idtr[9] ;
	wire \idtr[10] ;
	wire \idtr[11] ;
	wire \idtr[12] ;
	wire \idtr[13] ;
	wire \idtr[14] ;
	wire \idtr[15] ;
	wire \idtr[16] ;
	wire \idtr[17] ;
	wire \idtr[18] ;
	wire \idtr[19] ;
	wire \idtr[20] ;
	wire \idtr[21] ;
	wire \idtr[22] ;
	wire \idtr[23] ;
	wire \idtr[24] ;
	wire \idtr[25] ;
	wire \idtr[26] ;
	wire \idtr[27] ;
	wire \idtr[28] ;
	wire \idtr[29] ;
	wire \idtr[30] ;
	wire \idtr[31] ;


	assign O0[0] = idtr[0];
	assign O0[1] = idtr[1];
	assign O0[2] = idtr[2];
	assign \idtr[3]  = idtr[3];
	assign \idtr[4]  = idtr[4];
	assign \idtr[5]  = idtr[5];
	assign \idtr[6]  = idtr[6];
	assign \idtr[7]  = idtr[7];
	assign \idtr[8]  = idtr[8];
	assign \idtr[9]  = idtr[9];
	assign \idtr[10]  = idtr[10];
	assign \idtr[11]  = idtr[11];
	assign \idtr[12]  = idtr[12];
	assign \idtr[13]  = idtr[13];
	assign \idtr[14]  = idtr[14];
	assign \idtr[15]  = idtr[15];
	assign \idtr[16]  = idtr[16];
	assign \idtr[17]  = idtr[17];
	assign \idtr[18]  = idtr[18];
	assign \idtr[19]  = idtr[19];
	assign \idtr[20]  = idtr[20];
	assign \idtr[21]  = idtr[21];
	assign \idtr[22]  = idtr[22];
	assign \idtr[23]  = idtr[23];
	assign \idtr[24]  = idtr[24];
	assign \idtr[25]  = idtr[25];
	assign \idtr[26]  = idtr[26];
	assign \idtr[27]  = idtr[27];
	assign \idtr[28]  = idtr[28];
	assign \idtr[29]  = idtr[29];
	assign \idtr[30]  = idtr[30];
	assign \idtr[31]  = idtr[31];

	notech_ha2 i_28(.A(\idtr[31] ), .B(n_346), .Z(O0[31]));
	notech_ha2 i_27(.A(\idtr[30] ), .B(n_344), .Z(O0[30]), .CO(n_346));
	notech_ha2 i_26(.A(\idtr[29] ), .B(n_342), .Z(O0[29]), .CO(n_344));
	notech_ha2 i_25(.A(\idtr[28] ), .B(n_340), .Z(O0[28]), .CO(n_342));
	notech_ha2 i_24(.A(\idtr[27] ), .B(n_338), .Z(O0[27]), .CO(n_340));
	notech_ha2 i_23(.A(\idtr[26] ), .B(n_336), .Z(O0[26]), .CO(n_338));
	notech_ha2 i_22(.A(\idtr[25] ), .B(n_334), .Z(O0[25]), .CO(n_336));
	notech_ha2 i_21(.A(\idtr[24] ), .B(n_332), .Z(O0[24]), .CO(n_334));
	notech_ha2 i_20(.A(\idtr[23] ), .B(n_330), .Z(O0[23]), .CO(n_332));
	notech_ha2 i_19(.A(\idtr[22] ), .B(n_328), .Z(O0[22]), .CO(n_330));
	notech_ha2 i_18(.A(\idtr[21] ), .B(n_326), .Z(O0[21]), .CO(n_328));
	notech_ha2 i_17(.A(\idtr[20] ), .B(n_324), .Z(O0[20]), .CO(n_326));
	notech_ha2 i_16(.A(\idtr[19] ), .B(n_293), .Z(O0[19]), .CO(n_324));
	notech_fa2 i_15(.A(I0[18]), .B(n_291), .CI(\idtr[18] ), .Z(O0[18]), .CO(n_293
		));
	notech_fa2 i_14(.A(I0[17]), .B(n_289), .CI(\idtr[17] ), .Z(O0[17]), .CO(n_291
		));
	notech_fa2 i_13(.A(I0[16]), .B(n_287), .CI(\idtr[16] ), .Z(O0[16]), .CO(n_289
		));
	notech_fa2 i_12(.A(I0[15]), .B(n_285), .CI(\idtr[15] ), .Z(O0[15]), .CO(n_287
		));
	notech_fa2 i_11(.A(I0[14]), .B(n_283), .CI(\idtr[14] ), .Z(O0[14]), .CO(n_285
		));
	notech_fa2 i_10(.A(I0[13]), .B(n_281), .CI(\idtr[13] ), .Z(O0[13]), .CO(n_283
		));
	notech_fa2 i_9(.A(I0[12]), .B(n_279), .CI(\idtr[12] ), .Z(O0[12]), .CO(n_281
		));
	notech_fa2 i_8(.A(I0[11]), .B(n_277), .CI(\idtr[11] ), .Z(O0[11]), .CO(n_279
		));
	notech_fa2 i_7(.A(I0[10]), .B(n_275), .CI(\idtr[10] ), .Z(O0[10]), .CO(n_277
		));
	notech_fa2 i_6(.A(I0[9]), .B(n_273), .CI(\idtr[9] ), .Z(O0[9]), .CO(n_275
		));
	notech_fa2 i_5(.A(I0[8]), .B(n_271), .CI(\idtr[8] ), .Z(O0[8]), .CO(n_273
		));
	notech_fa2 i_4(.A(I0[7]), .B(n_269), .CI(\idtr[7] ), .Z(O0[7]), .CO(n_271
		));
	notech_fa2 i_3(.A(I0[6]), .B(n_267), .CI(\idtr[6] ), .Z(O0[6]), .CO(n_269
		));
	notech_fa2 i_2(.A(I0[5]), .B(n_265), .CI(\idtr[5] ), .Z(O0[5]), .CO(n_267
		));
	notech_fa2 i_1(.A(I0[4]), .B(n_322), .CI(\idtr[4] ), .Z(O0[4]), .CO(n_265
		));
	notech_ha2 i_0(.A(\idtr[3] ), .B(I0[3]), .Z(O0[3]), .CO(n_322));
endmodule
module AWDP_ADD_123(O0, opb, I0);

	output [32:0] O0;
	input [31:0] opb;
	input [31:0] I0;




	notech_inv i_10180(.A(n_58066), .Z(n_58071));
	notech_inv i_10176(.A(n_58066), .Z(n_58067));
	notech_inv i_10175(.A(I0[18]), .Z(n_58066));
	notech_fa2 i_31(.A(n_58071), .B(n_354), .CI(opb[31]), .Z(O0[31]), .CO(O0
		[32]));
	notech_fa2 i_30(.A(n_58071), .B(n_352), .CI(opb[30]), .Z(O0[30]), .CO(n_354
		));
	notech_fa2 i_29(.A(n_58071), .B(n_350), .CI(opb[29]), .Z(O0[29]), .CO(n_352
		));
	notech_fa2 i_28(.A(n_58071), .B(n_348), .CI(opb[28]), .Z(O0[28]), .CO(n_350
		));
	notech_fa2 i_27(.A(n_58071), .B(n_346), .CI(opb[27]), .Z(O0[27]), .CO(n_348
		));
	notech_fa2 i_26(.A(n_58071), .B(n_344), .CI(opb[26]), .Z(O0[26]), .CO(n_346
		));
	notech_fa2 i_25(.A(n_58071), .B(n_342), .CI(opb[25]), .Z(O0[25]), .CO(n_344
		));
	notech_fa2 i_24(.A(n_58071), .B(n_340), .CI(opb[24]), .Z(O0[24]), .CO(n_342
		));
	notech_fa2 i_23(.A(n_58071), .B(n_338), .CI(opb[23]), .Z(O0[23]), .CO(n_340
		));
	notech_fa2 i_22(.A(n_58071), .B(n_336), .CI(opb[22]), .Z(O0[22]), .CO(n_338
		));
	notech_fa2 i_21(.A(n_58071), .B(n_334), .CI(opb[21]), .Z(O0[21]), .CO(n_336
		));
	notech_fa2 i_20(.A(n_58071), .B(n_332), .CI(opb[20]), .Z(O0[20]), .CO(n_334
		));
	notech_fa2 i_19(.A(n_58071), .B(n_330), .CI(opb[19]), .Z(O0[19]), .CO(n_332
		));
	notech_fa2 i_18(.A(n_58071), .B(n_328), .CI(opb[18]), .Z(O0[18]), .CO(n_330
		));
	notech_fa2 i_17(.A(n_58071), .B(n_326), .CI(opb[17]), .Z(O0[17]), .CO(n_328
		));
	notech_fa2 i_16(.A(n_58067), .B(n_324), .CI(opb[16]), .Z(O0[16]), .CO(n_326
		));
	notech_fa2 i_15(.A(n_58067), .B(n_322), .CI(opb[15]), .Z(O0[15]), .CO(n_324
		));
	notech_fa2 i_14(.A(n_58067), .B(n_320), .CI(opb[14]), .Z(O0[14]), .CO(n_322
		));
	notech_fa2 i_13(.A(n_58067), .B(n_318), .CI(opb[13]), .Z(O0[13]), .CO(n_320
		));
	notech_fa2 i_12(.A(n_58067), .B(n_316), .CI(opb[12]), .Z(O0[12]), .CO(n_318
		));
	notech_fa2 i_11(.A(n_58067), .B(n_314), .CI(opb[11]), .Z(O0[11]), .CO(n_316
		));
	notech_fa2 i_10(.A(n_58067), .B(n_312), .CI(opb[10]), .Z(O0[10]), .CO(n_314
		));
	notech_fa2 i_9(.A(n_58067), .B(n_310), .CI(opb[9]), .Z(O0[9]), .CO(n_312
		));
	notech_fa2 i_8(.A(n_58071), .B(n_308), .CI(opb[8]), .Z(O0[8]), .CO(n_310
		));
	notech_fa2 i_7(.A(n_58071), .B(n_306), .CI(opb[7]), .Z(O0[7]), .CO(n_308
		));
	notech_fa2 i_6(.A(n_58071), .B(n_304), .CI(opb[6]), .Z(O0[6]), .CO(n_306
		));
	notech_fa2 i_5(.A(n_58071), .B(n_302), .CI(opb[5]), .Z(O0[5]), .CO(n_304
		));
	notech_fa2 i_4(.A(n_58067), .B(n_300), .CI(opb[4]), .Z(O0[4]), .CO(n_302
		));
	notech_fa2 i_3(.A(n_58067), .B(n_298), .CI(opb[3]), .Z(O0[3]), .CO(n_300
		));
	notech_fa2 i_2(.A(n_58071), .B(n_296), .CI(opb[2]), .Z(O0[2]), .CO(n_298
		));
	notech_fa2 i_1(.A(I0[1]), .B(n_361), .CI(opb[1]), .Z(O0[1]), .CO(n_296)
		);
	notech_ha2 i_0(.A(opb[0]), .B(I0[0]), .Z(O0[0]), .CO(n_361));
endmodule
module AWDP_ADD_135(O0, gdtr, I0);

	output [31:0] O0;
	input [31:0] gdtr;
	input [15:0] I0;

	wire \gdtr[1] ;
	wire \gdtr[2] ;
	wire \gdtr[3] ;
	wire \gdtr[4] ;
	wire \gdtr[5] ;
	wire \gdtr[6] ;
	wire \gdtr[7] ;
	wire \gdtr[8] ;
	wire \gdtr[9] ;
	wire \gdtr[10] ;
	wire \gdtr[11] ;
	wire \gdtr[12] ;
	wire \gdtr[13] ;
	wire \gdtr[14] ;
	wire \gdtr[15] ;
	wire \gdtr[16] ;
	wire \gdtr[17] ;
	wire \gdtr[18] ;
	wire \gdtr[19] ;
	wire \gdtr[20] ;
	wire \gdtr[21] ;
	wire \gdtr[22] ;
	wire \gdtr[23] ;
	wire \gdtr[24] ;
	wire \gdtr[25] ;
	wire \gdtr[26] ;
	wire \gdtr[27] ;
	wire \gdtr[28] ;
	wire \gdtr[29] ;
	wire \gdtr[30] ;
	wire \gdtr[31] ;


	assign O0[0] = gdtr[0];
	assign \gdtr[1]  = gdtr[1];
	assign \gdtr[2]  = gdtr[2];
	assign \gdtr[3]  = gdtr[3];
	assign \gdtr[4]  = gdtr[4];
	assign \gdtr[5]  = gdtr[5];
	assign \gdtr[6]  = gdtr[6];
	assign \gdtr[7]  = gdtr[7];
	assign \gdtr[8]  = gdtr[8];
	assign \gdtr[9]  = gdtr[9];
	assign \gdtr[10]  = gdtr[10];
	assign \gdtr[11]  = gdtr[11];
	assign \gdtr[12]  = gdtr[12];
	assign \gdtr[13]  = gdtr[13];
	assign \gdtr[14]  = gdtr[14];
	assign \gdtr[15]  = gdtr[15];
	assign \gdtr[16]  = gdtr[16];
	assign \gdtr[17]  = gdtr[17];
	assign \gdtr[18]  = gdtr[18];
	assign \gdtr[19]  = gdtr[19];
	assign \gdtr[20]  = gdtr[20];
	assign \gdtr[21]  = gdtr[21];
	assign \gdtr[22]  = gdtr[22];
	assign \gdtr[23]  = gdtr[23];
	assign \gdtr[24]  = gdtr[24];
	assign \gdtr[25]  = gdtr[25];
	assign \gdtr[26]  = gdtr[26];
	assign \gdtr[27]  = gdtr[27];
	assign \gdtr[28]  = gdtr[28];
	assign \gdtr[29]  = gdtr[29];
	assign \gdtr[30]  = gdtr[30];
	assign \gdtr[31]  = gdtr[31];

	notech_ha2 i_30(.A(\gdtr[31] ), .B(n_352), .Z(O0[31]));
	notech_ha2 i_29(.A(\gdtr[30] ), .B(n_350), .Z(O0[30]), .CO(n_352));
	notech_ha2 i_28(.A(\gdtr[29] ), .B(n_348), .Z(O0[29]), .CO(n_350));
	notech_ha2 i_27(.A(\gdtr[28] ), .B(n_346), .Z(O0[28]), .CO(n_348));
	notech_ha2 i_26(.A(\gdtr[27] ), .B(n_344), .Z(O0[27]), .CO(n_346));
	notech_ha2 i_25(.A(\gdtr[26] ), .B(n_342), .Z(O0[26]), .CO(n_344));
	notech_ha2 i_24(.A(\gdtr[25] ), .B(n_340), .Z(O0[25]), .CO(n_342));
	notech_ha2 i_23(.A(\gdtr[24] ), .B(n_338), .Z(O0[24]), .CO(n_340));
	notech_ha2 i_22(.A(\gdtr[23] ), .B(n_336), .Z(O0[23]), .CO(n_338));
	notech_ha2 i_21(.A(\gdtr[22] ), .B(n_334), .Z(O0[22]), .CO(n_336));
	notech_ha2 i_20(.A(\gdtr[21] ), .B(n_332), .Z(O0[21]), .CO(n_334));
	notech_ha2 i_19(.A(\gdtr[20] ), .B(n_330), .Z(O0[20]), .CO(n_332));
	notech_ha2 i_18(.A(\gdtr[19] ), .B(n_328), .Z(O0[19]), .CO(n_330));
	notech_ha2 i_17(.A(\gdtr[18] ), .B(n_326), .Z(O0[18]), .CO(n_328));
	notech_ha2 i_16(.A(\gdtr[17] ), .B(n_324), .Z(O0[17]), .CO(n_326));
	notech_ha2 i_15(.A(\gdtr[16] ), .B(n_285), .Z(O0[16]), .CO(n_324));
	notech_fa2 i_14(.A(I0[15]), .B(n_283), .CI(\gdtr[15] ), .Z(O0[15]), .CO(n_285
		));
	notech_fa2 i_13(.A(I0[14]), .B(n_281), .CI(\gdtr[14] ), .Z(O0[14]), .CO(n_283
		));
	notech_fa2 i_12(.A(I0[13]), .B(n_279), .CI(\gdtr[13] ), .Z(O0[13]), .CO(n_281
		));
	notech_fa2 i_11(.A(I0[12]), .B(n_277), .CI(\gdtr[12] ), .Z(O0[12]), .CO(n_279
		));
	notech_fa2 i_10(.A(I0[11]), .B(n_275), .CI(\gdtr[11] ), .Z(O0[11]), .CO(n_277
		));
	notech_fa2 i_9(.A(I0[10]), .B(n_273), .CI(\gdtr[10] ), .Z(O0[10]), .CO(n_275
		));
	notech_fa2 i_8(.A(I0[9]), .B(n_271), .CI(\gdtr[9] ), .Z(O0[9]), .CO(n_273
		));
	notech_fa2 i_7(.A(I0[8]), .B(n_269), .CI(\gdtr[8] ), .Z(O0[8]), .CO(n_271
		));
	notech_fa2 i_6(.A(I0[7]), .B(n_267), .CI(\gdtr[7] ), .Z(O0[7]), .CO(n_269
		));
	notech_fa2 i_5(.A(I0[6]), .B(n_265), .CI(\gdtr[6] ), .Z(O0[6]), .CO(n_267
		));
	notech_fa2 i_4(.A(I0[5]), .B(n_263), .CI(\gdtr[5] ), .Z(O0[5]), .CO(n_265
		));
	notech_fa2 i_3(.A(I0[4]), .B(n_261), .CI(\gdtr[4] ), .Z(O0[4]), .CO(n_263
		));
	notech_fa2 i_2(.A(I0[3]), .B(n_322), .CI(\gdtr[3] ), .Z(O0[3]), .CO(n_261
		));
	notech_ha2 i_1(.A(\gdtr[2] ), .B(\gdtr[1] ), .Z(O0[2]), .CO(n_322));
	notech_inv i_0(.A(\gdtr[1] ), .Z(O0[1]));
endmodule
module AWDP_ADD_160(O0, opb, I0);

	output [16:0] O0;
	input [15:0] opb;
	input [15:0] I0;




	notech_fa2 i_15(.A(I0[15]), .B(n_178), .CI(opb[15]), .Z(O0[15]), .CO(O0[
		16]));
	notech_fa2 i_14(.A(I0[15]), .B(n_176), .CI(opb[14]), .Z(O0[14]), .CO(n_178
		));
	notech_fa2 i_13(.A(I0[15]), .B(n_174), .CI(opb[13]), .Z(O0[13]), .CO(n_176
		));
	notech_fa2 i_12(.A(I0[15]), .B(n_172), .CI(opb[12]), .Z(O0[12]), .CO(n_174
		));
	notech_fa2 i_11(.A(I0[15]), .B(n_170), .CI(opb[11]), .Z(O0[11]), .CO(n_172
		));
	notech_fa2 i_10(.A(I0[15]), .B(n_168), .CI(opb[10]), .Z(O0[10]), .CO(n_170
		));
	notech_fa2 i_9(.A(I0[15]), .B(n_166), .CI(opb[9]), .Z(O0[9]), .CO(n_168)
		);
	notech_fa2 i_8(.A(I0[15]), .B(n_164), .CI(opb[8]), .Z(O0[8]), .CO(n_166)
		);
	notech_fa2 i_7(.A(I0[15]), .B(n_162), .CI(opb[7]), .Z(O0[7]), .CO(n_164)
		);
	notech_fa2 i_6(.A(I0[15]), .B(n_160), .CI(opb[6]), .Z(O0[6]), .CO(n_162)
		);
	notech_fa2 i_5(.A(I0[15]), .B(n_158), .CI(opb[5]), .Z(O0[5]), .CO(n_160)
		);
	notech_fa2 i_4(.A(I0[15]), .B(n_156), .CI(opb[4]), .Z(O0[4]), .CO(n_158)
		);
	notech_fa2 i_3(.A(I0[15]), .B(n_154), .CI(opb[3]), .Z(O0[3]), .CO(n_156)
		);
	notech_fa2 i_2(.A(I0[15]), .B(n_152), .CI(opb[2]), .Z(O0[2]), .CO(n_154)
		);
	notech_fa2 i_1(.A(I0[1]), .B(n_185), .CI(opb[1]), .Z(O0[1]), .CO(n_152)
		);
	notech_ha2 i_0(.A(opb[0]), .B(I0[0]), .Z(O0[0]), .CO(n_185));
endmodule
module AWDP_ADD_177(O0, opa, I0);

	output [32:0] O0;
	input [31:0] opa;
	input [31:0] I0;




	notech_inv i_10202(.A(n_58162), .Z(n_58167));
	notech_inv i_10198(.A(n_58162), .Z(n_58163));
	notech_inv i_10197(.A(I0[19]), .Z(n_58162));
	notech_fa2 i_31(.A(n_58167), .B(n_354), .CI(opa[31]), .Z(O0[31]), .CO(O0
		[32]));
	notech_fa2 i_30(.A(n_58167), .B(n_352), .CI(opa[30]), .Z(O0[30]), .CO(n_354
		));
	notech_fa2 i_29(.A(n_58167), .B(n_350), .CI(opa[29]), .Z(O0[29]), .CO(n_352
		));
	notech_fa2 i_28(.A(n_58167), .B(n_348), .CI(opa[28]), .Z(O0[28]), .CO(n_350
		));
	notech_fa2 i_27(.A(n_58167), .B(n_346), .CI(opa[27]), .Z(O0[27]), .CO(n_348
		));
	notech_fa2 i_26(.A(n_58167), .B(n_344), .CI(opa[26]), .Z(O0[26]), .CO(n_346
		));
	notech_fa2 i_25(.A(n_58167), .B(n_342), .CI(opa[25]), .Z(O0[25]), .CO(n_344
		));
	notech_fa2 i_24(.A(n_58167), .B(n_340), .CI(opa[24]), .Z(O0[24]), .CO(n_342
		));
	notech_fa2 i_23(.A(n_58167), .B(n_338), .CI(opa[23]), .Z(O0[23]), .CO(n_340
		));
	notech_fa2 i_22(.A(n_58167), .B(n_336), .CI(opa[22]), .Z(O0[22]), .CO(n_338
		));
	notech_fa2 i_21(.A(n_58167), .B(n_334), .CI(opa[21]), .Z(O0[21]), .CO(n_336
		));
	notech_fa2 i_20(.A(n_58167), .B(n_332), .CI(opa[20]), .Z(O0[20]), .CO(n_334
		));
	notech_fa2 i_19(.A(n_58167), .B(n_330), .CI(opa[19]), .Z(O0[19]), .CO(n_332
		));
	notech_fa2 i_18(.A(n_58167), .B(n_328), .CI(opa[18]), .Z(O0[18]), .CO(n_330
		));
	notech_fa2 i_17(.A(n_58167), .B(n_326), .CI(opa[17]), .Z(O0[17]), .CO(n_328
		));
	notech_fa2 i_16(.A(n_58163), .B(n_324), .CI(opa[16]), .Z(O0[16]), .CO(n_326
		));
	notech_fa2 i_15(.A(n_58163), .B(n_322), .CI(opa[15]), .Z(O0[15]), .CO(n_324
		));
	notech_fa2 i_14(.A(n_58163), .B(n_320), .CI(opa[14]), .Z(O0[14]), .CO(n_322
		));
	notech_fa2 i_13(.A(n_58163), .B(n_318), .CI(opa[13]), .Z(O0[13]), .CO(n_320
		));
	notech_fa2 i_12(.A(n_58163), .B(n_316), .CI(opa[12]), .Z(O0[12]), .CO(n_318
		));
	notech_fa2 i_11(.A(n_58163), .B(n_314), .CI(opa[11]), .Z(O0[11]), .CO(n_316
		));
	notech_fa2 i_10(.A(n_58163), .B(n_312), .CI(opa[10]), .Z(O0[10]), .CO(n_314
		));
	notech_fa2 i_9(.A(n_58163), .B(n_310), .CI(opa[9]), .Z(O0[9]), .CO(n_312
		));
	notech_fa2 i_8(.A(n_58167), .B(n_308), .CI(opa[8]), .Z(O0[8]), .CO(n_310
		));
	notech_fa2 i_7(.A(n_58167), .B(n_306), .CI(opa[7]), .Z(O0[7]), .CO(n_308
		));
	notech_fa2 i_6(.A(n_58167), .B(n_304), .CI(opa[6]), .Z(O0[6]), .CO(n_306
		));
	notech_fa2 i_5(.A(n_58167), .B(n_302), .CI(opa[5]), .Z(O0[5]), .CO(n_304
		));
	notech_fa2 i_4(.A(n_58163), .B(n_300), .CI(opa[4]), .Z(O0[4]), .CO(n_302
		));
	notech_fa2 i_3(.A(n_58163), .B(n_298), .CI(opa[3]), .Z(O0[3]), .CO(n_300
		));
	notech_fa2 i_2(.A(n_58167), .B(n_296), .CI(opa[2]), .Z(O0[2]), .CO(n_298
		));
	notech_fa2 i_1(.A(I0[1]), .B(n_361), .CI(opa[1]), .Z(O0[1]), .CO(n_296)
		);
	notech_ha2 i_0(.A(opa[0]), .B(I0[0]), .Z(O0[0]), .CO(n_361));
endmodule
module AWDP_ADD_189(O0, opd);

	output [31:0] O0;
	input [31:0] opd;

	wire \opd[2] ;
	wire \opd[3] ;
	wire \opd[4] ;
	wire \opd[5] ;
	wire \opd[6] ;
	wire \opd[7] ;
	wire \opd[8] ;
	wire \opd[9] ;
	wire \opd[10] ;
	wire \opd[11] ;
	wire \opd[12] ;
	wire \opd[13] ;
	wire \opd[14] ;
	wire \opd[15] ;
	wire \opd[16] ;
	wire \opd[17] ;
	wire \opd[18] ;
	wire \opd[19] ;
	wire \opd[20] ;
	wire \opd[21] ;
	wire \opd[22] ;
	wire \opd[23] ;
	wire \opd[24] ;
	wire \opd[25] ;
	wire \opd[26] ;
	wire \opd[27] ;
	wire \opd[28] ;
	wire \opd[29] ;
	wire \opd[30] ;
	wire \opd[31] ;


	assign O0[0] = opd[0];
	assign O0[1] = opd[1];
	assign \opd[2]  = opd[2];
	assign \opd[3]  = opd[3];
	assign \opd[4]  = opd[4];
	assign \opd[5]  = opd[5];
	assign \opd[6]  = opd[6];
	assign \opd[7]  = opd[7];
	assign \opd[8]  = opd[8];
	assign \opd[9]  = opd[9];
	assign \opd[10]  = opd[10];
	assign \opd[11]  = opd[11];
	assign \opd[12]  = opd[12];
	assign \opd[13]  = opd[13];
	assign \opd[14]  = opd[14];
	assign \opd[15]  = opd[15];
	assign \opd[16]  = opd[16];
	assign \opd[17]  = opd[17];
	assign \opd[18]  = opd[18];
	assign \opd[19]  = opd[19];
	assign \opd[20]  = opd[20];
	assign \opd[21]  = opd[21];
	assign \opd[22]  = opd[22];
	assign \opd[23]  = opd[23];
	assign \opd[24]  = opd[24];
	assign \opd[25]  = opd[25];
	assign \opd[26]  = opd[26];
	assign \opd[27]  = opd[27];
	assign \opd[28]  = opd[28];
	assign \opd[29]  = opd[29];
	assign \opd[30]  = opd[30];
	assign \opd[31]  = opd[31];

	notech_ha2 i_29(.A(\opd[31] ), .B(n_308), .Z(O0[31]));
	notech_ha2 i_28(.A(\opd[30] ), .B(n_306), .Z(O0[30]), .CO(n_308));
	notech_ha2 i_27(.A(\opd[29] ), .B(n_304), .Z(O0[29]), .CO(n_306));
	notech_ha2 i_26(.A(\opd[28] ), .B(n_302), .Z(O0[28]), .CO(n_304));
	notech_ha2 i_25(.A(\opd[27] ), .B(n_300), .Z(O0[27]), .CO(n_302));
	notech_ha2 i_24(.A(\opd[26] ), .B(n_298), .Z(O0[26]), .CO(n_300));
	notech_ha2 i_23(.A(\opd[25] ), .B(n_296), .Z(O0[25]), .CO(n_298));
	notech_ha2 i_22(.A(\opd[24] ), .B(n_294), .Z(O0[24]), .CO(n_296));
	notech_ha2 i_21(.A(\opd[23] ), .B(n_292), .Z(O0[23]), .CO(n_294));
	notech_ha2 i_20(.A(\opd[22] ), .B(n_290), .Z(O0[22]), .CO(n_292));
	notech_ha2 i_19(.A(\opd[21] ), .B(n_288), .Z(O0[21]), .CO(n_290));
	notech_ha2 i_18(.A(\opd[20] ), .B(n_286), .Z(O0[20]), .CO(n_288));
	notech_ha2 i_17(.A(\opd[19] ), .B(n_284), .Z(O0[19]), .CO(n_286));
	notech_ha2 i_16(.A(\opd[18] ), .B(n_282), .Z(O0[18]), .CO(n_284));
	notech_ha2 i_15(.A(\opd[17] ), .B(n_280), .Z(O0[17]), .CO(n_282));
	notech_ha2 i_14(.A(\opd[16] ), .B(n_278), .Z(O0[16]), .CO(n_280));
	notech_ha2 i_13(.A(\opd[15] ), .B(n_276), .Z(O0[15]), .CO(n_278));
	notech_ha2 i_12(.A(\opd[14] ), .B(n_274), .Z(O0[14]), .CO(n_276));
	notech_ha2 i_11(.A(\opd[13] ), .B(n_272), .Z(O0[13]), .CO(n_274));
	notech_ha2 i_10(.A(\opd[12] ), .B(n_270), .Z(O0[12]), .CO(n_272));
	notech_ha2 i_9(.A(\opd[11] ), .B(n_268), .Z(O0[11]), .CO(n_270));
	notech_ha2 i_8(.A(\opd[10] ), .B(n_266), .Z(O0[10]), .CO(n_268));
	notech_ha2 i_7(.A(\opd[9] ), .B(n_264), .Z(O0[9]), .CO(n_266));
	notech_ha2 i_6(.A(\opd[8] ), .B(n_262), .Z(O0[8]), .CO(n_264));
	notech_ha2 i_5(.A(\opd[7] ), .B(n_260), .Z(O0[7]), .CO(n_262));
	notech_ha2 i_4(.A(\opd[6] ), .B(n_258), .Z(O0[6]), .CO(n_260));
	notech_ha2 i_3(.A(\opd[5] ), .B(n_256), .Z(O0[5]), .CO(n_258));
	notech_ha2 i_2(.A(\opd[4] ), .B(n_254), .Z(O0[4]), .CO(n_256));
	notech_ha2 i_1(.A(\opd[3] ), .B(\opd[2] ), .Z(O0[3]), .CO(n_254));
	notech_inv i_0(.A(\opd[2] ), .Z(O0[2]));
endmodule
module AWDP_ADD_190(O0, I0, I1);

	output [31:0] O0;
	input [31:0] I0;
	input [31:0] I1;

	wire \I0[4] ;
	wire \I0[5] ;
	wire \I0[6] ;
	wire \I0[7] ;
	wire \I0[8] ;
	wire \I0[9] ;
	wire \I0[10] ;
	wire \I0[11] ;
	wire \I0[12] ;
	wire \I0[13] ;
	wire \I0[14] ;
	wire \I0[15] ;


	assign O0[0] = I0[0];
	assign O0[1] = I0[1];
	assign O0[2] = I0[2];
	assign O0[3] = I0[3];
	assign \I0[4]  = I0[4];
	assign \I0[5]  = I0[5];
	assign \I0[6]  = I0[6];
	assign \I0[7]  = I0[7];
	assign \I0[8]  = I0[8];
	assign \I0[9]  = I0[9];
	assign \I0[10]  = I0[10];
	assign \I0[11]  = I0[11];
	assign \I0[12]  = I0[12];
	assign \I0[13]  = I0[13];
	assign \I0[14]  = I0[14];
	assign \I0[15]  = I0[15];

	notech_ha2 i_27(.A(I1[31]), .B(n_376), .Z(O0[31]));
	notech_ha2 i_26(.A(I1[30]), .B(n_374), .Z(O0[30]), .CO(n_376));
	notech_ha2 i_25(.A(I1[29]), .B(n_372), .Z(O0[29]), .CO(n_374));
	notech_ha2 i_24(.A(I1[28]), .B(n_370), .Z(O0[28]), .CO(n_372));
	notech_ha2 i_23(.A(I1[27]), .B(n_368), .Z(O0[27]), .CO(n_370));
	notech_ha2 i_22(.A(I1[26]), .B(n_366), .Z(O0[26]), .CO(n_368));
	notech_ha2 i_21(.A(I1[25]), .B(n_364), .Z(O0[25]), .CO(n_366));
	notech_ha2 i_20(.A(I1[24]), .B(n_362), .Z(O0[24]), .CO(n_364));
	notech_ha2 i_19(.A(I1[23]), .B(n_360), .Z(O0[23]), .CO(n_362));
	notech_ha2 i_18(.A(I1[22]), .B(n_358), .Z(O0[22]), .CO(n_360));
	notech_ha2 i_17(.A(I1[21]), .B(n_356), .Z(O0[21]), .CO(n_358));
	notech_ha2 i_16(.A(I1[20]), .B(n_354), .Z(O0[20]), .CO(n_356));
	notech_ha2 i_15(.A(I1[19]), .B(n_352), .Z(O0[19]), .CO(n_354));
	notech_ha2 i_14(.A(I1[18]), .B(n_350), .Z(O0[18]), .CO(n_352));
	notech_ha2 i_13(.A(I1[17]), .B(n_348), .Z(O0[17]), .CO(n_350));
	notech_ha2 i_12(.A(I1[16]), .B(n_311), .Z(O0[16]), .CO(n_348));
	notech_fa2 i_11(.A(\I0[15] ), .B(n_309), .CI(I1[15]), .Z(O0[15]), .CO(n_311
		));
	notech_fa2 i_10(.A(\I0[14] ), .B(n_307), .CI(I1[14]), .Z(O0[14]), .CO(n_309
		));
	notech_fa2 i_9(.A(\I0[13] ), .B(n_305), .CI(I1[13]), .Z(O0[13]), .CO(n_307
		));
	notech_fa2 i_8(.A(\I0[12] ), .B(n_303), .CI(I1[12]), .Z(O0[12]), .CO(n_305
		));
	notech_fa2 i_7(.A(\I0[11] ), .B(n_301), .CI(I1[11]), .Z(O0[11]), .CO(n_303
		));
	notech_fa2 i_6(.A(\I0[10] ), .B(n_299), .CI(I1[10]), .Z(O0[10]), .CO(n_301
		));
	notech_fa2 i_5(.A(\I0[9] ), .B(n_297), .CI(I1[9]), .Z(O0[9]), .CO(n_299)
		);
	notech_fa2 i_4(.A(\I0[8] ), .B(n_295), .CI(I1[8]), .Z(O0[8]), .CO(n_297)
		);
	notech_fa2 i_3(.A(\I0[7] ), .B(n_293), .CI(I1[7]), .Z(O0[7]), .CO(n_295)
		);
	notech_fa2 i_2(.A(\I0[6] ), .B(n_291), .CI(I1[6]), .Z(O0[6]), .CO(n_293)
		);
	notech_fa2 i_1(.A(\I0[5] ), .B(n_346), .CI(I1[5]), .Z(O0[5]), .CO(n_291)
		);
	notech_ha2 i_0(.A(\I0[4] ), .B(I1[4]), .Z(O0[4]), .CO(n_346));
endmodule
module AWDP_ADD_198(O0, opd, I0);

	output [32:0] O0;
	input [31:0] opd;
	input [31:0] I0;




	notech_inv i_10168(.A(n_58028), .Z(n_58029));
	notech_inv i_10167(.A(I0[4]), .Z(n_58028));
	notech_fa2 i_31(.A(I0[4]), .B(n_354), .CI(opd[31]), .Z(O0[31]), .CO(O0[
		32]));
	notech_fa2 i_30(.A(I0[4]), .B(n_352), .CI(opd[30]), .Z(O0[30]), .CO(n_354
		));
	notech_fa2 i_29(.A(I0[4]), .B(n_350), .CI(opd[29]), .Z(O0[29]), .CO(n_352
		));
	notech_fa2 i_28(.A(I0[4]), .B(n_348), .CI(opd[28]), .Z(O0[28]), .CO(n_350
		));
	notech_fa2 i_27(.A(I0[4]), .B(n_346), .CI(opd[27]), .Z(O0[27]), .CO(n_348
		));
	notech_fa2 i_26(.A(I0[4]), .B(n_344), .CI(opd[26]), .Z(O0[26]), .CO(n_346
		));
	notech_fa2 i_25(.A(I0[4]), .B(n_342), .CI(opd[25]), .Z(O0[25]), .CO(n_344
		));
	notech_fa2 i_24(.A(I0[4]), .B(n_340), .CI(opd[24]), .Z(O0[24]), .CO(n_342
		));
	notech_fa2 i_23(.A(I0[4]), .B(n_338), .CI(opd[23]), .Z(O0[23]), .CO(n_340
		));
	notech_fa2 i_22(.A(I0[4]), .B(n_336), .CI(opd[22]), .Z(O0[22]), .CO(n_338
		));
	notech_fa2 i_21(.A(I0[4]), .B(n_334), .CI(opd[21]), .Z(O0[21]), .CO(n_336
		));
	notech_fa2 i_20(.A(I0[4]), .B(n_332), .CI(opd[20]), .Z(O0[20]), .CO(n_334
		));
	notech_fa2 i_19(.A(I0[4]), .B(n_330), .CI(opd[19]), .Z(O0[19]), .CO(n_332
		));
	notech_fa2 i_18(.A(I0[4]), .B(n_328), .CI(opd[18]), .Z(O0[18]), .CO(n_330
		));
	notech_fa2 i_17(.A(I0[4]), .B(n_326), .CI(opd[17]), .Z(O0[17]), .CO(n_328
		));
	notech_fa2 i_16(.A(n_58029), .B(n_324), .CI(opd[16]), .Z(O0[16]), .CO(n_326
		));
	notech_fa2 i_15(.A(n_58029), .B(n_322), .CI(opd[15]), .Z(O0[15]), .CO(n_324
		));
	notech_fa2 i_14(.A(n_58029), .B(n_320), .CI(opd[14]), .Z(O0[14]), .CO(n_322
		));
	notech_fa2 i_13(.A(n_58029), .B(n_318), .CI(opd[13]), .Z(O0[13]), .CO(n_320
		));
	notech_fa2 i_12(.A(n_58029), .B(n_316), .CI(opd[12]), .Z(O0[12]), .CO(n_318
		));
	notech_fa2 i_11(.A(n_58029), .B(n_314), .CI(opd[11]), .Z(O0[11]), .CO(n_316
		));
	notech_fa2 i_10(.A(n_58029), .B(n_312), .CI(opd[10]), .Z(O0[10]), .CO(n_314
		));
	notech_fa2 i_9(.A(n_58029), .B(n_310), .CI(opd[9]), .Z(O0[9]), .CO(n_312
		));
	notech_fa2 i_8(.A(n_58029), .B(n_308), .CI(opd[8]), .Z(O0[8]), .CO(n_310
		));
	notech_fa2 i_7(.A(n_58029), .B(n_306), .CI(opd[7]), .Z(O0[7]), .CO(n_308
		));
	notech_fa2 i_6(.A(n_58029), .B(n_304), .CI(opd[6]), .Z(O0[6]), .CO(n_306
		));
	notech_fa2 i_5(.A(n_58029), .B(n_302), .CI(opd[5]), .Z(O0[5]), .CO(n_304
		));
	notech_fa2 i_4(.A(n_58029), .B(n_300), .CI(opd[4]), .Z(O0[4]), .CO(n_302
		));
	notech_fa2 i_3(.A(n_58029), .B(n_298), .CI(opd[3]), .Z(O0[3]), .CO(n_300
		));
	notech_fa2 i_2(.A(n_58029), .B(n_296), .CI(opd[2]), .Z(O0[2]), .CO(n_298
		));
	notech_fa2 i_1(.A(I0[1]), .B(n_361), .CI(opd[1]), .Z(O0[1]), .CO(n_296)
		);
	notech_ha2 i_0(.A(opd[0]), .B(I0[0]), .Z(O0[0]), .CO(n_361));
endmodule
module AWDP_ADD_20(O0, opd, desc);
    output [31:0] O0;
    input [31:0] opd;
    input [31:0] desc;
    // Line 1146
    wire [31:0] N205;
    // Line 1144
    wire [31:0] O0;

    // Line 1146
    assign N205 = desc + opd;
    // Line 1144
    assign O0 = N205;
endmodule

module AWDP_ADD_201(O0, ldtr, I0);

	output [31:0] O0;
	input [31:0] ldtr;
	input [31:0] I0;

	wire \ldtr[1] ;
	wire \ldtr[2] ;
	wire \ldtr[3] ;
	wire \ldtr[4] ;
	wire \ldtr[5] ;
	wire \ldtr[6] ;
	wire \ldtr[7] ;
	wire \ldtr[8] ;
	wire \ldtr[9] ;
	wire \ldtr[10] ;
	wire \ldtr[11] ;
	wire \ldtr[12] ;
	wire \ldtr[13] ;
	wire \ldtr[14] ;
	wire \ldtr[15] ;
	wire \ldtr[16] ;
	wire \ldtr[17] ;
	wire \ldtr[18] ;
	wire \ldtr[19] ;
	wire \ldtr[20] ;
	wire \ldtr[21] ;
	wire \ldtr[22] ;
	wire \ldtr[23] ;
	wire \ldtr[24] ;
	wire \ldtr[25] ;
	wire \ldtr[26] ;
	wire \ldtr[27] ;
	wire \ldtr[28] ;
	wire \ldtr[29] ;
	wire \ldtr[30] ;
	wire \ldtr[31] ;


	assign O0[0] = ldtr[0];
	assign \ldtr[1]  = ldtr[1];
	assign \ldtr[2]  = ldtr[2];
	assign \ldtr[3]  = ldtr[3];
	assign \ldtr[4]  = ldtr[4];
	assign \ldtr[5]  = ldtr[5];
	assign \ldtr[6]  = ldtr[6];
	assign \ldtr[7]  = ldtr[7];
	assign \ldtr[8]  = ldtr[8];
	assign \ldtr[9]  = ldtr[9];
	assign \ldtr[10]  = ldtr[10];
	assign \ldtr[11]  = ldtr[11];
	assign \ldtr[12]  = ldtr[12];
	assign \ldtr[13]  = ldtr[13];
	assign \ldtr[14]  = ldtr[14];
	assign \ldtr[15]  = ldtr[15];
	assign \ldtr[16]  = ldtr[16];
	assign \ldtr[17]  = ldtr[17];
	assign \ldtr[18]  = ldtr[18];
	assign \ldtr[19]  = ldtr[19];
	assign \ldtr[20]  = ldtr[20];
	assign \ldtr[21]  = ldtr[21];
	assign \ldtr[22]  = ldtr[22];
	assign \ldtr[23]  = ldtr[23];
	assign \ldtr[24]  = ldtr[24];
	assign \ldtr[25]  = ldtr[25];
	assign \ldtr[26]  = ldtr[26];
	assign \ldtr[27]  = ldtr[27];
	assign \ldtr[28]  = ldtr[28];
	assign \ldtr[29]  = ldtr[29];
	assign \ldtr[30]  = ldtr[30];
	assign \ldtr[31]  = ldtr[31];

	notech_fa2 i_30(.A(I0[31]), .B(n_347), .CI(\ldtr[31] ), .Z(O0[31]));
	notech_fa2 i_29(.A(I0[30]), .B(n_345), .CI(\ldtr[30] ), .Z(O0[30]), .CO(n_347
		));
	notech_fa2 i_28(.A(I0[29]), .B(n_343), .CI(\ldtr[29] ), .Z(O0[29]), .CO(n_345
		));
	notech_fa2 i_27(.A(I0[28]), .B(n_341), .CI(\ldtr[28] ), .Z(O0[28]), .CO(n_343
		));
	notech_fa2 i_26(.A(I0[27]), .B(n_339), .CI(\ldtr[27] ), .Z(O0[27]), .CO(n_341
		));
	notech_fa2 i_25(.A(I0[26]), .B(n_337), .CI(\ldtr[26] ), .Z(O0[26]), .CO(n_339
		));
	notech_fa2 i_24(.A(I0[25]), .B(n_335), .CI(\ldtr[25] ), .Z(O0[25]), .CO(n_337
		));
	notech_fa2 i_23(.A(I0[24]), .B(n_333), .CI(\ldtr[24] ), .Z(O0[24]), .CO(n_335
		));
	notech_fa2 i_22(.A(I0[23]), .B(n_331), .CI(\ldtr[23] ), .Z(O0[23]), .CO(n_333
		));
	notech_fa2 i_21(.A(I0[22]), .B(n_329), .CI(\ldtr[22] ), .Z(O0[22]), .CO(n_331
		));
	notech_fa2 i_20(.A(I0[21]), .B(n_327), .CI(\ldtr[21] ), .Z(O0[21]), .CO(n_329
		));
	notech_fa2 i_19(.A(I0[20]), .B(n_325), .CI(\ldtr[20] ), .Z(O0[20]), .CO(n_327
		));
	notech_fa2 i_18(.A(I0[19]), .B(n_323), .CI(\ldtr[19] ), .Z(O0[19]), .CO(n_325
		));
	notech_fa2 i_17(.A(I0[18]), .B(n_321), .CI(\ldtr[18] ), .Z(O0[18]), .CO(n_323
		));
	notech_fa2 i_16(.A(I0[17]), .B(n_319), .CI(\ldtr[17] ), .Z(O0[17]), .CO(n_321
		));
	notech_fa2 i_15(.A(I0[16]), .B(n_317), .CI(\ldtr[16] ), .Z(O0[16]), .CO(n_319
		));
	notech_fa2 i_14(.A(I0[15]), .B(n_315), .CI(\ldtr[15] ), .Z(O0[15]), .CO(n_317
		));
	notech_fa2 i_13(.A(I0[14]), .B(n_313), .CI(\ldtr[14] ), .Z(O0[14]), .CO(n_315
		));
	notech_fa2 i_12(.A(I0[13]), .B(n_311), .CI(\ldtr[13] ), .Z(O0[13]), .CO(n_313
		));
	notech_fa2 i_11(.A(I0[12]), .B(n_309), .CI(\ldtr[12] ), .Z(O0[12]), .CO(n_311
		));
	notech_fa2 i_10(.A(I0[11]), .B(n_307), .CI(\ldtr[11] ), .Z(O0[11]), .CO(n_309
		));
	notech_fa2 i_9(.A(I0[10]), .B(n_305), .CI(\ldtr[10] ), .Z(O0[10]), .CO(n_307
		));
	notech_fa2 i_8(.A(I0[9]), .B(n_303), .CI(\ldtr[9] ), .Z(O0[9]), .CO(n_305
		));
	notech_fa2 i_7(.A(I0[8]), .B(n_301), .CI(\ldtr[8] ), .Z(O0[8]), .CO(n_303
		));
	notech_fa2 i_6(.A(I0[7]), .B(n_299), .CI(\ldtr[7] ), .Z(O0[7]), .CO(n_301
		));
	notech_fa2 i_5(.A(I0[6]), .B(n_297), .CI(\ldtr[6] ), .Z(O0[6]), .CO(n_299
		));
	notech_fa2 i_4(.A(I0[5]), .B(n_295), .CI(\ldtr[5] ), .Z(O0[5]), .CO(n_297
		));
	notech_fa2 i_3(.A(I0[4]), .B(n_293), .CI(\ldtr[4] ), .Z(O0[4]), .CO(n_295
		));
	notech_fa2 i_2(.A(I0[3]), .B(n_354), .CI(\ldtr[3] ), .Z(O0[3]), .CO(n_293
		));
	notech_ha2 i_1(.A(\ldtr[2] ), .B(\ldtr[1] ), .Z(O0[2]), .CO(n_354));
	notech_inv i_0(.A(\ldtr[1] ), .Z(O0[1]));
endmodule
module AWDP_ADD_216(O0, gdtr, I0);

	output [31:0] O0;
	input [31:0] gdtr;
	input [31:0] I0;

	wire \gdtr[1] ;
	wire \gdtr[2] ;
	wire \gdtr[3] ;
	wire \gdtr[4] ;
	wire \gdtr[5] ;
	wire \gdtr[6] ;
	wire \gdtr[7] ;
	wire \gdtr[8] ;
	wire \gdtr[9] ;
	wire \gdtr[10] ;
	wire \gdtr[11] ;
	wire \gdtr[12] ;
	wire \gdtr[13] ;
	wire \gdtr[14] ;
	wire \gdtr[15] ;
	wire \gdtr[16] ;
	wire \gdtr[17] ;
	wire \gdtr[18] ;
	wire \gdtr[19] ;
	wire \gdtr[20] ;
	wire \gdtr[21] ;
	wire \gdtr[22] ;
	wire \gdtr[23] ;
	wire \gdtr[24] ;
	wire \gdtr[25] ;
	wire \gdtr[26] ;
	wire \gdtr[27] ;
	wire \gdtr[28] ;
	wire \gdtr[29] ;
	wire \gdtr[30] ;
	wire \gdtr[31] ;


	assign O0[0] = gdtr[0];
	assign \gdtr[1]  = gdtr[1];
	assign \gdtr[2]  = gdtr[2];
	assign \gdtr[3]  = gdtr[3];
	assign \gdtr[4]  = gdtr[4];
	assign \gdtr[5]  = gdtr[5];
	assign \gdtr[6]  = gdtr[6];
	assign \gdtr[7]  = gdtr[7];
	assign \gdtr[8]  = gdtr[8];
	assign \gdtr[9]  = gdtr[9];
	assign \gdtr[10]  = gdtr[10];
	assign \gdtr[11]  = gdtr[11];
	assign \gdtr[12]  = gdtr[12];
	assign \gdtr[13]  = gdtr[13];
	assign \gdtr[14]  = gdtr[14];
	assign \gdtr[15]  = gdtr[15];
	assign \gdtr[16]  = gdtr[16];
	assign \gdtr[17]  = gdtr[17];
	assign \gdtr[18]  = gdtr[18];
	assign \gdtr[19]  = gdtr[19];
	assign \gdtr[20]  = gdtr[20];
	assign \gdtr[21]  = gdtr[21];
	assign \gdtr[22]  = gdtr[22];
	assign \gdtr[23]  = gdtr[23];
	assign \gdtr[24]  = gdtr[24];
	assign \gdtr[25]  = gdtr[25];
	assign \gdtr[26]  = gdtr[26];
	assign \gdtr[27]  = gdtr[27];
	assign \gdtr[28]  = gdtr[28];
	assign \gdtr[29]  = gdtr[29];
	assign \gdtr[30]  = gdtr[30];
	assign \gdtr[31]  = gdtr[31];

	notech_fa2 i_30(.A(I0[31]), .B(n_347), .CI(\gdtr[31] ), .Z(O0[31]));
	notech_fa2 i_29(.A(I0[30]), .B(n_345), .CI(\gdtr[30] ), .Z(O0[30]), .CO(n_347
		));
	notech_fa2 i_28(.A(I0[29]), .B(n_343), .CI(\gdtr[29] ), .Z(O0[29]), .CO(n_345
		));
	notech_fa2 i_27(.A(I0[28]), .B(n_341), .CI(\gdtr[28] ), .Z(O0[28]), .CO(n_343
		));
	notech_fa2 i_26(.A(I0[27]), .B(n_339), .CI(\gdtr[27] ), .Z(O0[27]), .CO(n_341
		));
	notech_fa2 i_25(.A(I0[26]), .B(n_337), .CI(\gdtr[26] ), .Z(O0[26]), .CO(n_339
		));
	notech_fa2 i_24(.A(I0[25]), .B(n_335), .CI(\gdtr[25] ), .Z(O0[25]), .CO(n_337
		));
	notech_fa2 i_23(.A(I0[24]), .B(n_333), .CI(\gdtr[24] ), .Z(O0[24]), .CO(n_335
		));
	notech_fa2 i_22(.A(I0[23]), .B(n_331), .CI(\gdtr[23] ), .Z(O0[23]), .CO(n_333
		));
	notech_fa2 i_21(.A(I0[22]), .B(n_329), .CI(\gdtr[22] ), .Z(O0[22]), .CO(n_331
		));
	notech_fa2 i_20(.A(I0[21]), .B(n_327), .CI(\gdtr[21] ), .Z(O0[21]), .CO(n_329
		));
	notech_fa2 i_19(.A(I0[20]), .B(n_325), .CI(\gdtr[20] ), .Z(O0[20]), .CO(n_327
		));
	notech_fa2 i_18(.A(I0[19]), .B(n_323), .CI(\gdtr[19] ), .Z(O0[19]), .CO(n_325
		));
	notech_fa2 i_17(.A(I0[18]), .B(n_321), .CI(\gdtr[18] ), .Z(O0[18]), .CO(n_323
		));
	notech_fa2 i_16(.A(I0[17]), .B(n_319), .CI(\gdtr[17] ), .Z(O0[17]), .CO(n_321
		));
	notech_fa2 i_15(.A(I0[16]), .B(n_317), .CI(\gdtr[16] ), .Z(O0[16]), .CO(n_319
		));
	notech_fa2 i_14(.A(I0[15]), .B(n_315), .CI(\gdtr[15] ), .Z(O0[15]), .CO(n_317
		));
	notech_fa2 i_13(.A(I0[14]), .B(n_313), .CI(\gdtr[14] ), .Z(O0[14]), .CO(n_315
		));
	notech_fa2 i_12(.A(I0[13]), .B(n_311), .CI(\gdtr[13] ), .Z(O0[13]), .CO(n_313
		));
	notech_fa2 i_11(.A(I0[12]), .B(n_309), .CI(\gdtr[12] ), .Z(O0[12]), .CO(n_311
		));
	notech_fa2 i_10(.A(I0[11]), .B(n_307), .CI(\gdtr[11] ), .Z(O0[11]), .CO(n_309
		));
	notech_fa2 i_9(.A(I0[10]), .B(n_305), .CI(\gdtr[10] ), .Z(O0[10]), .CO(n_307
		));
	notech_fa2 i_8(.A(I0[9]), .B(n_303), .CI(\gdtr[9] ), .Z(O0[9]), .CO(n_305
		));
	notech_fa2 i_7(.A(I0[8]), .B(n_301), .CI(\gdtr[8] ), .Z(O0[8]), .CO(n_303
		));
	notech_fa2 i_6(.A(I0[7]), .B(n_299), .CI(\gdtr[7] ), .Z(O0[7]), .CO(n_301
		));
	notech_fa2 i_5(.A(I0[6]), .B(n_297), .CI(\gdtr[6] ), .Z(O0[6]), .CO(n_299
		));
	notech_fa2 i_4(.A(I0[5]), .B(n_295), .CI(\gdtr[5] ), .Z(O0[5]), .CO(n_297
		));
	notech_fa2 i_3(.A(I0[4]), .B(n_293), .CI(\gdtr[4] ), .Z(O0[4]), .CO(n_295
		));
	notech_fa2 i_2(.A(I0[3]), .B(n_354), .CI(\gdtr[3] ), .Z(O0[3]), .CO(n_293
		));
	notech_ha2 i_1(.A(\gdtr[2] ), .B(\gdtr[1] ), .Z(O0[2]), .CO(n_354));
	notech_inv i_0(.A(\gdtr[1] ), .Z(O0[1]));
endmodule
module AWDP_ADD_222(add_len_pc16, regs_14, lenpc);
    output [15:0] add_len_pc16;
    input [15:0] regs_14;
    input [15:0] lenpc;
    // Line 154
    wire [15:0] N236;
    // Line 156
    wire [15:0] add_len_pc16;

    // Line 154
    assign N236 = lenpc + regs_14;
    // Line 156
    assign add_len_pc16 = N236;
endmodule

module AWDP_ADD_239(O0, opd, I0);

	output [16:0] O0;
	input [15:0] opd;
	input [15:0] I0;




	notech_fa2 i_15(.A(I0[4]), .B(n_178), .CI(opd[15]), .Z(O0[15]), .CO(O0[
		16]));
	notech_fa2 i_14(.A(I0[4]), .B(n_176), .CI(opd[14]), .Z(O0[14]), .CO(n_178
		));
	notech_fa2 i_13(.A(I0[4]), .B(n_174), .CI(opd[13]), .Z(O0[13]), .CO(n_176
		));
	notech_fa2 i_12(.A(I0[4]), .B(n_172), .CI(opd[12]), .Z(O0[12]), .CO(n_174
		));
	notech_fa2 i_11(.A(I0[4]), .B(n_170), .CI(opd[11]), .Z(O0[11]), .CO(n_172
		));
	notech_fa2 i_10(.A(I0[4]), .B(n_168), .CI(opd[10]), .Z(O0[10]), .CO(n_170
		));
	notech_fa2 i_9(.A(I0[4]), .B(n_166), .CI(opd[9]), .Z(O0[9]), .CO(n_168)
		);
	notech_fa2 i_8(.A(I0[4]), .B(n_164), .CI(opd[8]), .Z(O0[8]), .CO(n_166)
		);
	notech_fa2 i_7(.A(I0[4]), .B(n_162), .CI(opd[7]), .Z(O0[7]), .CO(n_164)
		);
	notech_fa2 i_6(.A(I0[4]), .B(n_160), .CI(opd[6]), .Z(O0[6]), .CO(n_162)
		);
	notech_fa2 i_5(.A(I0[4]), .B(n_158), .CI(opd[5]), .Z(O0[5]), .CO(n_160)
		);
	notech_fa2 i_4(.A(I0[4]), .B(n_156), .CI(opd[4]), .Z(O0[4]), .CO(n_158)
		);
	notech_fa2 i_3(.A(I0[4]), .B(n_154), .CI(opd[3]), .Z(O0[3]), .CO(n_156)
		);
	notech_fa2 i_2(.A(I0[4]), .B(n_152), .CI(opd[2]), .Z(O0[2]), .CO(n_154)
		);
	notech_fa2 i_1(.A(I0[1]), .B(n_185), .CI(opd[1]), .Z(O0[1]), .CO(n_152)
		);
	notech_ha2 i_0(.A(opd[0]), .B(I0[0]), .Z(O0[0]), .CO(n_185));
endmodule
module AWDP_ADD_242(O0, opb, I0);

	output [31:0] O0;
	input [31:0] opb;
	input [31:0] I0;




	notech_ha2 i_31(.A(opb[31]), .B(n_400), .Z(O0[31]));
	notech_ha2 i_30(.A(opb[30]), .B(n_398), .Z(O0[30]), .CO(n_400));
	notech_ha2 i_29(.A(opb[29]), .B(n_396), .Z(O0[29]), .CO(n_398));
	notech_ha2 i_28(.A(opb[28]), .B(n_394), .Z(O0[28]), .CO(n_396));
	notech_ha2 i_27(.A(opb[27]), .B(n_392), .Z(O0[27]), .CO(n_394));
	notech_ha2 i_26(.A(opb[26]), .B(n_390), .Z(O0[26]), .CO(n_392));
	notech_ha2 i_25(.A(opb[25]), .B(n_388), .Z(O0[25]), .CO(n_390));
	notech_ha2 i_24(.A(opb[24]), .B(n_386), .Z(O0[24]), .CO(n_388));
	notech_ha2 i_23(.A(opb[23]), .B(n_384), .Z(O0[23]), .CO(n_386));
	notech_ha2 i_22(.A(opb[22]), .B(n_382), .Z(O0[22]), .CO(n_384));
	notech_ha2 i_21(.A(opb[21]), .B(n_380), .Z(O0[21]), .CO(n_382));
	notech_ha2 i_20(.A(opb[20]), .B(n_378), .Z(O0[20]), .CO(n_380));
	notech_ha2 i_19(.A(opb[19]), .B(n_376), .Z(O0[19]), .CO(n_378));
	notech_ha2 i_18(.A(opb[18]), .B(n_374), .Z(O0[18]), .CO(n_376));
	notech_ha2 i_17(.A(opb[17]), .B(n_372), .Z(O0[17]), .CO(n_374));
	notech_ha2 i_16(.A(opb[16]), .B(n_370), .Z(O0[16]), .CO(n_372));
	notech_ha2 i_15(.A(opb[15]), .B(n_368), .Z(O0[15]), .CO(n_370));
	notech_ha2 i_14(.A(opb[14]), .B(n_366), .Z(O0[14]), .CO(n_368));
	notech_ha2 i_13(.A(opb[13]), .B(n_364), .Z(O0[13]), .CO(n_366));
	notech_ha2 i_12(.A(opb[12]), .B(n_362), .Z(O0[12]), .CO(n_364));
	notech_ha2 i_11(.A(opb[11]), .B(n_360), .Z(O0[11]), .CO(n_362));
	notech_ha2 i_10(.A(opb[10]), .B(n_358), .Z(O0[10]), .CO(n_360));
	notech_ha2 i_9(.A(opb[9]), .B(n_356), .Z(O0[9]), .CO(n_358));
	notech_ha2 i_8(.A(opb[8]), .B(n_303), .Z(O0[8]), .CO(n_356));
	notech_fa2 i_7(.A(I0[7]), .B(n_301), .CI(opb[7]), .Z(O0[7]), .CO(n_303)
		);
	notech_fa2 i_6(.A(I0[6]), .B(n_299), .CI(opb[6]), .Z(O0[6]), .CO(n_301)
		);
	notech_fa2 i_5(.A(I0[5]), .B(n_297), .CI(opb[5]), .Z(O0[5]), .CO(n_299)
		);
	notech_fa2 i_4(.A(I0[4]), .B(n_295), .CI(opb[4]), .Z(O0[4]), .CO(n_297)
		);
	notech_fa2 i_3(.A(I0[3]), .B(n_293), .CI(opb[3]), .Z(O0[3]), .CO(n_295)
		);
	notech_fa2 i_2(.A(I0[2]), .B(n_291), .CI(opb[2]), .Z(O0[2]), .CO(n_293)
		);
	notech_fa2 i_1(.A(I0[1]), .B(n_354), .CI(opb[1]), .Z(O0[1]), .CO(n_291)
		);
	notech_ha2 i_0(.A(I0[0]), .B(opb[0]), .Z(O0[0]), .CO(n_354));
endmodule
module AWDP_ADD_33(add_len_pc32, regs_14, lenpc);
    output [31:0] add_len_pc32;
    input [31:0] regs_14;
    input [31:0] lenpc;
    // Line 156
    wire [31:0] add_len_pc32;
    // Line 155
    wire [31:0] N262;

    // Line 156
    assign add_len_pc32 = N262;
    // Line 155
    assign N262 = lenpc + regs_14;
endmodule

module AWDP_ADD_43(O0, I0, add_len_pc);
    output [31:0] O0;
    input [31:0] I0;
    input [31:0] add_len_pc;
    // Line 879
    wire [31:0] N336;
    // Line 386
    wire [31:0] O0;

    // Line 879
    assign N336 = I0 + add_len_pc;
    // Line 386
    assign O0 = N336;
endmodule

module AWDP_ADD_45(O0, regs_6, opd);
    output [31:0] O0;
    input [31:0] regs_6;
    input [31:0] opd;
    // Line 348
    wire [31:0] O0;
    // Line 520
    wire [31:0] N346;

    // Line 348
    assign O0 = N346;
    // Line 520
    assign N346 = regs_6 + opd;
endmodule

module AWDP_ADD_47(O0, opa, I0);

	output [16:0] O0;
	input [15:0] opa;
	input [15:0] I0;




	notech_fa2 i_15(.A(I0[13]), .B(n_178), .CI(opa[15]), .Z(O0[15]), .CO(O0[
		16]));
	notech_fa2 i_14(.A(I0[13]), .B(n_176), .CI(opa[14]), .Z(O0[14]), .CO(n_178
		));
	notech_fa2 i_13(.A(I0[13]), .B(n_174), .CI(opa[13]), .Z(O0[13]), .CO(n_176
		));
	notech_fa2 i_12(.A(I0[13]), .B(n_172), .CI(opa[12]), .Z(O0[12]), .CO(n_174
		));
	notech_fa2 i_11(.A(I0[13]), .B(n_170), .CI(opa[11]), .Z(O0[11]), .CO(n_172
		));
	notech_fa2 i_10(.A(I0[13]), .B(n_168), .CI(opa[10]), .Z(O0[10]), .CO(n_170
		));
	notech_fa2 i_9(.A(I0[13]), .B(n_166), .CI(opa[9]), .Z(O0[9]), .CO(n_168)
		);
	notech_fa2 i_8(.A(I0[13]), .B(n_164), .CI(opa[8]), .Z(O0[8]), .CO(n_166)
		);
	notech_fa2 i_7(.A(I0[13]), .B(n_162), .CI(opa[7]), .Z(O0[7]), .CO(n_164)
		);
	notech_fa2 i_6(.A(I0[13]), .B(n_160), .CI(opa[6]), .Z(O0[6]), .CO(n_162)
		);
	notech_fa2 i_5(.A(I0[13]), .B(n_158), .CI(opa[5]), .Z(O0[5]), .CO(n_160)
		);
	notech_fa2 i_4(.A(I0[13]), .B(n_156), .CI(opa[4]), .Z(O0[4]), .CO(n_158)
		);
	notech_fa2 i_3(.A(I0[13]), .B(n_154), .CI(opa[3]), .Z(O0[3]), .CO(n_156)
		);
	notech_fa2 i_2(.A(I0[13]), .B(n_152), .CI(opa[2]), .Z(O0[2]), .CO(n_154)
		);
	notech_fa2 i_1(.A(I0[1]), .B(n_185), .CI(opa[1]), .Z(O0[1]), .CO(n_152)
		);
	notech_ha2 i_0(.A(opa[0]), .B(I0[0]), .Z(O0[0]), .CO(n_185));
endmodule
module AWDP_ADD_52(O0, regs_7, opd);
    output [31:0] O0;
    input [31:0] regs_7;
    input [31:0] opd;
    // Line 348
    wire [31:0] O0;
    // Line 520
    wire [31:0] N366;

    // Line 348
    assign O0 = N366;
    // Line 520
    assign N366 = regs_7 + opd;
endmodule

module AWDP_ADD_6(O0, opa, opd);
    output [32:0] O0;
    input [31:0] opa;
    input [31:0] opd;
    // Line 599
    wire [32:0] N376;
    // Line 599
    wire [32:0] O0;

    // Line 599
    assign N376 = opa + opd;
    // Line 599
    assign O0 = N376;
endmodule

module AWDP_ADD_74(O0, Daddrs);

	output [31:0] O0;
	input [31:0] Daddrs;

	wire \Daddrs[1] ;
	wire \Daddrs[2] ;
	wire \Daddrs[3] ;
	wire \Daddrs[4] ;
	wire \Daddrs[5] ;
	wire \Daddrs[6] ;
	wire \Daddrs[7] ;
	wire \Daddrs[8] ;
	wire \Daddrs[9] ;
	wire \Daddrs[10] ;
	wire \Daddrs[11] ;
	wire \Daddrs[12] ;
	wire \Daddrs[13] ;
	wire \Daddrs[14] ;
	wire \Daddrs[15] ;
	wire \Daddrs[16] ;
	wire \Daddrs[17] ;
	wire \Daddrs[18] ;
	wire \Daddrs[19] ;
	wire \Daddrs[20] ;
	wire \Daddrs[21] ;
	wire \Daddrs[22] ;
	wire \Daddrs[23] ;
	wire \Daddrs[24] ;
	wire \Daddrs[25] ;
	wire \Daddrs[26] ;
	wire \Daddrs[27] ;
	wire \Daddrs[28] ;
	wire \Daddrs[29] ;
	wire \Daddrs[30] ;
	wire \Daddrs[31] ;


	assign O0[0] = Daddrs[0];
	assign \Daddrs[1]  = Daddrs[1];
	assign \Daddrs[2]  = Daddrs[2];
	assign \Daddrs[3]  = Daddrs[3];
	assign \Daddrs[4]  = Daddrs[4];
	assign \Daddrs[5]  = Daddrs[5];
	assign \Daddrs[6]  = Daddrs[6];
	assign \Daddrs[7]  = Daddrs[7];
	assign \Daddrs[8]  = Daddrs[8];
	assign \Daddrs[9]  = Daddrs[9];
	assign \Daddrs[10]  = Daddrs[10];
	assign \Daddrs[11]  = Daddrs[11];
	assign \Daddrs[12]  = Daddrs[12];
	assign \Daddrs[13]  = Daddrs[13];
	assign \Daddrs[14]  = Daddrs[14];
	assign \Daddrs[15]  = Daddrs[15];
	assign \Daddrs[16]  = Daddrs[16];
	assign \Daddrs[17]  = Daddrs[17];
	assign \Daddrs[18]  = Daddrs[18];
	assign \Daddrs[19]  = Daddrs[19];
	assign \Daddrs[20]  = Daddrs[20];
	assign \Daddrs[21]  = Daddrs[21];
	assign \Daddrs[22]  = Daddrs[22];
	assign \Daddrs[23]  = Daddrs[23];
	assign \Daddrs[24]  = Daddrs[24];
	assign \Daddrs[25]  = Daddrs[25];
	assign \Daddrs[26]  = Daddrs[26];
	assign \Daddrs[27]  = Daddrs[27];
	assign \Daddrs[28]  = Daddrs[28];
	assign \Daddrs[29]  = Daddrs[29];
	assign \Daddrs[30]  = Daddrs[30];
	assign \Daddrs[31]  = Daddrs[31];

	notech_ha2 i_30(.A(\Daddrs[31] ), .B(n_312), .Z(O0[31]));
	notech_ha2 i_29(.A(\Daddrs[30] ), .B(n_310), .Z(O0[30]), .CO(n_312));
	notech_ha2 i_28(.A(\Daddrs[29] ), .B(n_308), .Z(O0[29]), .CO(n_310));
	notech_ha2 i_27(.A(\Daddrs[28] ), .B(n_306), .Z(O0[28]), .CO(n_308));
	notech_ha2 i_26(.A(\Daddrs[27] ), .B(n_304), .Z(O0[27]), .CO(n_306));
	notech_ha2 i_25(.A(\Daddrs[26] ), .B(n_302), .Z(O0[26]), .CO(n_304));
	notech_ha2 i_24(.A(\Daddrs[25] ), .B(n_300), .Z(O0[25]), .CO(n_302));
	notech_ha2 i_23(.A(\Daddrs[24] ), .B(n_298), .Z(O0[24]), .CO(n_300));
	notech_ha2 i_22(.A(\Daddrs[23] ), .B(n_296), .Z(O0[23]), .CO(n_298));
	notech_ha2 i_21(.A(\Daddrs[22] ), .B(n_294), .Z(O0[22]), .CO(n_296));
	notech_ha2 i_20(.A(\Daddrs[21] ), .B(n_292), .Z(O0[21]), .CO(n_294));
	notech_ha2 i_19(.A(\Daddrs[20] ), .B(n_290), .Z(O0[20]), .CO(n_292));
	notech_ha2 i_18(.A(\Daddrs[19] ), .B(n_288), .Z(O0[19]), .CO(n_290));
	notech_ha2 i_17(.A(\Daddrs[18] ), .B(n_286), .Z(O0[18]), .CO(n_288));
	notech_ha2 i_16(.A(\Daddrs[17] ), .B(n_284), .Z(O0[17]), .CO(n_286));
	notech_ha2 i_15(.A(\Daddrs[16] ), .B(n_282), .Z(O0[16]), .CO(n_284));
	notech_ha2 i_14(.A(\Daddrs[15] ), .B(n_280), .Z(O0[15]), .CO(n_282));
	notech_ha2 i_13(.A(\Daddrs[14] ), .B(n_278), .Z(O0[14]), .CO(n_280));
	notech_ha2 i_12(.A(\Daddrs[13] ), .B(n_276), .Z(O0[13]), .CO(n_278));
	notech_ha2 i_11(.A(\Daddrs[12] ), .B(n_274), .Z(O0[12]), .CO(n_276));
	notech_ha2 i_10(.A(\Daddrs[11] ), .B(n_272), .Z(O0[11]), .CO(n_274));
	notech_ha2 i_9(.A(\Daddrs[10] ), .B(n_270), .Z(O0[10]), .CO(n_272));
	notech_ha2 i_8(.A(\Daddrs[9] ), .B(n_268), .Z(O0[9]), .CO(n_270));
	notech_ha2 i_7(.A(\Daddrs[8] ), .B(n_266), .Z(O0[8]), .CO(n_268));
	notech_ha2 i_6(.A(\Daddrs[7] ), .B(n_264), .Z(O0[7]), .CO(n_266));
	notech_ha2 i_5(.A(\Daddrs[6] ), .B(n_262), .Z(O0[6]), .CO(n_264));
	notech_ha2 i_4(.A(\Daddrs[5] ), .B(n_260), .Z(O0[5]), .CO(n_262));
	notech_ha2 i_3(.A(\Daddrs[4] ), .B(n_258), .Z(O0[4]), .CO(n_260));
	notech_ha2 i_2(.A(\Daddrs[3] ), .B(n_256), .Z(O0[3]), .CO(n_258));
	notech_ha2 i_1(.A(\Daddrs[2] ), .B(\Daddrs[1] ), .Z(O0[2]), .CO(n_256)
		);
	notech_inv i_0(.A(\Daddrs[1] ), .Z(O0[1]));
endmodule
module AWDP_ADD_84(O0, Daddrs);

	output [31:0] O0;
	input [31:0] Daddrs;

	wire \Daddrs[2] ;
	wire \Daddrs[3] ;
	wire \Daddrs[4] ;
	wire \Daddrs[5] ;
	wire \Daddrs[6] ;
	wire \Daddrs[7] ;
	wire \Daddrs[8] ;
	wire \Daddrs[9] ;
	wire \Daddrs[10] ;
	wire \Daddrs[11] ;
	wire \Daddrs[12] ;
	wire \Daddrs[13] ;
	wire \Daddrs[14] ;
	wire \Daddrs[15] ;
	wire \Daddrs[16] ;
	wire \Daddrs[17] ;
	wire \Daddrs[18] ;
	wire \Daddrs[19] ;
	wire \Daddrs[20] ;
	wire \Daddrs[21] ;
	wire \Daddrs[22] ;
	wire \Daddrs[23] ;
	wire \Daddrs[24] ;
	wire \Daddrs[25] ;
	wire \Daddrs[26] ;
	wire \Daddrs[27] ;
	wire \Daddrs[28] ;
	wire \Daddrs[29] ;
	wire \Daddrs[30] ;
	wire \Daddrs[31] ;


	assign O0[0] = Daddrs[0];
	assign O0[1] = Daddrs[1];
	assign \Daddrs[2]  = Daddrs[2];
	assign \Daddrs[3]  = Daddrs[3];
	assign \Daddrs[4]  = Daddrs[4];
	assign \Daddrs[5]  = Daddrs[5];
	assign \Daddrs[6]  = Daddrs[6];
	assign \Daddrs[7]  = Daddrs[7];
	assign \Daddrs[8]  = Daddrs[8];
	assign \Daddrs[9]  = Daddrs[9];
	assign \Daddrs[10]  = Daddrs[10];
	assign \Daddrs[11]  = Daddrs[11];
	assign \Daddrs[12]  = Daddrs[12];
	assign \Daddrs[13]  = Daddrs[13];
	assign \Daddrs[14]  = Daddrs[14];
	assign \Daddrs[15]  = Daddrs[15];
	assign \Daddrs[16]  = Daddrs[16];
	assign \Daddrs[17]  = Daddrs[17];
	assign \Daddrs[18]  = Daddrs[18];
	assign \Daddrs[19]  = Daddrs[19];
	assign \Daddrs[20]  = Daddrs[20];
	assign \Daddrs[21]  = Daddrs[21];
	assign \Daddrs[22]  = Daddrs[22];
	assign \Daddrs[23]  = Daddrs[23];
	assign \Daddrs[24]  = Daddrs[24];
	assign \Daddrs[25]  = Daddrs[25];
	assign \Daddrs[26]  = Daddrs[26];
	assign \Daddrs[27]  = Daddrs[27];
	assign \Daddrs[28]  = Daddrs[28];
	assign \Daddrs[29]  = Daddrs[29];
	assign \Daddrs[30]  = Daddrs[30];
	assign \Daddrs[31]  = Daddrs[31];

	notech_ha2 i_29(.A(\Daddrs[31] ), .B(n_308), .Z(O0[31]));
	notech_ha2 i_28(.A(\Daddrs[30] ), .B(n_306), .Z(O0[30]), .CO(n_308));
	notech_ha2 i_27(.A(\Daddrs[29] ), .B(n_304), .Z(O0[29]), .CO(n_306));
	notech_ha2 i_26(.A(\Daddrs[28] ), .B(n_302), .Z(O0[28]), .CO(n_304));
	notech_ha2 i_25(.A(\Daddrs[27] ), .B(n_300), .Z(O0[27]), .CO(n_302));
	notech_ha2 i_24(.A(\Daddrs[26] ), .B(n_298), .Z(O0[26]), .CO(n_300));
	notech_ha2 i_23(.A(\Daddrs[25] ), .B(n_296), .Z(O0[25]), .CO(n_298));
	notech_ha2 i_22(.A(\Daddrs[24] ), .B(n_294), .Z(O0[24]), .CO(n_296));
	notech_ha2 i_21(.A(\Daddrs[23] ), .B(n_292), .Z(O0[23]), .CO(n_294));
	notech_ha2 i_20(.A(\Daddrs[22] ), .B(n_290), .Z(O0[22]), .CO(n_292));
	notech_ha2 i_19(.A(\Daddrs[21] ), .B(n_288), .Z(O0[21]), .CO(n_290));
	notech_ha2 i_18(.A(\Daddrs[20] ), .B(n_286), .Z(O0[20]), .CO(n_288));
	notech_ha2 i_17(.A(\Daddrs[19] ), .B(n_284), .Z(O0[19]), .CO(n_286));
	notech_ha2 i_16(.A(\Daddrs[18] ), .B(n_282), .Z(O0[18]), .CO(n_284));
	notech_ha2 i_15(.A(\Daddrs[17] ), .B(n_280), .Z(O0[17]), .CO(n_282));
	notech_ha2 i_14(.A(\Daddrs[16] ), .B(n_278), .Z(O0[16]), .CO(n_280));
	notech_ha2 i_13(.A(\Daddrs[15] ), .B(n_276), .Z(O0[15]), .CO(n_278));
	notech_ha2 i_12(.A(\Daddrs[14] ), .B(n_274), .Z(O0[14]), .CO(n_276));
	notech_ha2 i_11(.A(\Daddrs[13] ), .B(n_272), .Z(O0[13]), .CO(n_274));
	notech_ha2 i_10(.A(\Daddrs[12] ), .B(n_270), .Z(O0[12]), .CO(n_272));
	notech_ha2 i_9(.A(\Daddrs[11] ), .B(n_268), .Z(O0[11]), .CO(n_270));
	notech_ha2 i_8(.A(\Daddrs[10] ), .B(n_266), .Z(O0[10]), .CO(n_268));
	notech_ha2 i_7(.A(\Daddrs[9] ), .B(n_264), .Z(O0[9]), .CO(n_266));
	notech_ha2 i_6(.A(\Daddrs[8] ), .B(n_262), .Z(O0[8]), .CO(n_264));
	notech_ha2 i_5(.A(\Daddrs[7] ), .B(n_260), .Z(O0[7]), .CO(n_262));
	notech_ha2 i_4(.A(\Daddrs[6] ), .B(n_258), .Z(O0[6]), .CO(n_260));
	notech_ha2 i_3(.A(\Daddrs[5] ), .B(n_256), .Z(O0[5]), .CO(n_258));
	notech_ha2 i_2(.A(\Daddrs[4] ), .B(n_254), .Z(O0[4]), .CO(n_256));
	notech_ha2 i_1(.A(\Daddrs[3] ), .B(\Daddrs[2] ), .Z(O0[3]), .CO(n_254)
		);
	notech_inv i_0(.A(\Daddrs[2] ), .Z(O0[2]));
endmodule
module AWDP_DEC_143(O0, opc);

	output [31:0] O0;
	input [31:0] opc;




	notech_ha2 i_32(.A(n_192), .B(n_254), .Z(O0[31]));
	notech_inv i_1(.A(opc[0]), .Z(O0[0]));
	notech_inv i_0(.A(opc[31]), .Z(n_192));
	notech_xor2 i_54141(.A(opc[30]), .B(n_252), .Z(n_44785));
	notech_inv i_54142(.A(n_44785), .Z(O0[30]));
	notech_or2 i_54140(.A(opc[30]), .B(n_252), .Z(n_254));
	notech_xor2 i_48(.A(opc[29]), .B(n_250), .Z(n_44812));
	notech_inv i_49(.A(n_44812), .Z(O0[29]));
	notech_or2 i_47(.A(opc[29]), .B(n_250), .Z(n_252));
	notech_xor2 i_46(.A(opc[28]), .B(n_248), .Z(n_44839));
	notech_inv i_4798764(.A(n_44839), .Z(O0[28]));
	notech_or2 i_45(.A(opc[28]), .B(n_248), .Z(n_250));
	notech_xor2 i_4598765(.A(opc[27]), .B(n_246), .Z(n_44866));
	notech_inv i_4698766(.A(n_44866), .Z(O0[27]));
	notech_or2 i_44(.A(opc[27]), .B(n_246), .Z(n_248));
	notech_xor2 i_4498767(.A(opc[26]), .B(n_244), .Z(n_44893));
	notech_inv i_4598768(.A(n_44893), .Z(O0[26]));
	notech_or2 i_43(.A(opc[26]), .B(n_244), .Z(n_246));
	notech_xor2 i_4398769(.A(opc[25]), .B(n_242), .Z(n_44920));
	notech_inv i_4498770(.A(n_44920), .Z(O0[25]));
	notech_or2 i_42(.A(opc[25]), .B(n_242), .Z(n_244));
	notech_xor2 i_4298771(.A(opc[24]), .B(n_240), .Z(n_44947));
	notech_inv i_4398772(.A(n_44947), .Z(O0[24]));
	notech_or2 i_41(.A(opc[24]), .B(n_240), .Z(n_242));
	notech_xor2 i_4198773(.A(opc[23]), .B(n_238), .Z(n_44974));
	notech_inv i_4298774(.A(n_44974), .Z(O0[23]));
	notech_or2 i_40(.A(opc[23]), .B(n_238), .Z(n_240));
	notech_xor2 i_4098775(.A(opc[22]), .B(n_236), .Z(n_45001));
	notech_inv i_4198776(.A(n_45001), .Z(O0[22]));
	notech_or2 i_39(.A(opc[22]), .B(n_236), .Z(n_238));
	notech_xor2 i_3998777(.A(opc[21]), .B(n_234), .Z(n_45028));
	notech_inv i_4098778(.A(n_45028), .Z(O0[21]));
	notech_or2 i_38(.A(opc[21]), .B(n_234), .Z(n_236));
	notech_xor2 i_3898779(.A(opc[20]), .B(n_232), .Z(n_45055));
	notech_inv i_3998780(.A(n_45055), .Z(O0[20]));
	notech_or2 i_37(.A(opc[20]), .B(n_232), .Z(n_234));
	notech_xor2 i_3798781(.A(opc[19]), .B(n_230), .Z(n_45082));
	notech_inv i_3898782(.A(n_45082), .Z(O0[19]));
	notech_or2 i_36(.A(opc[19]), .B(n_230), .Z(n_232));
	notech_xor2 i_3698783(.A(opc[18]), .B(n_228), .Z(n_45109));
	notech_inv i_3798784(.A(n_45109), .Z(O0[18]));
	notech_or2 i_35(.A(opc[18]), .B(n_228), .Z(n_230));
	notech_xor2 i_3598785(.A(opc[17]), .B(n_226), .Z(n_45136));
	notech_inv i_3698786(.A(n_45136), .Z(O0[17]));
	notech_or2 i_34(.A(opc[17]), .B(n_226), .Z(n_228));
	notech_xor2 i_3498787(.A(opc[16]), .B(n_224), .Z(n_45163));
	notech_inv i_3598788(.A(n_45163), .Z(O0[16]));
	notech_or2 i_33(.A(opc[16]), .B(n_224), .Z(n_226));
	notech_xor2 i_3398789(.A(opc[15]), .B(n_222), .Z(n_45190));
	notech_inv i_3498790(.A(n_45190), .Z(O0[15]));
	notech_or2 i_3298791(.A(opc[15]), .B(n_222), .Z(n_224));
	notech_xor2 i_3298792(.A(opc[14]), .B(n_220), .Z(n_45217));
	notech_inv i_3398793(.A(n_45217), .Z(O0[14]));
	notech_or2 i_31(.A(opc[14]), .B(n_220), .Z(n_222));
	notech_xor2 i_3198794(.A(opc[13]), .B(n_218), .Z(n_45244));
	notech_inv i_3298795(.A(n_45244), .Z(O0[13]));
	notech_or2 i_30(.A(opc[13]), .B(n_218), .Z(n_220));
	notech_xor2 i_3098796(.A(opc[12]), .B(n_216), .Z(n_45271));
	notech_inv i_3198797(.A(n_45271), .Z(O0[12]));
	notech_or2 i_29(.A(opc[12]), .B(n_216), .Z(n_218));
	notech_xor2 i_2998798(.A(opc[11]), .B(n_214), .Z(n_45298));
	notech_inv i_3098799(.A(n_45298), .Z(O0[11]));
	notech_or2 i_28(.A(opc[11]), .B(n_214), .Z(n_216));
	notech_xor2 i_2898800(.A(opc[10]), .B(n_212), .Z(n_45325));
	notech_inv i_2998801(.A(n_45325), .Z(O0[10]));
	notech_or2 i_27(.A(opc[10]), .B(n_212), .Z(n_214));
	notech_xor2 i_2798802(.A(opc[9]), .B(n_210), .Z(n_45352));
	notech_inv i_2898803(.A(n_45352), .Z(O0[9]));
	notech_or2 i_26(.A(opc[9]), .B(n_210), .Z(n_212));
	notech_xor2 i_2798804(.A(opc[8]), .B(n_208), .Z(n_45379));
	notech_inv i_2898805(.A(n_45379), .Z(O0[8]));
	notech_or2 i_2698806(.A(opc[8]), .B(n_208), .Z(n_210));
	notech_xor2 i_2798807(.A(opc[7]), .B(n_206), .Z(n_45406));
	notech_inv i_2898808(.A(n_45406), .Z(O0[7]));
	notech_or2 i_2698809(.A(opc[7]), .B(n_206), .Z(n_208));
	notech_xor2 i_2798810(.A(opc[6]), .B(n_204), .Z(n_45433));
	notech_inv i_2898811(.A(n_45433), .Z(O0[6]));
	notech_or2 i_2698812(.A(opc[6]), .B(n_204), .Z(n_206));
	notech_xor2 i_2798813(.A(opc[5]), .B(n_202), .Z(n_45460));
	notech_inv i_2898814(.A(n_45460), .Z(O0[5]));
	notech_or2 i_2698815(.A(opc[5]), .B(n_202), .Z(n_204));
	notech_xor2 i_2798816(.A(opc[4]), .B(n_200), .Z(n_45487));
	notech_inv i_2898817(.A(n_45487), .Z(O0[4]));
	notech_or2 i_2698818(.A(opc[4]), .B(n_200), .Z(n_202));
	notech_xor2 i_2798819(.A(opc[3]), .B(n_198), .Z(n_45514));
	notech_inv i_2898820(.A(n_45514), .Z(O0[3]));
	notech_or2 i_2698821(.A(opc[3]), .B(n_198), .Z(n_200));
	notech_xor2 i_2798822(.A(opc[2]), .B(n_196), .Z(n_45541));
	notech_inv i_2898823(.A(n_45541), .Z(O0[2]));
	notech_or2 i_2698824(.A(opc[2]), .B(n_196), .Z(n_198));
	notech_xor2 i_2798825(.A(opc[1]), .B(opc[0]), .Z(n_45569));
	notech_inv i_2898826(.A(n_45569), .Z(O0[1]));
	notech_or2 i_2698827(.A(opc[1]), .B(opc[0]), .Z(n_196));
endmodule
module AWDP_DEC_206(O0, cx);

	output [15:0] O0;
	input [15:0] cx;




	notech_ha2 i_16(.A(n_96), .B(n_126), .Z(O0[15]));
	notech_inv i_1(.A(cx[0]), .Z(O0[0]));
	notech_inv i_0(.A(cx[15]), .Z(n_96));
	notech_xor2 i_33(.A(cx[14]), .B(n_124), .Z(n_45596));
	notech_inv i_34(.A(n_45596), .Z(O0[14]));
	notech_or2 i_32(.A(cx[14]), .B(n_124), .Z(n_126));
	notech_xor2 i_3298828(.A(cx[13]), .B(n_122), .Z(n_45623));
	notech_inv i_3398829(.A(n_45623), .Z(O0[13]));
	notech_or2 i_31(.A(cx[13]), .B(n_122), .Z(n_124));
	notech_xor2 i_30(.A(cx[12]), .B(n_120), .Z(n_45650));
	notech_inv i_3198830(.A(n_45650), .Z(O0[12]));
	notech_or2 i_29(.A(cx[12]), .B(n_120), .Z(n_122));
	notech_xor2 i_2998831(.A(cx[11]), .B(n_118), .Z(n_45677));
	notech_inv i_3098832(.A(n_45677), .Z(O0[11]));
	notech_or2 i_28(.A(cx[11]), .B(n_118), .Z(n_120));
	notech_xor2 i_2898833(.A(cx[10]), .B(n_116), .Z(n_45704));
	notech_inv i_2998834(.A(n_45704), .Z(O0[10]));
	notech_or2 i_27(.A(cx[10]), .B(n_116), .Z(n_118));
	notech_xor2 i_2798835(.A(cx[9]), .B(n_114), .Z(n_45731));
	notech_inv i_2898836(.A(n_45731), .Z(O0[9]));
	notech_or2 i_26(.A(cx[9]), .B(n_114), .Z(n_116));
	notech_xor2 i_2798837(.A(cx[8]), .B(n_112), .Z(n_45758));
	notech_inv i_2898838(.A(n_45758), .Z(O0[8]));
	notech_or2 i_2698839(.A(cx[8]), .B(n_112), .Z(n_114));
	notech_xor2 i_2798840(.A(cx[7]), .B(n_110), .Z(n_45785));
	notech_inv i_2898841(.A(n_45785), .Z(O0[7]));
	notech_or2 i_2698842(.A(cx[7]), .B(n_110), .Z(n_112));
	notech_xor2 i_2798843(.A(cx[6]), .B(n_108), .Z(n_45812));
	notech_inv i_2898844(.A(n_45812), .Z(O0[6]));
	notech_or2 i_2698845(.A(cx[6]), .B(n_108), .Z(n_110));
	notech_xor2 i_2798846(.A(cx[5]), .B(n_106), .Z(n_45839));
	notech_inv i_2898847(.A(n_45839), .Z(O0[5]));
	notech_or2 i_2698848(.A(cx[5]), .B(n_106), .Z(n_108));
	notech_xor2 i_2798849(.A(cx[4]), .B(n_104), .Z(n_45866));
	notech_inv i_2898850(.A(n_45866), .Z(O0[4]));
	notech_or2 i_2698851(.A(cx[4]), .B(n_104), .Z(n_106));
	notech_xor2 i_2798852(.A(cx[3]), .B(n_102), .Z(n_45893));
	notech_inv i_2898853(.A(n_45893), .Z(O0[3]));
	notech_or2 i_2698854(.A(cx[3]), .B(n_102), .Z(n_104));
	notech_xor2 i_2798855(.A(cx[2]), .B(n_100), .Z(n_45920));
	notech_inv i_2898856(.A(n_45920), .Z(O0[2]));
	notech_or2 i_2698857(.A(cx[2]), .B(n_100), .Z(n_102));
	notech_xor2 i_2798858(.A(cx[1]), .B(cx[0]), .Z(n_45948));
	notech_inv i_2898859(.A(n_45948), .Z(O0[1]));
	notech_or2 i_2698860(.A(cx[1]), .B(cx[0]), .Z(n_100));
endmodule
module AWDP_DEC_236(O0, ecx);

	output [31:0] O0;
	input [31:0] ecx;




	notech_ha2 i_32(.A(n_192), .B(n_254), .Z(O0[31]));
	notech_inv i_1(.A(ecx[0]), .Z(O0[0]));
	notech_inv i_0(.A(ecx[31]), .Z(n_192));
	notech_xor2 i_49(.A(ecx[30]), .B(n_252), .Z(n_45975));
	notech_inv i_50(.A(n_45975), .Z(O0[30]));
	notech_or2 i_48(.A(ecx[30]), .B(n_252), .Z(n_254));
	notech_xor2 i_4898861(.A(ecx[29]), .B(n_250), .Z(n_46002));
	notech_inv i_4998862(.A(n_46002), .Z(O0[29]));
	notech_or2 i_47(.A(ecx[29]), .B(n_250), .Z(n_252));
	notech_xor2 i_46(.A(ecx[28]), .B(n_248), .Z(n_46029));
	notech_inv i_4798863(.A(n_46029), .Z(O0[28]));
	notech_or2 i_45(.A(ecx[28]), .B(n_248), .Z(n_250));
	notech_xor2 i_4598864(.A(ecx[27]), .B(n_246), .Z(n_46056));
	notech_inv i_4698865(.A(n_46056), .Z(O0[27]));
	notech_or2 i_44(.A(ecx[27]), .B(n_246), .Z(n_248));
	notech_xor2 i_4498866(.A(ecx[26]), .B(n_244), .Z(n_46083));
	notech_inv i_4598867(.A(n_46083), .Z(O0[26]));
	notech_or2 i_43(.A(ecx[26]), .B(n_244), .Z(n_246));
	notech_xor2 i_4398868(.A(ecx[25]), .B(n_242), .Z(n_46110));
	notech_inv i_4498869(.A(n_46110), .Z(O0[25]));
	notech_or2 i_42(.A(ecx[25]), .B(n_242), .Z(n_244));
	notech_xor2 i_4298870(.A(ecx[24]), .B(n_240), .Z(n_46137));
	notech_inv i_4398871(.A(n_46137), .Z(O0[24]));
	notech_or2 i_41(.A(ecx[24]), .B(n_240), .Z(n_242));
	notech_xor2 i_4198872(.A(ecx[23]), .B(n_238), .Z(n_46164));
	notech_inv i_4298873(.A(n_46164), .Z(O0[23]));
	notech_or2 i_40(.A(ecx[23]), .B(n_238), .Z(n_240));
	notech_xor2 i_4098874(.A(ecx[22]), .B(n_236), .Z(n_46191));
	notech_inv i_4198875(.A(n_46191), .Z(O0[22]));
	notech_or2 i_39(.A(ecx[22]), .B(n_236), .Z(n_238));
	notech_xor2 i_3998876(.A(ecx[21]), .B(n_234), .Z(n_46218));
	notech_inv i_4098877(.A(n_46218), .Z(O0[21]));
	notech_or2 i_38(.A(ecx[21]), .B(n_234), .Z(n_236));
	notech_xor2 i_3898878(.A(ecx[20]), .B(n_232), .Z(n_46245));
	notech_inv i_3998879(.A(n_46245), .Z(O0[20]));
	notech_or2 i_37(.A(ecx[20]), .B(n_232), .Z(n_234));
	notech_xor2 i_3798880(.A(ecx[19]), .B(n_230), .Z(n_46272));
	notech_inv i_3898881(.A(n_46272), .Z(O0[19]));
	notech_or2 i_36(.A(ecx[19]), .B(n_230), .Z(n_232));
	notech_xor2 i_3698882(.A(ecx[18]), .B(n_228), .Z(n_46299));
	notech_inv i_3798883(.A(n_46299), .Z(O0[18]));
	notech_or2 i_35(.A(ecx[18]), .B(n_228), .Z(n_230));
	notech_xor2 i_3598884(.A(ecx[17]), .B(n_226), .Z(n_46326));
	notech_inv i_3698885(.A(n_46326), .Z(O0[17]));
	notech_or2 i_34(.A(ecx[17]), .B(n_226), .Z(n_228));
	notech_xor2 i_3498886(.A(ecx[16]), .B(n_224), .Z(n_46353));
	notech_inv i_3598887(.A(n_46353), .Z(O0[16]));
	notech_or2 i_33(.A(ecx[16]), .B(n_224), .Z(n_226));
	notech_xor2 i_3398888(.A(ecx[15]), .B(n_222), .Z(n_46380));
	notech_inv i_3498889(.A(n_46380), .Z(O0[15]));
	notech_or2 i_3298890(.A(ecx[15]), .B(n_222), .Z(n_224));
	notech_xor2 i_3298891(.A(ecx[14]), .B(n_220), .Z(n_46407));
	notech_inv i_3398892(.A(n_46407), .Z(O0[14]));
	notech_or2 i_31(.A(ecx[14]), .B(n_220), .Z(n_222));
	notech_xor2 i_3198893(.A(ecx[13]), .B(n_218), .Z(n_46434));
	notech_inv i_3298894(.A(n_46434), .Z(O0[13]));
	notech_or2 i_30(.A(ecx[13]), .B(n_218), .Z(n_220));
	notech_xor2 i_3098895(.A(ecx[12]), .B(n_216), .Z(n_46461));
	notech_inv i_3198896(.A(n_46461), .Z(O0[12]));
	notech_or2 i_29(.A(ecx[12]), .B(n_216), .Z(n_218));
	notech_xor2 i_2998897(.A(ecx[11]), .B(n_214), .Z(n_46488));
	notech_inv i_3098898(.A(n_46488), .Z(O0[11]));
	notech_or2 i_28(.A(ecx[11]), .B(n_214), .Z(n_216));
	notech_xor2 i_2898899(.A(ecx[10]), .B(n_212), .Z(n_46515));
	notech_inv i_2998900(.A(n_46515), .Z(O0[10]));
	notech_or2 i_27(.A(ecx[10]), .B(n_212), .Z(n_214));
	notech_xor2 i_2798901(.A(ecx[9]), .B(n_210), .Z(n_46542));
	notech_inv i_2898902(.A(n_46542), .Z(O0[9]));
	notech_or2 i_26(.A(ecx[9]), .B(n_210), .Z(n_212));
	notech_xor2 i_2798903(.A(ecx[8]), .B(n_208), .Z(n_46569));
	notech_inv i_2898904(.A(n_46569), .Z(O0[8]));
	notech_or2 i_2698905(.A(ecx[8]), .B(n_208), .Z(n_210));
	notech_xor2 i_2798906(.A(ecx[7]), .B(n_206), .Z(n_46596));
	notech_inv i_2898907(.A(n_46596), .Z(O0[7]));
	notech_or2 i_2698908(.A(ecx[7]), .B(n_206), .Z(n_208));
	notech_xor2 i_2798909(.A(ecx[6]), .B(n_204), .Z(n_46623));
	notech_inv i_2898910(.A(n_46623), .Z(O0[6]));
	notech_or2 i_2698911(.A(ecx[6]), .B(n_204), .Z(n_206));
	notech_xor2 i_2798912(.A(ecx[5]), .B(n_202), .Z(n_46650));
	notech_inv i_2898913(.A(n_46650), .Z(O0[5]));
	notech_or2 i_2698914(.A(ecx[5]), .B(n_202), .Z(n_204));
	notech_xor2 i_2798915(.A(ecx[4]), .B(n_200), .Z(n_46677));
	notech_inv i_2898916(.A(n_46677), .Z(O0[4]));
	notech_or2 i_2698917(.A(ecx[4]), .B(n_200), .Z(n_202));
	notech_xor2 i_2798918(.A(ecx[3]), .B(n_198), .Z(n_46704));
	notech_inv i_2898919(.A(n_46704), .Z(O0[3]));
	notech_or2 i_2698920(.A(ecx[3]), .B(n_198), .Z(n_200));
	notech_xor2 i_2798921(.A(ecx[2]), .B(n_196), .Z(n_46731));
	notech_inv i_2898922(.A(n_46731), .Z(O0[2]));
	notech_or2 i_2698923(.A(ecx[2]), .B(n_196), .Z(n_198));
	notech_xor2 i_2798924(.A(ecx[1]), .B(ecx[0]), .Z(n_46759));
	notech_inv i_2898925(.A(n_46759), .Z(O0[1]));
	notech_or2 i_2698926(.A(ecx[1]), .B(ecx[0]), .Z(n_196));
endmodule
module AWDP_DEC_7(O0, opc);

	output [7:0] O0;
	input [7:0] opc;




	notech_ha2 i_8(.A(n_48), .B(n_62), .Z(O0[7]));
	notech_inv i_1(.A(opc[0]), .Z(O0[0]));
	notech_inv i_0(.A(opc[7]), .Z(n_48));
	notech_xor2 i_30(.A(opc[6]), .B(n_60), .Z(n_46786));
	notech_inv i_31(.A(n_46786), .Z(O0[6]));
	notech_or2 i_29(.A(opc[6]), .B(n_60), .Z(n_62));
	notech_xor2 i_27(.A(opc[5]), .B(n_58), .Z(n_46813));
	notech_inv i_28(.A(n_46813), .Z(O0[5]));
	notech_or2 i_26(.A(opc[5]), .B(n_58), .Z(n_60));
	notech_xor2 i_2798927(.A(opc[4]), .B(n_56), .Z(n_46840));
	notech_inv i_2898928(.A(n_46840), .Z(O0[4]));
	notech_or2 i_2698929(.A(opc[4]), .B(n_56), .Z(n_58));
	notech_xor2 i_2798930(.A(opc[3]), .B(n_54), .Z(n_46867));
	notech_inv i_2898931(.A(n_46867), .Z(O0[3]));
	notech_or2 i_2698932(.A(opc[3]), .B(n_54), .Z(n_56));
	notech_xor2 i_2798933(.A(opc[2]), .B(n_52), .Z(n_46894));
	notech_inv i_2898934(.A(n_46894), .Z(O0[2]));
	notech_or2 i_2698935(.A(opc[2]), .B(n_52), .Z(n_54));
	notech_xor2 i_2798936(.A(opc[1]), .B(opc[0]), .Z(n_46922));
	notech_inv i_2898937(.A(n_46922), .Z(O0[1]));
	notech_or2 i_2698938(.A(opc[1]), .B(opc[0]), .Z(n_52));
endmodule
module AWDP_EQ_138(O0, I0, I1);
    output [0:0] O0;
    input [63:0] I0;
    input [63:0] I1;
    // Line 790
    wire [0:0] N524;
    // Line 790
    wire [0:0] O0;

    // Line 790
    assign N524 = I0 == I1;
    // Line 790
    assign O0 = N524;
endmodule

module AWDP_EQ_174(O0, mul64);
    output [0:0] O0;
    input [63:16] mul64;
    // Line 126
    wire [0:0] N555;
    // Line 126
    wire [0:0] O0;

    // Line 126
    assign N555 = mul64 == 48'h0;
    // Line 126
    assign O0 = N555;
endmodule

module AWDP_EQ_205(O0, mul64);
    output [0:0] O0;
    input [63:32] mul64;
    // Line 131
    wire [0:0] N564;
    // Line 131
    wire [0:0] O0;

    // Line 131
    assign N564 = mul64 == 32'hffffffff;
    // Line 131
    assign O0 = N564;
endmodule

module AWDP_EQ_24111880(O0, mul64);
    output [0:0] O0;
    input [63:16] mul64;
    // Line 130
    wire [0:0] N577;
    // Line 130
    wire [0:0] O0;

    // Line 130
    assign N577 = mul64 == 48'hffffffff;
    // Line 130
    assign O0 = N577;
endmodule

module AWDP_EQ_85(O0, mul64);
    output [0:0] O0;
    input [63:8] mul64;
    // Line 125
    wire [0:0] O0;
    // Line 125
    wire [0:0] N607;

    // Line 125
    assign O0 = N607;
    // Line 125
    assign N607 = mul64 == 56'h0;
endmodule

module AWDP_EQ_91(O0, mul64);
    output [0:0] O0;
    input [63:8] mul64;
    // Line 129
    wire [0:0] N620;
    // Line 129
    wire [0:0] O0;

    // Line 129
    assign N620 = mul64 == 56'hffffffff;
    // Line 129
    assign O0 = N620;
endmodule

module AWDP_GE_13(O0, divr, divq);
    output [0:0] O0;
    input [63:0] divr;
    input [63:0] divq;
    // Line 1006
    wire [0:0] N627;
    // Line 1006
    wire [0:0] O0;

    // Line 1006
    assign N627 = divr >= divq;
    // Line 1006
    assign O0 = N627;
endmodule

module AWDP_INC_0(O0, tsc);

	output [63:0] O0;
	input [63:0] tsc;




	notech_ha2 i_63(.A(tsc[63]), .B(n_636), .Z(O0[63]));
	notech_ha2 i_62(.A(tsc[62]), .B(n_634), .Z(O0[62]), .CO(n_636));
	notech_ha2 i_61(.A(tsc[61]), .B(n_632), .Z(O0[61]), .CO(n_634));
	notech_ha2 i_60(.A(tsc[60]), .B(n_630), .Z(O0[60]), .CO(n_632));
	notech_ha2 i_59(.A(tsc[59]), .B(n_628), .Z(O0[59]), .CO(n_630));
	notech_ha2 i_58(.A(tsc[58]), .B(n_626), .Z(O0[58]), .CO(n_628));
	notech_ha2 i_57(.A(tsc[57]), .B(n_624), .Z(O0[57]), .CO(n_626));
	notech_ha2 i_56(.A(tsc[56]), .B(n_622), .Z(O0[56]), .CO(n_624));
	notech_ha2 i_55(.A(tsc[55]), .B(n_620), .Z(O0[55]), .CO(n_622));
	notech_ha2 i_54(.A(tsc[54]), .B(n_618), .Z(O0[54]), .CO(n_620));
	notech_ha2 i_53(.A(tsc[53]), .B(n_616), .Z(O0[53]), .CO(n_618));
	notech_ha2 i_52(.A(tsc[52]), .B(n_614), .Z(O0[52]), .CO(n_616));
	notech_ha2 i_51(.A(tsc[51]), .B(n_612), .Z(O0[51]), .CO(n_614));
	notech_ha2 i_50(.A(tsc[50]), .B(n_610), .Z(O0[50]), .CO(n_612));
	notech_ha2 i_49(.A(tsc[49]), .B(n_608), .Z(O0[49]), .CO(n_610));
	notech_ha2 i_48(.A(tsc[48]), .B(n_606), .Z(O0[48]), .CO(n_608));
	notech_ha2 i_47(.A(tsc[47]), .B(n_604), .Z(O0[47]), .CO(n_606));
	notech_ha2 i_46(.A(tsc[46]), .B(n_602), .Z(O0[46]), .CO(n_604));
	notech_ha2 i_45(.A(tsc[45]), .B(n_600), .Z(O0[45]), .CO(n_602));
	notech_ha2 i_44(.A(tsc[44]), .B(n_598), .Z(O0[44]), .CO(n_600));
	notech_ha2 i_43(.A(tsc[43]), .B(n_596), .Z(O0[43]), .CO(n_598));
	notech_ha2 i_42(.A(tsc[42]), .B(n_594), .Z(O0[42]), .CO(n_596));
	notech_ha2 i_41(.A(tsc[41]), .B(n_592), .Z(O0[41]), .CO(n_594));
	notech_ha2 i_40(.A(tsc[40]), .B(n_590), .Z(O0[40]), .CO(n_592));
	notech_ha2 i_39(.A(tsc[39]), .B(n_588), .Z(O0[39]), .CO(n_590));
	notech_ha2 i_38(.A(tsc[38]), .B(n_586), .Z(O0[38]), .CO(n_588));
	notech_ha2 i_37(.A(tsc[37]), .B(n_584), .Z(O0[37]), .CO(n_586));
	notech_ha2 i_36(.A(tsc[36]), .B(n_582), .Z(O0[36]), .CO(n_584));
	notech_ha2 i_35(.A(tsc[35]), .B(n_580), .Z(O0[35]), .CO(n_582));
	notech_ha2 i_34(.A(tsc[34]), .B(n_578), .Z(O0[34]), .CO(n_580));
	notech_ha2 i_33(.A(tsc[33]), .B(n_576), .Z(O0[33]), .CO(n_578));
	notech_ha2 i_32(.A(tsc[32]), .B(n_574), .Z(O0[32]), .CO(n_576));
	notech_ha2 i_31(.A(tsc[31]), .B(n_572), .Z(O0[31]), .CO(n_574));
	notech_ha2 i_30(.A(tsc[30]), .B(n_570), .Z(O0[30]), .CO(n_572));
	notech_ha2 i_29(.A(tsc[29]), .B(n_568), .Z(O0[29]), .CO(n_570));
	notech_ha2 i_28(.A(tsc[28]), .B(n_566), .Z(O0[28]), .CO(n_568));
	notech_ha2 i_27(.A(tsc[27]), .B(n_564), .Z(O0[27]), .CO(n_566));
	notech_ha2 i_26(.A(tsc[26]), .B(n_562), .Z(O0[26]), .CO(n_564));
	notech_ha2 i_25(.A(tsc[25]), .B(n_560), .Z(O0[25]), .CO(n_562));
	notech_ha2 i_24(.A(tsc[24]), .B(n_558), .Z(O0[24]), .CO(n_560));
	notech_ha2 i_23(.A(tsc[23]), .B(n_556), .Z(O0[23]), .CO(n_558));
	notech_ha2 i_22(.A(tsc[22]), .B(n_554), .Z(O0[22]), .CO(n_556));
	notech_ha2 i_21(.A(tsc[21]), .B(n_552), .Z(O0[21]), .CO(n_554));
	notech_ha2 i_20(.A(tsc[20]), .B(n_550), .Z(O0[20]), .CO(n_552));
	notech_ha2 i_19(.A(tsc[19]), .B(n_548), .Z(O0[19]), .CO(n_550));
	notech_ha2 i_18(.A(tsc[18]), .B(n_546), .Z(O0[18]), .CO(n_548));
	notech_ha2 i_17(.A(tsc[17]), .B(n_544), .Z(O0[17]), .CO(n_546));
	notech_ha2 i_16(.A(tsc[16]), .B(n_542), .Z(O0[16]), .CO(n_544));
	notech_ha2 i_15(.A(tsc[15]), .B(n_540), .Z(O0[15]), .CO(n_542));
	notech_ha2 i_14(.A(tsc[14]), .B(n_538), .Z(O0[14]), .CO(n_540));
	notech_ha2 i_13(.A(tsc[13]), .B(n_536), .Z(O0[13]), .CO(n_538));
	notech_ha2 i_12(.A(tsc[12]), .B(n_534), .Z(O0[12]), .CO(n_536));
	notech_ha2 i_11(.A(tsc[11]), .B(n_532), .Z(O0[11]), .CO(n_534));
	notech_ha2 i_10(.A(tsc[10]), .B(n_530), .Z(O0[10]), .CO(n_532));
	notech_ha2 i_9(.A(tsc[9]), .B(n_528), .Z(O0[9]), .CO(n_530));
	notech_ha2 i_8(.A(tsc[8]), .B(n_526), .Z(O0[8]), .CO(n_528));
	notech_ha2 i_7(.A(tsc[7]), .B(n_524), .Z(O0[7]), .CO(n_526));
	notech_ha2 i_6(.A(tsc[6]), .B(n_522), .Z(O0[6]), .CO(n_524));
	notech_ha2 i_5(.A(tsc[5]), .B(n_520), .Z(O0[5]), .CO(n_522));
	notech_ha2 i_4(.A(tsc[4]), .B(n_518), .Z(O0[4]), .CO(n_520));
	notech_ha2 i_3(.A(tsc[3]), .B(n_516), .Z(O0[3]), .CO(n_518));
	notech_ha2 i_2(.A(tsc[2]), .B(n_514), .Z(O0[2]), .CO(n_516));
	notech_ha2 i_1(.A(tsc[1]), .B(tsc[0]), .Z(O0[1]), .CO(n_514));
	notech_inv i_0(.A(tsc[0]), .Z(O0[0]));
endmodule
module AWDP_INC_125(O0, I0);

	output [63:0] O0;
	input [63:0] I0;




	notech_ha2 i_63(.A(I0[63]), .B(n_636), .Z(O0[63]));
	notech_ha2 i_62(.A(I0[62]), .B(n_634), .Z(O0[62]), .CO(n_636));
	notech_ha2 i_61(.A(I0[61]), .B(n_632), .Z(O0[61]), .CO(n_634));
	notech_ha2 i_60(.A(I0[60]), .B(n_630), .Z(O0[60]), .CO(n_632));
	notech_ha2 i_59(.A(I0[59]), .B(n_628), .Z(O0[59]), .CO(n_630));
	notech_ha2 i_58(.A(I0[58]), .B(n_626), .Z(O0[58]), .CO(n_628));
	notech_ha2 i_57(.A(I0[57]), .B(n_624), .Z(O0[57]), .CO(n_626));
	notech_ha2 i_56(.A(I0[56]), .B(n_622), .Z(O0[56]), .CO(n_624));
	notech_ha2 i_55(.A(I0[55]), .B(n_620), .Z(O0[55]), .CO(n_622));
	notech_ha2 i_54(.A(I0[54]), .B(n_618), .Z(O0[54]), .CO(n_620));
	notech_ha2 i_53(.A(I0[53]), .B(n_616), .Z(O0[53]), .CO(n_618));
	notech_ha2 i_52(.A(I0[52]), .B(n_614), .Z(O0[52]), .CO(n_616));
	notech_ha2 i_51(.A(I0[51]), .B(n_612), .Z(O0[51]), .CO(n_614));
	notech_ha2 i_50(.A(I0[50]), .B(n_610), .Z(O0[50]), .CO(n_612));
	notech_ha2 i_49(.A(I0[49]), .B(n_608), .Z(O0[49]), .CO(n_610));
	notech_ha2 i_48(.A(I0[48]), .B(n_606), .Z(O0[48]), .CO(n_608));
	notech_ha2 i_47(.A(I0[47]), .B(n_604), .Z(O0[47]), .CO(n_606));
	notech_ha2 i_46(.A(I0[46]), .B(n_602), .Z(O0[46]), .CO(n_604));
	notech_ha2 i_45(.A(I0[45]), .B(n_600), .Z(O0[45]), .CO(n_602));
	notech_ha2 i_44(.A(I0[44]), .B(n_598), .Z(O0[44]), .CO(n_600));
	notech_ha2 i_43(.A(I0[43]), .B(n_596), .Z(O0[43]), .CO(n_598));
	notech_ha2 i_42(.A(I0[42]), .B(n_594), .Z(O0[42]), .CO(n_596));
	notech_ha2 i_41(.A(I0[41]), .B(n_592), .Z(O0[41]), .CO(n_594));
	notech_ha2 i_40(.A(I0[40]), .B(n_590), .Z(O0[40]), .CO(n_592));
	notech_ha2 i_39(.A(I0[39]), .B(n_588), .Z(O0[39]), .CO(n_590));
	notech_ha2 i_38(.A(I0[38]), .B(n_586), .Z(O0[38]), .CO(n_588));
	notech_ha2 i_37(.A(I0[37]), .B(n_584), .Z(O0[37]), .CO(n_586));
	notech_ha2 i_36(.A(I0[36]), .B(n_582), .Z(O0[36]), .CO(n_584));
	notech_ha2 i_35(.A(I0[35]), .B(n_580), .Z(O0[35]), .CO(n_582));
	notech_ha2 i_34(.A(I0[34]), .B(n_578), .Z(O0[34]), .CO(n_580));
	notech_ha2 i_33(.A(I0[33]), .B(n_576), .Z(O0[33]), .CO(n_578));
	notech_ha2 i_32(.A(I0[32]), .B(n_574), .Z(O0[32]), .CO(n_576));
	notech_ha2 i_31(.A(I0[31]), .B(n_572), .Z(O0[31]), .CO(n_574));
	notech_ha2 i_30(.A(I0[30]), .B(n_570), .Z(O0[30]), .CO(n_572));
	notech_ha2 i_29(.A(I0[29]), .B(n_568), .Z(O0[29]), .CO(n_570));
	notech_ha2 i_28(.A(I0[28]), .B(n_566), .Z(O0[28]), .CO(n_568));
	notech_ha2 i_27(.A(I0[27]), .B(n_564), .Z(O0[27]), .CO(n_566));
	notech_ha2 i_26(.A(I0[26]), .B(n_562), .Z(O0[26]), .CO(n_564));
	notech_ha2 i_25(.A(I0[25]), .B(n_560), .Z(O0[25]), .CO(n_562));
	notech_ha2 i_24(.A(I0[24]), .B(n_558), .Z(O0[24]), .CO(n_560));
	notech_ha2 i_23(.A(I0[23]), .B(n_556), .Z(O0[23]), .CO(n_558));
	notech_ha2 i_22(.A(I0[22]), .B(n_554), .Z(O0[22]), .CO(n_556));
	notech_ha2 i_21(.A(I0[21]), .B(n_552), .Z(O0[21]), .CO(n_554));
	notech_ha2 i_20(.A(I0[20]), .B(n_550), .Z(O0[20]), .CO(n_552));
	notech_ha2 i_19(.A(I0[19]), .B(n_548), .Z(O0[19]), .CO(n_550));
	notech_ha2 i_18(.A(I0[18]), .B(n_546), .Z(O0[18]), .CO(n_548));
	notech_ha2 i_17(.A(I0[17]), .B(n_544), .Z(O0[17]), .CO(n_546));
	notech_ha2 i_16(.A(I0[16]), .B(n_542), .Z(O0[16]), .CO(n_544));
	notech_ha2 i_15(.A(I0[15]), .B(n_540), .Z(O0[15]), .CO(n_542));
	notech_ha2 i_14(.A(I0[14]), .B(n_538), .Z(O0[14]), .CO(n_540));
	notech_ha2 i_13(.A(I0[13]), .B(n_536), .Z(O0[13]), .CO(n_538));
	notech_ha2 i_12(.A(I0[12]), .B(n_534), .Z(O0[12]), .CO(n_536));
	notech_ha2 i_11(.A(I0[11]), .B(n_532), .Z(O0[11]), .CO(n_534));
	notech_ha2 i_10(.A(I0[10]), .B(n_530), .Z(O0[10]), .CO(n_532));
	notech_ha2 i_9(.A(I0[9]), .B(n_528), .Z(O0[9]), .CO(n_530));
	notech_ha2 i_8(.A(I0[8]), .B(n_526), .Z(O0[8]), .CO(n_528));
	notech_ha2 i_7(.A(I0[7]), .B(n_524), .Z(O0[7]), .CO(n_526));
	notech_ha2 i_6(.A(I0[6]), .B(n_522), .Z(O0[6]), .CO(n_524));
	notech_ha2 i_5(.A(I0[5]), .B(n_520), .Z(O0[5]), .CO(n_522));
	notech_ha2 i_4(.A(I0[4]), .B(n_518), .Z(O0[4]), .CO(n_520));
	notech_ha2 i_3(.A(I0[3]), .B(n_516), .Z(O0[3]), .CO(n_518));
	notech_ha2 i_2(.A(I0[2]), .B(n_514), .Z(O0[2]), .CO(n_516));
	notech_ha2 i_1(.A(I0[0]), .B(I0[1]), .Z(O0[1]), .CO(n_514));
	notech_inv i_0(.A(I0[0]), .Z(O0[0]));
endmodule
module AWDP_INC_153(O0, I0);

	output [31:0] O0;
	input [31:0] I0;




	notech_ha2 i_31(.A(I0[31]), .B(n_316), .Z(O0[31]));
	notech_ha2 i_30(.A(I0[30]), .B(n_314), .Z(O0[30]), .CO(n_316));
	notech_ha2 i_29(.A(I0[29]), .B(n_312), .Z(O0[29]), .CO(n_314));
	notech_ha2 i_28(.A(I0[28]), .B(n_310), .Z(O0[28]), .CO(n_312));
	notech_ha2 i_27(.A(I0[27]), .B(n_308), .Z(O0[27]), .CO(n_310));
	notech_ha2 i_26(.A(I0[26]), .B(n_306), .Z(O0[26]), .CO(n_308));
	notech_ha2 i_25(.A(I0[25]), .B(n_304), .Z(O0[25]), .CO(n_306));
	notech_ha2 i_24(.A(I0[24]), .B(n_302), .Z(O0[24]), .CO(n_304));
	notech_ha2 i_23(.A(I0[23]), .B(n_300), .Z(O0[23]), .CO(n_302));
	notech_ha2 i_22(.A(I0[22]), .B(n_298), .Z(O0[22]), .CO(n_300));
	notech_ha2 i_21(.A(I0[21]), .B(n_296), .Z(O0[21]), .CO(n_298));
	notech_ha2 i_20(.A(I0[20]), .B(n_294), .Z(O0[20]), .CO(n_296));
	notech_ha2 i_19(.A(I0[19]), .B(n_292), .Z(O0[19]), .CO(n_294));
	notech_ha2 i_18(.A(I0[18]), .B(n_290), .Z(O0[18]), .CO(n_292));
	notech_ha2 i_17(.A(I0[17]), .B(n_288), .Z(O0[17]), .CO(n_290));
	notech_ha2 i_16(.A(I0[16]), .B(n_286), .Z(O0[16]), .CO(n_288));
	notech_ha2 i_15(.A(I0[15]), .B(n_284), .Z(O0[15]), .CO(n_286));
	notech_ha2 i_14(.A(I0[14]), .B(n_282), .Z(O0[14]), .CO(n_284));
	notech_ha2 i_13(.A(I0[13]), .B(n_280), .Z(O0[13]), .CO(n_282));
	notech_ha2 i_12(.A(I0[12]), .B(n_278), .Z(O0[12]), .CO(n_280));
	notech_ha2 i_11(.A(I0[11]), .B(n_276), .Z(O0[11]), .CO(n_278));
	notech_ha2 i_10(.A(I0[10]), .B(n_274), .Z(O0[10]), .CO(n_276));
	notech_ha2 i_9(.A(I0[9]), .B(n_272), .Z(O0[9]), .CO(n_274));
	notech_ha2 i_8(.A(I0[8]), .B(n_270), .Z(O0[8]), .CO(n_272));
	notech_ha2 i_7(.A(I0[7]), .B(n_268), .Z(O0[7]), .CO(n_270));
	notech_ha2 i_6(.A(I0[6]), .B(n_266), .Z(O0[6]), .CO(n_268));
	notech_ha2 i_5(.A(I0[5]), .B(n_264), .Z(O0[5]), .CO(n_266));
	notech_ha2 i_4(.A(I0[4]), .B(n_262), .Z(O0[4]), .CO(n_264));
	notech_ha2 i_3(.A(I0[3]), .B(n_260), .Z(O0[3]), .CO(n_262));
	notech_ha2 i_2(.A(I0[2]), .B(n_258), .Z(O0[2]), .CO(n_260));
	notech_ha2 i_1(.A(I0[0]), .B(I0[1]), .Z(O0[1]), .CO(n_258));
	notech_inv i_0(.A(I0[0]), .Z(O0[0]));
endmodule
module AWDP_INC_163(O0, I0);

	output [63:0] O0;
	input [63:0] I0;




	notech_ha2 i_31(.A(I0[31]), .B(n_573), .Z(O0[31]), .CO(O0[32]));
	notech_ha2 i_30(.A(I0[30]), .B(n_571), .Z(O0[30]), .CO(n_573));
	notech_ha2 i_29(.A(I0[29]), .B(n_569), .Z(O0[29]), .CO(n_571));
	notech_ha2 i_28(.A(I0[28]), .B(n_567), .Z(O0[28]), .CO(n_569));
	notech_ha2 i_27(.A(I0[27]), .B(n_565), .Z(O0[27]), .CO(n_567));
	notech_ha2 i_26(.A(I0[26]), .B(n_563), .Z(O0[26]), .CO(n_565));
	notech_ha2 i_25(.A(I0[25]), .B(n_561), .Z(O0[25]), .CO(n_563));
	notech_ha2 i_24(.A(I0[24]), .B(n_559), .Z(O0[24]), .CO(n_561));
	notech_ha2 i_23(.A(I0[23]), .B(n_557), .Z(O0[23]), .CO(n_559));
	notech_ha2 i_22(.A(I0[22]), .B(n_555), .Z(O0[22]), .CO(n_557));
	notech_ha2 i_21(.A(I0[21]), .B(n_553), .Z(O0[21]), .CO(n_555));
	notech_ha2 i_20(.A(I0[20]), .B(n_551), .Z(O0[20]), .CO(n_553));
	notech_ha2 i_19(.A(I0[19]), .B(n_549), .Z(O0[19]), .CO(n_551));
	notech_ha2 i_18(.A(I0[18]), .B(n_547), .Z(O0[18]), .CO(n_549));
	notech_ha2 i_17(.A(I0[17]), .B(n_545), .Z(O0[17]), .CO(n_547));
	notech_ha2 i_16(.A(I0[16]), .B(n_543), .Z(O0[16]), .CO(n_545));
	notech_ha2 i_15(.A(I0[15]), .B(n_541), .Z(O0[15]), .CO(n_543));
	notech_ha2 i_14(.A(I0[14]), .B(n_539), .Z(O0[14]), .CO(n_541));
	notech_ha2 i_13(.A(I0[13]), .B(n_537), .Z(O0[13]), .CO(n_539));
	notech_ha2 i_12(.A(I0[12]), .B(n_535), .Z(O0[12]), .CO(n_537));
	notech_ha2 i_11(.A(I0[11]), .B(n_533), .Z(O0[11]), .CO(n_535));
	notech_ha2 i_10(.A(I0[10]), .B(n_531), .Z(O0[10]), .CO(n_533));
	notech_ha2 i_9(.A(I0[9]), .B(n_529), .Z(O0[9]), .CO(n_531));
	notech_ha2 i_8(.A(I0[8]), .B(n_527), .Z(O0[8]), .CO(n_529));
	notech_ha2 i_7(.A(I0[7]), .B(n_525), .Z(O0[7]), .CO(n_527));
	notech_ha2 i_6(.A(I0[6]), .B(n_523), .Z(O0[6]), .CO(n_525));
	notech_ha2 i_5(.A(I0[5]), .B(n_521), .Z(O0[5]), .CO(n_523));
	notech_ha2 i_4(.A(I0[4]), .B(n_519), .Z(O0[4]), .CO(n_521));
	notech_ha2 i_3(.A(I0[3]), .B(n_517), .Z(O0[3]), .CO(n_519));
	notech_ha2 i_2(.A(I0[2]), .B(n_515), .Z(O0[2]), .CO(n_517));
	notech_ha2 i_1(.A(I0[0]), .B(I0[1]), .Z(O0[1]), .CO(n_515));
	notech_inv i_0(.A(I0[0]), .Z(O0[0]));
endmodule
module AWDP_INC_200(O0, I0);

	output [31:0] O0;
	input [31:0] I0;




	notech_ha2 i_31(.A(I0[31]), .B(n_316), .Z(O0[31]));
	notech_ha2 i_30(.A(I0[30]), .B(n_314), .Z(O0[30]), .CO(n_316));
	notech_ha2 i_29(.A(I0[29]), .B(n_312), .Z(O0[29]), .CO(n_314));
	notech_ha2 i_28(.A(I0[28]), .B(n_310), .Z(O0[28]), .CO(n_312));
	notech_ha2 i_27(.A(I0[27]), .B(n_308), .Z(O0[27]), .CO(n_310));
	notech_ha2 i_26(.A(I0[26]), .B(n_306), .Z(O0[26]), .CO(n_308));
	notech_ha2 i_25(.A(I0[25]), .B(n_304), .Z(O0[25]), .CO(n_306));
	notech_ha2 i_24(.A(I0[24]), .B(n_302), .Z(O0[24]), .CO(n_304));
	notech_ha2 i_23(.A(I0[23]), .B(n_300), .Z(O0[23]), .CO(n_302));
	notech_ha2 i_22(.A(I0[22]), .B(n_298), .Z(O0[22]), .CO(n_300));
	notech_ha2 i_21(.A(I0[21]), .B(n_296), .Z(O0[21]), .CO(n_298));
	notech_ha2 i_20(.A(I0[20]), .B(n_294), .Z(O0[20]), .CO(n_296));
	notech_ha2 i_19(.A(I0[19]), .B(n_292), .Z(O0[19]), .CO(n_294));
	notech_ha2 i_18(.A(I0[18]), .B(n_290), .Z(O0[18]), .CO(n_292));
	notech_ha2 i_17(.A(I0[17]), .B(n_288), .Z(O0[17]), .CO(n_290));
	notech_ha2 i_16(.A(I0[16]), .B(n_286), .Z(O0[16]), .CO(n_288));
	notech_ha2 i_15(.A(I0[15]), .B(n_284), .Z(O0[15]), .CO(n_286));
	notech_ha2 i_14(.A(I0[14]), .B(n_282), .Z(O0[14]), .CO(n_284));
	notech_ha2 i_13(.A(I0[13]), .B(n_280), .Z(O0[13]), .CO(n_282));
	notech_ha2 i_12(.A(I0[12]), .B(n_278), .Z(O0[12]), .CO(n_280));
	notech_ha2 i_11(.A(I0[11]), .B(n_276), .Z(O0[11]), .CO(n_278));
	notech_ha2 i_10(.A(I0[10]), .B(n_274), .Z(O0[10]), .CO(n_276));
	notech_ha2 i_9(.A(I0[9]), .B(n_272), .Z(O0[9]), .CO(n_274));
	notech_ha2 i_8(.A(I0[8]), .B(n_270), .Z(O0[8]), .CO(n_272));
	notech_ha2 i_7(.A(I0[7]), .B(n_268), .Z(O0[7]), .CO(n_270));
	notech_ha2 i_6(.A(I0[6]), .B(n_266), .Z(O0[6]), .CO(n_268));
	notech_ha2 i_5(.A(I0[5]), .B(n_264), .Z(O0[5]), .CO(n_266));
	notech_ha2 i_4(.A(I0[4]), .B(n_262), .Z(O0[4]), .CO(n_264));
	notech_ha2 i_3(.A(I0[3]), .B(n_260), .Z(O0[3]), .CO(n_262));
	notech_ha2 i_2(.A(I0[2]), .B(n_258), .Z(O0[2]), .CO(n_260));
	notech_ha2 i_1(.A(I0[1]), .B(I0[0]), .Z(O0[1]), .CO(n_258));
	notech_inv i_0(.A(I0[0]), .Z(O0[0]));
endmodule
module AWDP_INC_210(O0, I0);

	output [31:0] O0;
	input [31:0] I0;




	notech_ha2 i_31(.A(I0[31]), .B(n_316), .Z(O0[31]));
	notech_ha2 i_30(.A(I0[30]), .B(n_314), .Z(O0[30]), .CO(n_316));
	notech_ha2 i_29(.A(I0[29]), .B(n_312), .Z(O0[29]), .CO(n_314));
	notech_ha2 i_28(.A(I0[28]), .B(n_310), .Z(O0[28]), .CO(n_312));
	notech_ha2 i_27(.A(I0[27]), .B(n_308), .Z(O0[27]), .CO(n_310));
	notech_ha2 i_26(.A(I0[26]), .B(n_306), .Z(O0[26]), .CO(n_308));
	notech_ha2 i_25(.A(I0[25]), .B(n_304), .Z(O0[25]), .CO(n_306));
	notech_ha2 i_24(.A(I0[24]), .B(n_302), .Z(O0[24]), .CO(n_304));
	notech_ha2 i_23(.A(I0[23]), .B(n_300), .Z(O0[23]), .CO(n_302));
	notech_ha2 i_22(.A(I0[22]), .B(n_298), .Z(O0[22]), .CO(n_300));
	notech_ha2 i_21(.A(I0[21]), .B(n_296), .Z(O0[21]), .CO(n_298));
	notech_ha2 i_20(.A(I0[20]), .B(n_294), .Z(O0[20]), .CO(n_296));
	notech_ha2 i_19(.A(I0[19]), .B(n_292), .Z(O0[19]), .CO(n_294));
	notech_ha2 i_18(.A(I0[18]), .B(n_290), .Z(O0[18]), .CO(n_292));
	notech_ha2 i_17(.A(I0[17]), .B(n_288), .Z(O0[17]), .CO(n_290));
	notech_ha2 i_16(.A(I0[16]), .B(n_286), .Z(O0[16]), .CO(n_288));
	notech_ha2 i_15(.A(I0[15]), .B(n_284), .Z(O0[15]), .CO(n_286));
	notech_ha2 i_14(.A(I0[14]), .B(n_282), .Z(O0[14]), .CO(n_284));
	notech_ha2 i_13(.A(I0[13]), .B(n_280), .Z(O0[13]), .CO(n_282));
	notech_ha2 i_12(.A(I0[12]), .B(n_278), .Z(O0[12]), .CO(n_280));
	notech_ha2 i_11(.A(I0[11]), .B(n_276), .Z(O0[11]), .CO(n_278));
	notech_ha2 i_10(.A(I0[10]), .B(n_274), .Z(O0[10]), .CO(n_276));
	notech_ha2 i_9(.A(I0[9]), .B(n_272), .Z(O0[9]), .CO(n_274));
	notech_ha2 i_8(.A(I0[8]), .B(n_270), .Z(O0[8]), .CO(n_272));
	notech_ha2 i_7(.A(I0[7]), .B(n_268), .Z(O0[7]), .CO(n_270));
	notech_ha2 i_6(.A(I0[6]), .B(n_266), .Z(O0[6]), .CO(n_268));
	notech_ha2 i_5(.A(I0[5]), .B(n_264), .Z(O0[5]), .CO(n_266));
	notech_ha2 i_4(.A(I0[4]), .B(n_262), .Z(O0[4]), .CO(n_264));
	notech_ha2 i_3(.A(I0[3]), .B(n_260), .Z(O0[3]), .CO(n_262));
	notech_ha2 i_2(.A(I0[2]), .B(n_258), .Z(O0[2]), .CO(n_260));
	notech_ha2 i_1(.A(I0[1]), .B(I0[0]), .Z(O0[1]), .CO(n_258));
	notech_inv i_0(.A(I0[0]), .Z(O0[0]));
endmodule
module AWDP_INC_26111934(O0, I0);

	output [15:0] O0;
	input [15:0] I0;




	notech_ha2 i_15(.A(I0[15]), .B(n_156), .Z(O0[15]));
	notech_ha2 i_14(.A(I0[14]), .B(n_154), .Z(O0[14]), .CO(n_156));
	notech_ha2 i_13(.A(I0[13]), .B(n_152), .Z(O0[13]), .CO(n_154));
	notech_ha2 i_12(.A(I0[12]), .B(n_150), .Z(O0[12]), .CO(n_152));
	notech_ha2 i_11(.A(I0[11]), .B(n_148), .Z(O0[11]), .CO(n_150));
	notech_ha2 i_10(.A(I0[10]), .B(n_146), .Z(O0[10]), .CO(n_148));
	notech_ha2 i_9(.A(I0[9]), .B(n_144), .Z(O0[9]), .CO(n_146));
	notech_ha2 i_8(.A(I0[8]), .B(n_142), .Z(O0[8]), .CO(n_144));
	notech_ha2 i_7(.A(I0[7]), .B(n_140), .Z(O0[7]), .CO(n_142));
	notech_ha2 i_6(.A(I0[6]), .B(n_138), .Z(O0[6]), .CO(n_140));
	notech_ha2 i_5(.A(I0[5]), .B(n_136), .Z(O0[5]), .CO(n_138));
	notech_ha2 i_4(.A(I0[4]), .B(n_134), .Z(O0[4]), .CO(n_136));
	notech_ha2 i_3(.A(I0[3]), .B(n_132), .Z(O0[3]), .CO(n_134));
	notech_ha2 i_2(.A(I0[2]), .B(n_130), .Z(O0[2]), .CO(n_132));
	notech_ha2 i_1(.A(I0[0]), .B(I0[1]), .Z(O0[1]), .CO(n_130));
	notech_inv i_0(.A(I0[0]), .Z(O0[0]));
endmodule
module AWDP_LE_211(O0, divq, I0);

	output [0:0] O0;
	input [63:0] divq;
	input [63:0] I0;




	notech_inv i_320(.A(n_710), .Z(O0[0]));
	notech_nand2 i_317(.A(n_703), .B(n_709), .Z(n_710));
	notech_inv i_506(.A(n_835), .Z(n_703));
	notech_or2 i_505(.A(n_834), .B(n_701), .Z(n_835));
	notech_and2 i_504(.A(n_702), .B(n_700), .Z(n_834));
	notech_inv i_315(.A(n_512), .Z(n_702));
	notech_inv i_314(.A(n_577), .Z(n_701));
	notech_inv i_503(.A(n_928), .Z(n_700));
	notech_nor2 i_502(.A(n_927), .B(n_866), .Z(n_928));
	notech_nor2 i_501(.A(n_699), .B(n_511), .Z(n_927));
	notech_inv i_500(.A(n_831), .Z(n_699));
	notech_or2 i_499(.A(n_830), .B(n_697), .Z(n_831));
	notech_and2 i_498(.A(n_698), .B(n_696), .Z(n_830));
	notech_inv i_311(.A(n_510), .Z(n_698));
	notech_inv i_310(.A(n_575), .Z(n_697));
	notech_inv i_497(.A(n_926), .Z(n_696));
	notech_nor2 i_496(.A(n_925), .B(n_865), .Z(n_926));
	notech_nor2 i_495(.A(n_695), .B(n_509), .Z(n_925));
	notech_inv i_494(.A(n_827), .Z(n_695));
	notech_or2 i_493(.A(n_826), .B(n_693), .Z(n_827));
	notech_and2 i_492(.A(n_694), .B(n_692), .Z(n_826));
	notech_inv i_307(.A(n_508), .Z(n_694));
	notech_inv i_306(.A(n_573), .Z(n_693));
	notech_inv i_491(.A(n_924), .Z(n_692));
	notech_nor2 i_490(.A(n_923), .B(n_864), .Z(n_924));
	notech_nor2 i_489(.A(n_691), .B(n_507), .Z(n_923));
	notech_inv i_488(.A(n_823), .Z(n_691));
	notech_or2 i_487(.A(n_822), .B(n_689), .Z(n_823));
	notech_and2 i_486(.A(n_690), .B(n_688), .Z(n_822));
	notech_inv i_303(.A(n_506), .Z(n_690));
	notech_inv i_302(.A(n_571), .Z(n_689));
	notech_inv i_485(.A(n_922), .Z(n_688));
	notech_nor2 i_484(.A(n_921), .B(n_863), .Z(n_922));
	notech_nor2 i_483(.A(n_687), .B(n_505), .Z(n_921));
	notech_inv i_482(.A(n_819), .Z(n_687));
	notech_or2 i_481(.A(n_818), .B(n_685), .Z(n_819));
	notech_and2 i_480(.A(n_686), .B(n_684), .Z(n_818));
	notech_inv i_299(.A(n_504), .Z(n_686));
	notech_inv i_298(.A(n_569), .Z(n_685));
	notech_inv i_479(.A(n_920), .Z(n_684));
	notech_nor2 i_478(.A(n_919), .B(n_862), .Z(n_920));
	notech_nor2 i_477(.A(n_683), .B(n_503), .Z(n_919));
	notech_inv i_476(.A(n_815), .Z(n_683));
	notech_or2 i_475(.A(n_814), .B(n_681), .Z(n_815));
	notech_and2 i_474(.A(n_682), .B(n_680), .Z(n_814));
	notech_inv i_295(.A(n_502), .Z(n_682));
	notech_inv i_294(.A(n_567), .Z(n_681));
	notech_inv i_473(.A(n_918), .Z(n_680));
	notech_nor2 i_472(.A(n_917), .B(n_861), .Z(n_918));
	notech_nor2 i_471(.A(n_679), .B(n_501), .Z(n_917));
	notech_inv i_470(.A(n_811), .Z(n_679));
	notech_or2 i_469(.A(n_810), .B(n_677), .Z(n_811));
	notech_and2 i_468(.A(n_678), .B(n_676), .Z(n_810));
	notech_inv i_291(.A(n_500), .Z(n_678));
	notech_inv i_290(.A(n_565), .Z(n_677));
	notech_inv i_467(.A(n_916), .Z(n_676));
	notech_nor2 i_466(.A(n_915), .B(n_860), .Z(n_916));
	notech_nor2 i_465(.A(n_675), .B(n_499), .Z(n_915));
	notech_inv i_464(.A(n_807), .Z(n_675));
	notech_or2 i_463(.A(n_806), .B(n_673), .Z(n_807));
	notech_and2 i_462(.A(n_674), .B(n_672), .Z(n_806));
	notech_inv i_287(.A(n_498), .Z(n_674));
	notech_inv i_286(.A(n_563), .Z(n_673));
	notech_inv i_461(.A(n_914), .Z(n_672));
	notech_nor2 i_460(.A(n_913), .B(n_859), .Z(n_914));
	notech_nor2 i_459(.A(n_671), .B(n_497), .Z(n_913));
	notech_inv i_458(.A(n_803), .Z(n_671));
	notech_or2 i_457(.A(n_802), .B(n_669), .Z(n_803));
	notech_and2 i_456(.A(n_670), .B(n_668), .Z(n_802));
	notech_inv i_283(.A(n_496), .Z(n_670));
	notech_inv i_282(.A(n_561), .Z(n_669));
	notech_inv i_455(.A(n_912), .Z(n_668));
	notech_nor2 i_454(.A(n_911), .B(n_858), .Z(n_912));
	notech_nor2 i_453(.A(n_667), .B(n_495), .Z(n_911));
	notech_inv i_452(.A(n_799), .Z(n_667));
	notech_or2 i_451(.A(n_798), .B(n_665), .Z(n_799));
	notech_and2 i_450(.A(n_666), .B(n_664), .Z(n_798));
	notech_inv i_279(.A(n_494), .Z(n_666));
	notech_inv i_278(.A(n_559), .Z(n_665));
	notech_inv i_449(.A(n_910), .Z(n_664));
	notech_nor2 i_448(.A(n_909), .B(n_857), .Z(n_910));
	notech_nor2 i_447(.A(n_663), .B(n_493), .Z(n_909));
	notech_inv i_446(.A(n_795), .Z(n_663));
	notech_or2 i_445(.A(n_794), .B(n_661), .Z(n_795));
	notech_and2 i_444(.A(n_662), .B(n_660), .Z(n_794));
	notech_inv i_275(.A(n_492), .Z(n_662));
	notech_inv i_274(.A(n_557), .Z(n_661));
	notech_inv i_443(.A(n_908), .Z(n_660));
	notech_nor2 i_442(.A(n_907), .B(n_856), .Z(n_908));
	notech_nor2 i_441(.A(n_659), .B(n_491), .Z(n_907));
	notech_inv i_440(.A(n_791), .Z(n_659));
	notech_or2 i_439(.A(n_790), .B(n_657), .Z(n_791));
	notech_and2 i_438(.A(n_658), .B(n_656), .Z(n_790));
	notech_inv i_271(.A(n_490), .Z(n_658));
	notech_inv i_270(.A(n_555), .Z(n_657));
	notech_inv i_437(.A(n_906), .Z(n_656));
	notech_nor2 i_436(.A(n_905), .B(n_855), .Z(n_906));
	notech_nor2 i_435(.A(n_655), .B(n_489), .Z(n_905));
	notech_inv i_434(.A(n_787), .Z(n_655));
	notech_or2 i_433(.A(n_786), .B(n_653), .Z(n_787));
	notech_and2 i_432(.A(n_654), .B(n_652), .Z(n_786));
	notech_inv i_267(.A(n_488), .Z(n_654));
	notech_inv i_266(.A(n_553), .Z(n_653));
	notech_inv i_431(.A(n_904), .Z(n_652));
	notech_nor2 i_430(.A(n_903), .B(n_854), .Z(n_904));
	notech_nor2 i_429(.A(n_651), .B(n_487), .Z(n_903));
	notech_inv i_428(.A(n_783), .Z(n_651));
	notech_or2 i_427(.A(n_782), .B(n_649), .Z(n_783));
	notech_and2 i_426(.A(n_650), .B(n_648), .Z(n_782));
	notech_inv i_263(.A(n_486), .Z(n_650));
	notech_inv i_262(.A(n_551), .Z(n_649));
	notech_inv i_425(.A(n_902), .Z(n_648));
	notech_nor2 i_424(.A(n_901), .B(n_853), .Z(n_902));
	notech_nor2 i_423(.A(n_647), .B(n_485), .Z(n_901));
	notech_inv i_422(.A(n_779), .Z(n_647));
	notech_or2 i_421(.A(n_778), .B(n_645), .Z(n_779));
	notech_and2 i_420(.A(n_646), .B(n_644), .Z(n_778));
	notech_inv i_259(.A(n_484), .Z(n_646));
	notech_inv i_258(.A(n_549), .Z(n_645));
	notech_inv i_419(.A(n_900), .Z(n_644));
	notech_nor2 i_418(.A(n_899), .B(n_852), .Z(n_900));
	notech_nor2 i_417(.A(n_643), .B(n_483), .Z(n_899));
	notech_inv i_416(.A(n_775), .Z(n_643));
	notech_or2 i_415(.A(n_774), .B(n_641), .Z(n_775));
	notech_and2 i_414(.A(n_642), .B(n_640), .Z(n_774));
	notech_inv i_255(.A(n_482), .Z(n_642));
	notech_inv i_254(.A(n_547), .Z(n_641));
	notech_inv i_413(.A(n_898), .Z(n_640));
	notech_nor2 i_412(.A(n_897), .B(n_851), .Z(n_898));
	notech_nor2 i_411(.A(n_639), .B(n_481), .Z(n_897));
	notech_inv i_410(.A(n_771), .Z(n_639));
	notech_or2 i_409(.A(n_770), .B(n_637), .Z(n_771));
	notech_and2 i_408(.A(n_638), .B(n_636), .Z(n_770));
	notech_inv i_251(.A(n_480), .Z(n_638));
	notech_inv i_250(.A(n_545), .Z(n_637));
	notech_inv i_407(.A(n_896), .Z(n_636));
	notech_nor2 i_406(.A(n_895), .B(n_850), .Z(n_896));
	notech_nor2 i_405(.A(n_635), .B(n_479), .Z(n_895));
	notech_inv i_404(.A(n_767), .Z(n_635));
	notech_or2 i_403(.A(n_766), .B(n_633), .Z(n_767));
	notech_and2 i_402(.A(n_634), .B(n_632), .Z(n_766));
	notech_inv i_247(.A(n_478), .Z(n_634));
	notech_inv i_246(.A(n_543), .Z(n_633));
	notech_inv i_401(.A(n_894), .Z(n_632));
	notech_nor2 i_400(.A(n_893), .B(n_849), .Z(n_894));
	notech_nor2 i_399(.A(n_631), .B(n_477), .Z(n_893));
	notech_inv i_398(.A(n_763), .Z(n_631));
	notech_or2 i_397(.A(n_762), .B(n_629), .Z(n_763));
	notech_and2 i_396(.A(n_630), .B(n_628), .Z(n_762));
	notech_inv i_243(.A(n_476), .Z(n_630));
	notech_inv i_242(.A(n_541), .Z(n_629));
	notech_inv i_395(.A(n_892), .Z(n_628));
	notech_nor2 i_394(.A(n_891), .B(n_848), .Z(n_892));
	notech_nor2 i_393(.A(n_627), .B(n_475), .Z(n_891));
	notech_inv i_392(.A(n_759), .Z(n_627));
	notech_or2 i_391(.A(n_758), .B(n_625), .Z(n_759));
	notech_and2 i_390(.A(n_626), .B(n_624), .Z(n_758));
	notech_inv i_239(.A(n_474), .Z(n_626));
	notech_inv i_238(.A(n_539), .Z(n_625));
	notech_inv i_389(.A(n_890), .Z(n_624));
	notech_nor2 i_388(.A(n_889), .B(n_847), .Z(n_890));
	notech_nor2 i_387(.A(n_623), .B(n_473), .Z(n_889));
	notech_inv i_386(.A(n_755), .Z(n_623));
	notech_or2 i_385(.A(n_754), .B(n_621), .Z(n_755));
	notech_and2 i_384(.A(n_622), .B(n_620), .Z(n_754));
	notech_inv i_235(.A(n_472), .Z(n_622));
	notech_inv i_234(.A(n_537), .Z(n_621));
	notech_inv i_383(.A(n_888), .Z(n_620));
	notech_nor2 i_382(.A(n_887), .B(n_846), .Z(n_888));
	notech_nor2 i_381(.A(n_619), .B(n_471), .Z(n_887));
	notech_inv i_380(.A(n_751), .Z(n_619));
	notech_or2 i_379(.A(n_750), .B(n_617), .Z(n_751));
	notech_and2 i_378(.A(n_618), .B(n_616), .Z(n_750));
	notech_inv i_231(.A(n_470), .Z(n_618));
	notech_inv i_230(.A(n_535), .Z(n_617));
	notech_inv i_377(.A(n_886), .Z(n_616));
	notech_nor2 i_376(.A(n_885), .B(n_845), .Z(n_886));
	notech_nor2 i_375(.A(n_615), .B(n_469), .Z(n_885));
	notech_inv i_374(.A(n_747), .Z(n_615));
	notech_or2 i_373(.A(n_746), .B(n_613), .Z(n_747));
	notech_and2 i_372(.A(n_614), .B(n_612), .Z(n_746));
	notech_inv i_227(.A(n_468), .Z(n_614));
	notech_inv i_226(.A(n_533), .Z(n_613));
	notech_inv i_371(.A(n_884), .Z(n_612));
	notech_nor2 i_370(.A(n_883), .B(n_844), .Z(n_884));
	notech_nor2 i_369(.A(n_611), .B(n_467), .Z(n_883));
	notech_inv i_368(.A(n_743), .Z(n_611));
	notech_or2 i_367(.A(n_742), .B(n_609), .Z(n_743));
	notech_and2 i_366(.A(n_610), .B(n_608), .Z(n_742));
	notech_inv i_223(.A(n_466), .Z(n_610));
	notech_inv i_222(.A(n_531), .Z(n_609));
	notech_inv i_365(.A(n_882), .Z(n_608));
	notech_nor2 i_364(.A(n_881), .B(n_843), .Z(n_882));
	notech_nor2 i_363(.A(n_607), .B(n_465), .Z(n_881));
	notech_inv i_362(.A(n_739), .Z(n_607));
	notech_or2 i_361(.A(n_738), .B(n_605), .Z(n_739));
	notech_and2 i_360(.A(n_606), .B(n_604), .Z(n_738));
	notech_inv i_219(.A(n_464), .Z(n_606));
	notech_inv i_218(.A(n_529), .Z(n_605));
	notech_inv i_359(.A(n_880), .Z(n_604));
	notech_nor2 i_358(.A(n_879), .B(n_842), .Z(n_880));
	notech_nor2 i_357(.A(n_603), .B(n_463), .Z(n_879));
	notech_inv i_356(.A(n_735), .Z(n_603));
	notech_or2 i_355(.A(n_734), .B(n_601), .Z(n_735));
	notech_and2 i_354(.A(n_602), .B(n_600), .Z(n_734));
	notech_inv i_215(.A(n_462), .Z(n_602));
	notech_inv i_214(.A(n_527), .Z(n_601));
	notech_inv i_353(.A(n_878), .Z(n_600));
	notech_nor2 i_352(.A(n_877), .B(n_841), .Z(n_878));
	notech_nor2 i_351(.A(n_599), .B(n_461), .Z(n_877));
	notech_inv i_350(.A(n_731), .Z(n_599));
	notech_or2 i_349(.A(n_730), .B(n_597), .Z(n_731));
	notech_and2 i_348(.A(n_598), .B(n_596), .Z(n_730));
	notech_inv i_211(.A(n_460), .Z(n_598));
	notech_inv i_210(.A(n_525), .Z(n_597));
	notech_inv i_347(.A(n_876), .Z(n_596));
	notech_nor2 i_346(.A(n_875), .B(n_840), .Z(n_876));
	notech_nor2 i_345(.A(n_595), .B(n_459), .Z(n_875));
	notech_inv i_344(.A(n_727), .Z(n_595));
	notech_or2 i_343(.A(n_726), .B(n_593), .Z(n_727));
	notech_and2 i_342(.A(n_594), .B(n_592), .Z(n_726));
	notech_inv i_207(.A(n_458), .Z(n_594));
	notech_inv i_206(.A(n_523), .Z(n_593));
	notech_inv i_341(.A(n_874), .Z(n_592));
	notech_nor2 i_340(.A(n_873), .B(n_839), .Z(n_874));
	notech_nor2 i_339(.A(n_591), .B(n_457), .Z(n_873));
	notech_inv i_338(.A(n_723), .Z(n_591));
	notech_or2 i_337(.A(n_722), .B(n_589), .Z(n_723));
	notech_and2 i_336(.A(n_590), .B(n_588), .Z(n_722));
	notech_inv i_203(.A(n_456), .Z(n_590));
	notech_inv i_202(.A(n_521), .Z(n_589));
	notech_inv i_335(.A(n_872), .Z(n_588));
	notech_nor2 i_334(.A(n_871), .B(n_838), .Z(n_872));
	notech_nor2 i_333(.A(n_587), .B(n_455), .Z(n_871));
	notech_inv i_332(.A(n_719), .Z(n_587));
	notech_or2 i_331(.A(n_718), .B(n_585), .Z(n_719));
	notech_and2 i_330(.A(n_586), .B(n_584), .Z(n_718));
	notech_inv i_199(.A(n_454), .Z(n_586));
	notech_inv i_198(.A(n_519), .Z(n_585));
	notech_inv i_329(.A(n_870), .Z(n_584));
	notech_nor2 i_328(.A(n_869), .B(n_837), .Z(n_870));
	notech_nor2 i_327(.A(n_583), .B(n_453), .Z(n_869));
	notech_inv i_326(.A(n_715), .Z(n_583));
	notech_or2 i_325(.A(n_714), .B(n_581), .Z(n_715));
	notech_and2 i_324(.A(n_582), .B(n_580), .Z(n_714));
	notech_inv i_195(.A(n_452), .Z(n_582));
	notech_inv i_194(.A(n_517), .Z(n_581));
	notech_inv i_323(.A(n_868), .Z(n_580));
	notech_nor2 i_322(.A(n_867), .B(n_836), .Z(n_868));
	notech_nor2 i_321(.A(n_451), .B(n_515), .Z(n_867));
	notech_inv i_191(.A(divq[63]), .Z(n_709));
	notech_nand2 i_190(.A(n_449), .B(divq[62]), .Z(n_577));
	notech_and2 i_189(.A(n_448), .B(divq[61]), .Z(n_866));
	notech_nand2 i_188(.A(n_447), .B(divq[60]), .Z(n_575));
	notech_and2 i_187(.A(n_446), .B(divq[59]), .Z(n_865));
	notech_nand2 i_186(.A(n_445), .B(divq[58]), .Z(n_573));
	notech_and2 i_185(.A(n_444), .B(divq[57]), .Z(n_864));
	notech_nand2 i_184(.A(n_443), .B(divq[56]), .Z(n_571));
	notech_and2 i_183(.A(n_442), .B(divq[55]), .Z(n_863));
	notech_nand2 i_182(.A(n_441), .B(divq[54]), .Z(n_569));
	notech_and2 i_181(.A(n_440), .B(divq[53]), .Z(n_862));
	notech_nand2 i_180(.A(n_439), .B(divq[52]), .Z(n_567));
	notech_and2 i_179(.A(n_438), .B(divq[51]), .Z(n_861));
	notech_nand2 i_178(.A(n_437), .B(divq[50]), .Z(n_565));
	notech_and2 i_177(.A(n_436), .B(divq[49]), .Z(n_860));
	notech_nand2 i_176(.A(n_435), .B(divq[48]), .Z(n_563));
	notech_and2 i_175(.A(n_434), .B(divq[47]), .Z(n_859));
	notech_nand2 i_174(.A(n_433), .B(divq[46]), .Z(n_561));
	notech_and2 i_173(.A(n_432), .B(divq[45]), .Z(n_858));
	notech_nand2 i_172(.A(n_431), .B(divq[44]), .Z(n_559));
	notech_and2 i_171(.A(n_430), .B(divq[43]), .Z(n_857));
	notech_nand2 i_170(.A(n_429), .B(divq[42]), .Z(n_557));
	notech_and2 i_169(.A(n_428), .B(divq[41]), .Z(n_856));
	notech_nand2 i_168(.A(n_427), .B(divq[40]), .Z(n_555));
	notech_and2 i_167(.A(n_426), .B(divq[39]), .Z(n_855));
	notech_nand2 i_166(.A(n_425), .B(divq[38]), .Z(n_553));
	notech_and2 i_165(.A(n_424), .B(divq[37]), .Z(n_854));
	notech_nand2 i_164(.A(n_423), .B(divq[36]), .Z(n_551));
	notech_and2 i_163(.A(n_422), .B(divq[35]), .Z(n_853));
	notech_nand2 i_162(.A(n_421), .B(divq[34]), .Z(n_549));
	notech_and2 i_161(.A(n_420), .B(divq[33]), .Z(n_852));
	notech_nand2 i_160(.A(n_419), .B(divq[32]), .Z(n_547));
	notech_and2 i_159(.A(n_418), .B(divq[31]), .Z(n_851));
	notech_nand2 i_158(.A(n_417), .B(divq[30]), .Z(n_545));
	notech_and2 i_157(.A(n_416), .B(divq[29]), .Z(n_850));
	notech_nand2 i_156(.A(n_415), .B(divq[28]), .Z(n_543));
	notech_and2 i_155(.A(n_414), .B(divq[27]), .Z(n_849));
	notech_nand2 i_154(.A(n_413), .B(divq[26]), .Z(n_541));
	notech_and2 i_153(.A(n_412), .B(divq[25]), .Z(n_848));
	notech_nand2 i_152(.A(n_411), .B(divq[24]), .Z(n_539));
	notech_and2 i_151(.A(n_410), .B(divq[23]), .Z(n_847));
	notech_nand2 i_150(.A(n_409), .B(divq[22]), .Z(n_537));
	notech_and2 i_149(.A(n_408), .B(divq[21]), .Z(n_846));
	notech_nand2 i_148(.A(n_407), .B(divq[20]), .Z(n_535));
	notech_and2 i_147(.A(n_406), .B(divq[19]), .Z(n_845));
	notech_nand2 i_146(.A(n_405), .B(divq[18]), .Z(n_533));
	notech_and2 i_145(.A(n_404), .B(divq[17]), .Z(n_844));
	notech_nand2 i_144(.A(n_403), .B(divq[16]), .Z(n_531));
	notech_and2 i_143(.A(n_402), .B(divq[15]), .Z(n_843));
	notech_nand2 i_142(.A(n_401), .B(divq[14]), .Z(n_529));
	notech_and2 i_141(.A(n_400), .B(divq[13]), .Z(n_842));
	notech_nand2 i_140(.A(n_399), .B(divq[12]), .Z(n_527));
	notech_and2 i_139(.A(n_398), .B(divq[11]), .Z(n_841));
	notech_nand2 i_138(.A(n_397), .B(divq[10]), .Z(n_525));
	notech_and2 i_137(.A(n_396), .B(divq[9]), .Z(n_840));
	notech_nand2 i_136(.A(n_395), .B(divq[8]), .Z(n_523));
	notech_and2 i_135(.A(n_394), .B(divq[7]), .Z(n_839));
	notech_nand2 i_134(.A(n_393), .B(divq[6]), .Z(n_521));
	notech_and2 i_133(.A(n_392), .B(divq[5]), .Z(n_838));
	notech_nand2 i_132(.A(n_391), .B(divq[4]), .Z(n_519));
	notech_and2 i_131(.A(n_390), .B(divq[3]), .Z(n_837));
	notech_nand2 i_130(.A(n_389), .B(divq[2]), .Z(n_517));
	notech_and2 i_129(.A(n_388), .B(divq[1]), .Z(n_836));
	notech_nand2 i_128(.A(n_387), .B(divq[0]), .Z(n_515));
	notech_nor2 i_125(.A(n_449), .B(divq[62]), .Z(n_512));
	notech_nor2 i_124(.A(n_448), .B(divq[61]), .Z(n_511));
	notech_nor2 i_123(.A(n_447), .B(divq[60]), .Z(n_510));
	notech_nor2 i_122(.A(n_446), .B(divq[59]), .Z(n_509));
	notech_nor2 i_121(.A(n_445), .B(divq[58]), .Z(n_508));
	notech_nor2 i_120(.A(n_444), .B(divq[57]), .Z(n_507));
	notech_nor2 i_119(.A(n_443), .B(divq[56]), .Z(n_506));
	notech_nor2 i_118(.A(n_442), .B(divq[55]), .Z(n_505));
	notech_nor2 i_117(.A(n_441), .B(divq[54]), .Z(n_504));
	notech_nor2 i_116(.A(n_440), .B(divq[53]), .Z(n_503));
	notech_nor2 i_115(.A(n_439), .B(divq[52]), .Z(n_502));
	notech_nor2 i_114(.A(n_438), .B(divq[51]), .Z(n_501));
	notech_nor2 i_113(.A(n_437), .B(divq[50]), .Z(n_500));
	notech_nor2 i_112(.A(n_436), .B(divq[49]), .Z(n_499));
	notech_nor2 i_111(.A(n_435), .B(divq[48]), .Z(n_498));
	notech_nor2 i_110(.A(n_434), .B(divq[47]), .Z(n_497));
	notech_nor2 i_109(.A(n_433), .B(divq[46]), .Z(n_496));
	notech_nor2 i_108(.A(n_432), .B(divq[45]), .Z(n_495));
	notech_nor2 i_107(.A(n_431), .B(divq[44]), .Z(n_494));
	notech_nor2 i_106(.A(n_430), .B(divq[43]), .Z(n_493));
	notech_nor2 i_105(.A(n_429), .B(divq[42]), .Z(n_492));
	notech_nor2 i_104(.A(n_428), .B(divq[41]), .Z(n_491));
	notech_nor2 i_103(.A(n_427), .B(divq[40]), .Z(n_490));
	notech_nor2 i_102(.A(n_426), .B(divq[39]), .Z(n_489));
	notech_nor2 i_101(.A(n_425), .B(divq[38]), .Z(n_488));
	notech_nor2 i_100(.A(n_424), .B(divq[37]), .Z(n_487));
	notech_nor2 i_99(.A(n_423), .B(divq[36]), .Z(n_486));
	notech_nor2 i_98(.A(n_422), .B(divq[35]), .Z(n_485));
	notech_nor2 i_97(.A(n_421), .B(divq[34]), .Z(n_484));
	notech_nor2 i_96(.A(n_420), .B(divq[33]), .Z(n_483));
	notech_nor2 i_95(.A(n_419), .B(divq[32]), .Z(n_482));
	notech_nor2 i_94(.A(n_418), .B(divq[31]), .Z(n_481));
	notech_nor2 i_93(.A(n_417), .B(divq[30]), .Z(n_480));
	notech_nor2 i_92(.A(n_416), .B(divq[29]), .Z(n_479));
	notech_nor2 i_91(.A(n_415), .B(divq[28]), .Z(n_478));
	notech_nor2 i_90(.A(n_414), .B(divq[27]), .Z(n_477));
	notech_nor2 i_89(.A(n_413), .B(divq[26]), .Z(n_476));
	notech_nor2 i_88(.A(n_412), .B(divq[25]), .Z(n_475));
	notech_nor2 i_87(.A(n_411), .B(divq[24]), .Z(n_474));
	notech_nor2 i_86(.A(n_410), .B(divq[23]), .Z(n_473));
	notech_nor2 i_85(.A(n_409), .B(divq[22]), .Z(n_472));
	notech_nor2 i_84(.A(n_408), .B(divq[21]), .Z(n_471));
	notech_nor2 i_83(.A(n_407), .B(divq[20]), .Z(n_470));
	notech_nor2 i_82(.A(n_406), .B(divq[19]), .Z(n_469));
	notech_nor2 i_81(.A(n_405), .B(divq[18]), .Z(n_468));
	notech_nor2 i_80(.A(n_404), .B(divq[17]), .Z(n_467));
	notech_nor2 i_79(.A(n_403), .B(divq[16]), .Z(n_466));
	notech_nor2 i_78(.A(n_402), .B(divq[15]), .Z(n_465));
	notech_nor2 i_77(.A(n_401), .B(divq[14]), .Z(n_464));
	notech_nor2 i_76(.A(n_400), .B(divq[13]), .Z(n_463));
	notech_nor2 i_75(.A(n_399), .B(divq[12]), .Z(n_462));
	notech_nor2 i_74(.A(n_398), .B(divq[11]), .Z(n_461));
	notech_nor2 i_73(.A(n_397), .B(divq[10]), .Z(n_460));
	notech_nor2 i_72(.A(n_396), .B(divq[9]), .Z(n_459));
	notech_nor2 i_71(.A(n_395), .B(divq[8]), .Z(n_458));
	notech_nor2 i_70(.A(n_394), .B(divq[7]), .Z(n_457));
	notech_nor2 i_69(.A(n_393), .B(divq[6]), .Z(n_456));
	notech_nor2 i_68(.A(n_392), .B(divq[5]), .Z(n_455));
	notech_nor2 i_67(.A(n_391), .B(divq[4]), .Z(n_454));
	notech_nor2 i_66(.A(n_390), .B(divq[3]), .Z(n_453));
	notech_nor2 i_65(.A(n_389), .B(divq[2]), .Z(n_452));
	notech_nor2 i_64(.A(n_388), .B(divq[1]), .Z(n_451));
	notech_inv i_62(.A(I0[62]), .Z(n_449));
	notech_inv i_61(.A(I0[61]), .Z(n_448));
	notech_inv i_60(.A(I0[60]), .Z(n_447));
	notech_inv i_59(.A(I0[59]), .Z(n_446));
	notech_inv i_58(.A(I0[58]), .Z(n_445));
	notech_inv i_57(.A(I0[57]), .Z(n_444));
	notech_inv i_56(.A(I0[56]), .Z(n_443));
	notech_inv i_55(.A(I0[55]), .Z(n_442));
	notech_inv i_54(.A(I0[54]), .Z(n_441));
	notech_inv i_53(.A(I0[53]), .Z(n_440));
	notech_inv i_52(.A(I0[52]), .Z(n_439));
	notech_inv i_51(.A(I0[51]), .Z(n_438));
	notech_inv i_50(.A(I0[50]), .Z(n_437));
	notech_inv i_49(.A(I0[49]), .Z(n_436));
	notech_inv i_48(.A(I0[48]), .Z(n_435));
	notech_inv i_47(.A(I0[47]), .Z(n_434));
	notech_inv i_46(.A(I0[46]), .Z(n_433));
	notech_inv i_45(.A(I0[45]), .Z(n_432));
	notech_inv i_44(.A(I0[44]), .Z(n_431));
	notech_inv i_43(.A(I0[43]), .Z(n_430));
	notech_inv i_42(.A(I0[42]), .Z(n_429));
	notech_inv i_41(.A(I0[41]), .Z(n_428));
	notech_inv i_40(.A(I0[40]), .Z(n_427));
	notech_inv i_39(.A(I0[39]), .Z(n_426));
	notech_inv i_38(.A(I0[38]), .Z(n_425));
	notech_inv i_37(.A(I0[37]), .Z(n_424));
	notech_inv i_36(.A(I0[36]), .Z(n_423));
	notech_inv i_35(.A(I0[35]), .Z(n_422));
	notech_inv i_34(.A(I0[34]), .Z(n_421));
	notech_inv i_33(.A(I0[33]), .Z(n_420));
	notech_inv i_32(.A(I0[32]), .Z(n_419));
	notech_inv i_31(.A(I0[31]), .Z(n_418));
	notech_inv i_30(.A(I0[30]), .Z(n_417));
	notech_inv i_29(.A(I0[29]), .Z(n_416));
	notech_inv i_28(.A(I0[28]), .Z(n_415));
	notech_inv i_27(.A(I0[27]), .Z(n_414));
	notech_inv i_26(.A(I0[26]), .Z(n_413));
	notech_inv i_25(.A(I0[25]), .Z(n_412));
	notech_inv i_24(.A(I0[24]), .Z(n_411));
	notech_inv i_23(.A(I0[23]), .Z(n_410));
	notech_inv i_22(.A(I0[22]), .Z(n_409));
	notech_inv i_21(.A(I0[21]), .Z(n_408));
	notech_inv i_20(.A(I0[20]), .Z(n_407));
	notech_inv i_19(.A(I0[19]), .Z(n_406));
	notech_inv i_18(.A(I0[18]), .Z(n_405));
	notech_inv i_17(.A(I0[17]), .Z(n_404));
	notech_inv i_16(.A(I0[16]), .Z(n_403));
	notech_inv i_15(.A(I0[15]), .Z(n_402));
	notech_inv i_14(.A(I0[14]), .Z(n_401));
	notech_inv i_13(.A(I0[13]), .Z(n_400));
	notech_inv i_12(.A(I0[12]), .Z(n_399));
	notech_inv i_11(.A(I0[11]), .Z(n_398));
	notech_inv i_10(.A(I0[10]), .Z(n_397));
	notech_inv i_9(.A(I0[9]), .Z(n_396));
	notech_inv i_8(.A(I0[8]), .Z(n_395));
	notech_inv i_7(.A(I0[7]), .Z(n_394));
	notech_inv i_6(.A(I0[6]), .Z(n_393));
	notech_inv i_5(.A(I0[5]), .Z(n_392));
	notech_inv i_4(.A(I0[4]), .Z(n_391));
	notech_inv i_3(.A(I0[3]), .Z(n_390));
	notech_inv i_2(.A(I0[2]), .Z(n_389));
	notech_inv i_1(.A(I0[1]), .Z(n_388));
	notech_inv i_0(.A(I0[0]), .Z(n_387));
endmodule
module AWDP_LSH_10(O0, opd);
    output [31:0] O0;
    input [5:0] opd;
    // Line 1006
    wire [31:0] N745;
    wire [31:0] O0;

    // Line 1006
    assign N745 = 6'h1 << opd;
    assign O0 = N745;
endmodule

module AWDP_LSH_40(O0, opb);
    output [31:0] O0;
    input [4:0] opb;
    // Line 636
    wire [31:0] N755;
    // Line 348
    wire [31:0] O0;

    // Line 636
    assign N755 = 5'h1 << opb;
    // Line 348
    assign O0 = N755;
endmodule

module AWDP_SUB_129(O0, regs_7, opd);
    output [31:0] O0;
    input [31:0] regs_7;
    input [31:0] opd;
    // Line 521
    wire [31:0] N771;
    // Line 348
    wire [31:0] O0;

    // Line 521
    assign N771 = regs_7 - opd;
    // Line 348
    assign O0 = N771;
endmodule

module AWDP_SUB_139(O0, regs_6, opd);
    output [31:0] O0;
    input [31:0] regs_6;
    input [31:0] opd;
    // Line 348
    wire [31:0] O0;
    // Line 521
    wire [31:0] N785;

    // Line 348
    assign O0 = N785;
    // Line 521
    assign N785 = regs_6 - opd;
endmodule

module AWDP_SUB_176(O0, opa, I0);

	output [32:0] O0;
	input [31:0] opa;
	input [31:0] I0;




	notech_inv i_10184(.A(n_58104), .Z(n_58105));
	notech_inv i_10183(.A(I0[19]), .Z(n_58104));
	notech_inv i_64(.A(n_454), .Z(O0[32]));
	notech_fa2 i_63(.A(n_58104), .B(n_452), .CI(opa[31]), .Z(O0[31]), .CO(n_454
		));
	notech_fa2 i_62(.A(n_58104), .B(n_450), .CI(opa[30]), .Z(O0[30]), .CO(n_452
		));
	notech_fa2 i_61(.A(n_58104), .B(n_448), .CI(opa[29]), .Z(O0[29]), .CO(n_450
		));
	notech_fa2 i_60(.A(n_58104), .B(n_446), .CI(opa[28]), .Z(O0[28]), .CO(n_448
		));
	notech_fa2 i_59(.A(n_58104), .B(n_444), .CI(opa[27]), .Z(O0[27]), .CO(n_446
		));
	notech_fa2 i_58(.A(n_58104), .B(n_442), .CI(opa[26]), .Z(O0[26]), .CO(n_444
		));
	notech_fa2 i_57(.A(n_58104), .B(n_440), .CI(opa[25]), .Z(O0[25]), .CO(n_442
		));
	notech_fa2 i_56(.A(n_58104), .B(n_438), .CI(opa[24]), .Z(O0[24]), .CO(n_440
		));
	notech_fa2 i_55(.A(n_58104), .B(n_436), .CI(opa[23]), .Z(O0[23]), .CO(n_438
		));
	notech_fa2 i_54(.A(n_58104), .B(n_434), .CI(opa[22]), .Z(O0[22]), .CO(n_436
		));
	notech_fa2 i_53(.A(n_58104), .B(n_432), .CI(opa[21]), .Z(O0[21]), .CO(n_434
		));
	notech_fa2 i_52(.A(n_58104), .B(n_430), .CI(opa[20]), .Z(O0[20]), .CO(n_432
		));
	notech_fa2 i_51(.A(n_58104), .B(n_428), .CI(opa[19]), .Z(O0[19]), .CO(n_430
		));
	notech_fa2 i_50(.A(n_58104), .B(n_426), .CI(opa[18]), .Z(O0[18]), .CO(n_428
		));
	notech_fa2 i_49(.A(n_58104), .B(n_424), .CI(opa[17]), .Z(O0[17]), .CO(n_426
		));
	notech_fa2 i_48(.A(n_361), .B(n_422), .CI(opa[16]), .Z(O0[16]), .CO(n_424
		));
	notech_fa2 i_47(.A(n_361), .B(n_420), .CI(opa[15]), .Z(O0[15]), .CO(n_422
		));
	notech_fa2 i_46(.A(n_361), .B(n_418), .CI(opa[14]), .Z(O0[14]), .CO(n_420
		));
	notech_fa2 i_45(.A(n_361), .B(n_416), .CI(opa[13]), .Z(O0[13]), .CO(n_418
		));
	notech_fa2 i_44(.A(n_361), .B(n_414), .CI(opa[12]), .Z(O0[12]), .CO(n_416
		));
	notech_fa2 i_43(.A(n_361), .B(n_412), .CI(opa[11]), .Z(O0[11]), .CO(n_414
		));
	notech_fa2 i_42(.A(n_361), .B(n_410), .CI(opa[10]), .Z(O0[10]), .CO(n_412
		));
	notech_fa2 i_41(.A(n_361), .B(n_408), .CI(opa[9]), .Z(O0[9]), .CO(n_410)
		);
	notech_fa2 i_40(.A(n_361), .B(n_406), .CI(opa[8]), .Z(O0[8]), .CO(n_408)
		);
	notech_fa2 i_39(.A(n_361), .B(n_404), .CI(opa[7]), .Z(O0[7]), .CO(n_406)
		);
	notech_fa2 i_38(.A(n_361), .B(n_402), .CI(opa[6]), .Z(O0[6]), .CO(n_404)
		);
	notech_fa2 i_37(.A(n_361), .B(n_400), .CI(opa[5]), .Z(O0[5]), .CO(n_402)
		);
	notech_fa2 i_36(.A(n_361), .B(n_398), .CI(opa[4]), .Z(O0[4]), .CO(n_400)
		);
	notech_fa2 i_35(.A(n_361), .B(n_396), .CI(opa[3]), .Z(O0[3]), .CO(n_398)
		);
	notech_fa2 i_34(.A(n_361), .B(n_394), .CI(opa[2]), .Z(O0[2]), .CO(n_396)
		);
	notech_fa2 i_33(.A(n_360), .B(n_392), .CI(opa[1]), .Z(O0[1]), .CO(n_394)
		);
	notech_inv i_2(.A(n_58105), .Z(n_361));
	notech_inv i_1(.A(I0[1]), .Z(n_360));
	notech_inv i_0(.A(I0[0]), .Z(n_359));
	notech_xor2 i_81(.A(opa[0]), .B(n_359), .Z(n_47003));
	notech_inv i_82(.A(n_47003), .Z(O0[0]));
	notech_or2 i_80(.A(opa[0]), .B(n_359), .Z(n_392));
endmodule
module AWDP_SUB_192(O0, opd);

	output [31:0] O0;
	input [31:0] opd;

	wire \opd[2] ;
	wire \opd[3] ;
	wire \opd[4] ;
	wire \opd[5] ;
	wire \opd[6] ;
	wire \opd[7] ;
	wire \opd[8] ;
	wire \opd[9] ;
	wire \opd[10] ;
	wire \opd[11] ;
	wire \opd[12] ;
	wire \opd[13] ;
	wire \opd[14] ;
	wire \opd[15] ;
	wire \opd[16] ;
	wire \opd[17] ;
	wire \opd[18] ;
	wire \opd[19] ;
	wire \opd[20] ;
	wire \opd[21] ;
	wire \opd[22] ;
	wire \opd[23] ;
	wire \opd[24] ;
	wire \opd[25] ;
	wire \opd[26] ;
	wire \opd[27] ;
	wire \opd[28] ;
	wire \opd[29] ;
	wire \opd[30] ;
	wire \opd[31] ;


	assign O0[0] = opd[0];
	assign O0[1] = opd[1];
	assign \opd[2]  = opd[2];
	assign \opd[3]  = opd[3];
	assign \opd[4]  = opd[4];
	assign \opd[5]  = opd[5];
	assign \opd[6]  = opd[6];
	assign \opd[7]  = opd[7];
	assign \opd[8]  = opd[8];
	assign \opd[9]  = opd[9];
	assign \opd[10]  = opd[10];
	assign \opd[11]  = opd[11];
	assign \opd[12]  = opd[12];
	assign \opd[13]  = opd[13];
	assign \opd[14]  = opd[14];
	assign \opd[15]  = opd[15];
	assign \opd[16]  = opd[16];
	assign \opd[17]  = opd[17];
	assign \opd[18]  = opd[18];
	assign \opd[19]  = opd[19];
	assign \opd[20]  = opd[20];
	assign \opd[21]  = opd[21];
	assign \opd[22]  = opd[22];
	assign \opd[23]  = opd[23];
	assign \opd[24]  = opd[24];
	assign \opd[25]  = opd[25];
	assign \opd[26]  = opd[26];
	assign \opd[27]  = opd[27];
	assign \opd[28]  = opd[28];
	assign \opd[29]  = opd[29];
	assign \opd[30]  = opd[30];
	assign \opd[31]  = opd[31];

	notech_ha2 i_30(.A(n_192), .B(n_250), .Z(O0[31]));
	notech_inv i_1(.A(\opd[2] ), .Z(O0[2]));
	notech_inv i_0(.A(\opd[31] ), .Z(n_192));
	notech_xor2 i_47(.A(\opd[30] ), .B(n_248), .Z(n_47030));
	notech_inv i_48(.A(n_47030), .Z(O0[30]));
	notech_or2 i_46(.A(\opd[30] ), .B(n_248), .Z(n_250));
	notech_xor2 i_4698939(.A(\opd[29] ), .B(n_246), .Z(n_47057));
	notech_inv i_4798940(.A(n_47057), .Z(O0[29]));
	notech_or2 i_45(.A(\opd[29] ), .B(n_246), .Z(n_248));
	notech_xor2 i_44(.A(\opd[28] ), .B(n_244), .Z(n_47084));
	notech_inv i_4598941(.A(n_47084), .Z(O0[28]));
	notech_or2 i_43(.A(\opd[28] ), .B(n_244), .Z(n_246));
	notech_xor2 i_4398942(.A(\opd[27] ), .B(n_242), .Z(n_47111));
	notech_inv i_4498943(.A(n_47111), .Z(O0[27]));
	notech_or2 i_42(.A(\opd[27] ), .B(n_242), .Z(n_244));
	notech_xor2 i_4298944(.A(\opd[26] ), .B(n_240), .Z(n_47138));
	notech_inv i_4398945(.A(n_47138), .Z(O0[26]));
	notech_or2 i_41(.A(\opd[26] ), .B(n_240), .Z(n_242));
	notech_xor2 i_4198946(.A(\opd[25] ), .B(n_238), .Z(n_47165));
	notech_inv i_4298947(.A(n_47165), .Z(O0[25]));
	notech_or2 i_40(.A(\opd[25] ), .B(n_238), .Z(n_240));
	notech_xor2 i_4098948(.A(\opd[24] ), .B(n_236), .Z(n_47192));
	notech_inv i_4198949(.A(n_47192), .Z(O0[24]));
	notech_or2 i_39(.A(\opd[24] ), .B(n_236), .Z(n_238));
	notech_xor2 i_3998950(.A(\opd[23] ), .B(n_234), .Z(n_47219));
	notech_inv i_4098951(.A(n_47219), .Z(O0[23]));
	notech_or2 i_38(.A(\opd[23] ), .B(n_234), .Z(n_236));
	notech_xor2 i_3898952(.A(\opd[22] ), .B(n_232), .Z(n_47246));
	notech_inv i_3998953(.A(n_47246), .Z(O0[22]));
	notech_or2 i_37(.A(\opd[22] ), .B(n_232), .Z(n_234));
	notech_xor2 i_3798954(.A(\opd[21] ), .B(n_230), .Z(n_47273));
	notech_inv i_3898955(.A(n_47273), .Z(O0[21]));
	notech_or2 i_36(.A(\opd[21] ), .B(n_230), .Z(n_232));
	notech_xor2 i_3698956(.A(\opd[20] ), .B(n_228), .Z(n_47300));
	notech_inv i_3798957(.A(n_47300), .Z(O0[20]));
	notech_or2 i_35(.A(\opd[20] ), .B(n_228), .Z(n_230));
	notech_xor2 i_3598958(.A(\opd[19] ), .B(n_226), .Z(n_47327));
	notech_inv i_3698959(.A(n_47327), .Z(O0[19]));
	notech_or2 i_34(.A(\opd[19] ), .B(n_226), .Z(n_228));
	notech_xor2 i_3498960(.A(\opd[18] ), .B(n_224), .Z(n_47354));
	notech_inv i_3598961(.A(n_47354), .Z(O0[18]));
	notech_or2 i_33(.A(\opd[18] ), .B(n_224), .Z(n_226));
	notech_xor2 i_3398962(.A(\opd[17] ), .B(n_222), .Z(n_47381));
	notech_inv i_3498963(.A(n_47381), .Z(O0[17]));
	notech_or2 i_32(.A(\opd[17] ), .B(n_222), .Z(n_224));
	notech_xor2 i_3298964(.A(\opd[16] ), .B(n_220), .Z(n_47408));
	notech_inv i_3398965(.A(n_47408), .Z(O0[16]));
	notech_or2 i_31(.A(\opd[16] ), .B(n_220), .Z(n_222));
	notech_xor2 i_3198966(.A(\opd[15] ), .B(n_218), .Z(n_47435));
	notech_inv i_3298967(.A(n_47435), .Z(O0[15]));
	notech_or2 i_3098968(.A(\opd[15] ), .B(n_218), .Z(n_220));
	notech_xor2 i_3098969(.A(\opd[14] ), .B(n_216), .Z(n_47462));
	notech_inv i_3198970(.A(n_47462), .Z(O0[14]));
	notech_or2 i_29(.A(\opd[14] ), .B(n_216), .Z(n_218));
	notech_xor2 i_2998971(.A(\opd[13] ), .B(n_214), .Z(n_47489));
	notech_inv i_3098972(.A(n_47489), .Z(O0[13]));
	notech_or2 i_28(.A(\opd[13] ), .B(n_214), .Z(n_216));
	notech_xor2 i_2898973(.A(\opd[12] ), .B(n_212), .Z(n_47516));
	notech_inv i_2998974(.A(n_47516), .Z(O0[12]));
	notech_or2 i_27(.A(\opd[12] ), .B(n_212), .Z(n_214));
	notech_xor2 i_2798975(.A(\opd[11] ), .B(n_210), .Z(n_47543));
	notech_inv i_2898976(.A(n_47543), .Z(O0[11]));
	notech_or2 i_26(.A(\opd[11] ), .B(n_210), .Z(n_212));
	notech_xor2 i_2798977(.A(\opd[10] ), .B(n_208), .Z(n_47570));
	notech_inv i_2898978(.A(n_47570), .Z(O0[10]));
	notech_or2 i_2698979(.A(\opd[10] ), .B(n_208), .Z(n_210));
	notech_xor2 i_2798980(.A(\opd[9] ), .B(n_206), .Z(n_47597));
	notech_inv i_2898981(.A(n_47597), .Z(O0[9]));
	notech_or2 i_2698982(.A(\opd[9] ), .B(n_206), .Z(n_208));
	notech_xor2 i_2798983(.A(\opd[8] ), .B(n_204), .Z(n_47624));
	notech_inv i_2898984(.A(n_47624), .Z(O0[8]));
	notech_or2 i_2698985(.A(\opd[8] ), .B(n_204), .Z(n_206));
	notech_xor2 i_2798986(.A(\opd[7] ), .B(n_202), .Z(n_47651));
	notech_inv i_2898987(.A(n_47651), .Z(O0[7]));
	notech_or2 i_2698988(.A(\opd[7] ), .B(n_202), .Z(n_204));
	notech_xor2 i_2798989(.A(\opd[6] ), .B(n_200), .Z(n_47678));
	notech_inv i_2898990(.A(n_47678), .Z(O0[6]));
	notech_or2 i_2698991(.A(\opd[6] ), .B(n_200), .Z(n_202));
	notech_xor2 i_2798992(.A(\opd[5] ), .B(n_198), .Z(n_47705));
	notech_inv i_2898993(.A(n_47705), .Z(O0[5]));
	notech_or2 i_2698994(.A(\opd[5] ), .B(n_198), .Z(n_200));
	notech_xor2 i_2798995(.A(\opd[4] ), .B(n_196), .Z(n_47732));
	notech_inv i_2898996(.A(n_47732), .Z(O0[4]));
	notech_or2 i_2698997(.A(\opd[4] ), .B(n_196), .Z(n_198));
	notech_xor2 i_2798998(.A(\opd[3] ), .B(\opd[2] ), .Z(n_47760));
	notech_inv i_2898999(.A(n_47760), .Z(O0[3]));
	notech_or2 i_2699000(.A(\opd[3] ), .B(\opd[2] ), .Z(n_196));
endmodule
module AWDP_SUB_237(O0, opa, I0);

	output [16:0] O0;
	input [15:0] opa;
	input [15:0] I0;




	notech_inv i_10191(.A(I0[13]), .Z(n_58142));
	notech_inv i_32(.A(n_230), .Z(O0[16]));
	notech_fa2 i_31(.A(n_58142), .B(n_228), .CI(opa[15]), .Z(O0[15]), .CO(n_230
		));
	notech_fa2 i_30(.A(n_58142), .B(n_226), .CI(opa[14]), .Z(O0[14]), .CO(n_228
		));
	notech_fa2 i_29(.A(n_58142), .B(n_224), .CI(opa[13]), .Z(O0[13]), .CO(n_226
		));
	notech_fa2 i_28(.A(n_58142), .B(n_222), .CI(opa[12]), .Z(O0[12]), .CO(n_224
		));
	notech_fa2 i_27(.A(n_58142), .B(n_220), .CI(opa[11]), .Z(O0[11]), .CO(n_222
		));
	notech_fa2 i_26(.A(n_58142), .B(n_218), .CI(opa[10]), .Z(O0[10]), .CO(n_220
		));
	notech_fa2 i_25(.A(n_58142), .B(n_216), .CI(opa[9]), .Z(O0[9]), .CO(n_218
		));
	notech_fa2 i_24(.A(n_58142), .B(n_214), .CI(opa[8]), .Z(O0[8]), .CO(n_216
		));
	notech_fa2 i_23(.A(n_58142), .B(n_212), .CI(opa[7]), .Z(O0[7]), .CO(n_214
		));
	notech_fa2 i_22(.A(n_58142), .B(n_210), .CI(opa[6]), .Z(O0[6]), .CO(n_212
		));
	notech_fa2 i_21(.A(n_58142), .B(n_208), .CI(opa[5]), .Z(O0[5]), .CO(n_210
		));
	notech_fa2 i_20(.A(n_58142), .B(n_206), .CI(opa[4]), .Z(O0[4]), .CO(n_208
		));
	notech_fa2 i_19(.A(n_58142), .B(n_204), .CI(opa[3]), .Z(O0[3]), .CO(n_206
		));
	notech_fa2 i_18(.A(n_58142), .B(n_202), .CI(opa[2]), .Z(O0[2]), .CO(n_204
		));
	notech_fa2 i_17(.A(n_184), .B(n_200), .CI(opa[1]), .Z(O0[1]), .CO(n_202)
		);
	notech_inv i_1(.A(I0[1]), .Z(n_184));
	notech_inv i_0(.A(I0[0]), .Z(n_183));
	notech_xor2 i_49(.A(opa[0]), .B(n_183), .Z(n_47787));
	notech_inv i_50(.A(n_47787), .Z(O0[0]));
	notech_or2 i_48(.A(opa[0]), .B(n_183), .Z(n_200));
endmodule
module AWDP_SUB_37(O0, regs_4, calc_sz);
    output [31:0] O0;
    input [31:0] regs_4;
    input [2:0] calc_sz;
    // Line 348
    wire [31:0] O0;
    // Line 456
    wire [31:0] N831;

    // Line 348
    assign O0 = N831;
    // Line 456
    assign N831 = regs_4 - calc_sz;
endmodule

module AWDP_SUB_39(O0, divr, divq);
    output [63:0] O0;
    input [63:0] divr;
    input [63:0] divq;
    // Line 1006
    wire [63:0] O0;
    // Line 1006
    wire [63:0] N843;

    // Line 1006
    assign O0 = N843;
    // Line 1006
    assign N843 = divr - divq;
endmodule

module AWMUX_16_1(I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14
		, I15, S, O0);

	input I0;
	input I1;
	input I2;
	input I3;
	input I4;
	input I5;
	input I6;
	input I7;
	input I8;
	input I9;
	input I10;
	input I11;
	input I12;
	input I13;
	input I14;
	input I15;
	input [3:0] S;
	output O0;




	notech_inv i_15554(.A(n_63721), .Z(n_63722));
	notech_inv i_15553(.A(S[1]), .Z(n_63721));
	notech_mux4 i_14(.S0(S[2]), .S1(S[3]), .A(n_23), .B(n_26), .C(n_29), .D(n_32
		), .Z(O0));
	notech_mux4 i_11(.S0(S[0]), .S1(n_63722), .A(I12), .B(n_18767), .C(I14),
		 .D(n_18766), .Z(n_32));
	notech_mux4 i_8(.S0(S[0]), .S1(n_63722), .A(I8), .B(n_18769), .C(I10), .D
		(n_18768), .Z(n_29));
	notech_mux4 i_5(.S0(S[0]), .S1(n_63722), .A(I4), .B(n_18771), .C(I6), .D
		(n_18770), .Z(n_26));
	notech_mux4 i_2(.S0(S[0]), .S1(n_63722), .A(I0), .B(n_18773), .C(I2), .D
		(n_18772), .Z(n_23));
	notech_inv i_19(.A(I14), .Z(n_18766));
	notech_inv i_20(.A(I12), .Z(n_18767));
	notech_inv i_21(.A(I10), .Z(n_18768));
	notech_inv i_22(.A(I8), .Z(n_18769));
	notech_inv i_23(.A(I6), .Z(n_18770));
	notech_inv i_24(.A(I4), .Z(n_18771));
	notech_inv i_25(.A(I2), .Z(n_18772));
	notech_inv i_26(.A(I0), .Z(n_18773));
endmodule
module AWMUX_16_32_0(I0 , I1 , I2 , I3 , I4 , I5 , I6 , I7 , I8 , I9 , I10 , I11 , I12 , I13 , I14 , I15 , S , O0);
input  [31:0] I0;
input  [31:0] I1;
input  [31:0] I2;
input  [31:0] I3;
input  [31:0] I4;
input  [31:0] I5;
input  [31:0] I6;
input  [31:0] I7;
input  [31:0] I8;
input  [31:0] I9;
input  [31:0] I10;
input  [31:0] I11;
input  [31:0] I12;
input  [31:0] I13;
input  [31:0] I14;
input  [31:0] I15;
input  [3:0] S;
output  [31:0] O0;
reg [31:0] O0;

always @(I0 or I1 or I2 or I3 or I4 or I5 or I6 or I7 or I8 or I9 or I10 or I11 or I12 or I13 or I14 or I15 or S or O0)
begin
	case(S)
	4'h0 : O0 = I0;
	4'h1 : O0 = I1;
	4'h2 : O0 = I2;
	4'h3 : O0 = I3;
	4'h4 : O0 = I4;
	4'h5 : O0 = I5;
	4'h6 : O0 = I6;
	4'h7 : O0 = I7;
	4'h8 : O0 = I8;
	4'h9 : O0 = I9;
	4'ha : O0 = I10;
	4'hb : O0 = I11;
	4'hc : O0 = I12;
	4'hd : O0 = I13;
	4'he : O0 = I14;
	default : O0 = I15;
	endcase
end
endmodule

module AWMUX_16_32_1(I0 , I1 , I2 , I3 , I4 , I5 , I6 , I7 , I8 , I9 , I10 , I11 , I12 , I13 , I14 , I15 , S , O0);
input  [31:0] I0;
input  [31:0] I1;
input  [31:0] I2;
input  [31:0] I3;
input  [31:0] I4;
input  [31:0] I5;
input  [31:0] I6;
input  [31:0] I7;
input  [31:0] I8;
input  [31:0] I9;
input  [31:0] I10;
input  [31:0] I11;
input  [31:0] I12;
input  [31:0] I13;
input  [31:0] I14;
input  [31:0] I15;
input  [3:0] S;
output  [31:0] O0;
reg [31:0] O0;

always @(I0 or I1 or I2 or I3 or I4 or I5 or I6 or I7 or I8 or I9 or I10 or I11 or I12 or I13 or I14 or I15 or S or O0)
begin
	case(S)
	4'h0 : O0 = I0;
	4'h1 : O0 = I1;
	4'h2 : O0 = I2;
	4'h3 : O0 = I3;
	4'h4 : O0 = I4;
	4'h5 : O0 = I5;
	4'h6 : O0 = I6;
	4'h7 : O0 = I7;
	4'h8 : O0 = I8;
	4'h9 : O0 = I9;
	4'ha : O0 = I10;
	4'hb : O0 = I11;
	4'hc : O0 = I12;
	4'hd : O0 = I13;
	4'he : O0 = I14;
	default : O0 = I15;
	endcase
end
endmodule

module AWMUX_16_32_2(I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13,
		 I14, I15, S, O0);

	input [31:0] I0;
	input [31:0] I1;
	input [31:0] I2;
	input [31:0] I3;
	input [31:0] I4;
	input [31:0] I5;
	input [31:0] I6;
	input [31:0] I7;
	input [31:0] I8;
	input [31:0] I9;
	input [31:0] I10;
	input [31:0] I11;
	input [31:0] I12;
	input [31:0] I13;
	input [31:0] I14;
	input [31:0] I15;
	input [3:0] S;
	output [31:0] O0;




	notech_inv i_7696(.A(n_54998), .Z(n_55283));
	notech_inv i_7691(.A(n_54998), .Z(n_55278));
	notech_inv i_7686(.A(n_54987), .Z(n_55272));
	notech_inv i_7681(.A(n_54987), .Z(n_55267));
	notech_inv i_7445(.A(n_55020), .Z(n_55021));
	notech_inv i_7444(.A(n_18765), .Z(n_55020));
	notech_inv i_7442(.A(n_723), .Z(n_55017));
	notech_inv i_7440(.A(n_723), .Z(n_55015));
	notech_inv i_7437(.A(n_723), .Z(n_55012));
	notech_inv i_7435(.A(n_723), .Z(n_55010));
	notech_inv i_7425(.A(n_54998), .Z(n_54999));
	notech_inv i_7424(.A(n_548), .Z(n_54998));
	notech_inv i_7415(.A(n_54987), .Z(n_54988));
	notech_inv i_7414(.A(n_549), .Z(n_54987));
	notech_inv i_180(.A(S[3]), .Z(n_723));
	notech_inv i_179(.A(n_722), .Z(n_684));
	notech_inv i_178(.A(S[2]), .Z(n_722));
	notech_mux4 i_67(.S0(n_548), .S1(n_549), .A(I4[31]), .B(I5[31]), .C(I6[
		31]), .D(I7[31]), .Z(n_615));
	notech_mux4 i_66(.S0(n_548), .S1(n_549), .A(I4[30]), .B(I5[30]), .C(I6[
		30]), .D(I7[30]), .Z(n_614));
	notech_mux4 i_65(.S0(n_548), .S1(n_549), .A(I4[29]), .B(I5[29]), .C(I6[
		29]), .D(I7[29]), .Z(n_613));
	notech_mux4 i_64(.S0(n_548), .S1(n_549), .A(I4[28]), .B(I5[28]), .C(I6[
		28]), .D(I7[28]), .Z(n_612));
	notech_mux4 i_63(.S0(n_548), .S1(n_549), .A(I4[27]), .B(I5[27]), .C(I6[
		27]), .D(I7[27]), .Z(n_611));
	notech_mux4 i_62(.S0(n_548), .S1(n_549), .A(I4[26]), .B(I5[26]), .C(I6[
		26]), .D(I7[26]), .Z(n_610));
	notech_mux4 i_61(.S0(n_548), .S1(n_549), .A(I4[25]), .B(I5[25]), .C(I6[
		25]), .D(I7[25]), .Z(n_609));
	notech_mux4 i_60(.S0(n_548), .S1(n_549), .A(I4[24]), .B(I5[24]), .C(I6[
		24]), .D(I7[24]), .Z(n_608));
	notech_mux4 i_59(.S0(n_548), .S1(n_549), .A(I4[23]), .B(I5[23]), .C(I6[
		23]), .D(I7[23]), .Z(n_607));
	notech_mux4 i_58(.S0(n_548), .S1(n_549), .A(I4[22]), .B(I5[22]), .C(I6[
		22]), .D(I7[22]), .Z(n_606));
	notech_mux4 i_57(.S0(n_548), .S1(n_549), .A(I4[21]), .B(I5[21]), .C(I6[
		21]), .D(I7[21]), .Z(n_605));
	notech_mux4 i_56(.S0(n_548), .S1(n_549), .A(I4[20]), .B(I5[20]), .C(I6[
		20]), .D(I7[20]), .Z(n_604));
	notech_mux4 i_55(.S0(n_548), .S1(n_549), .A(I4[19]), .B(I5[19]), .C(I6[
		19]), .D(I7[19]), .Z(n_603));
	notech_mux4 i_54(.S0(n_548), .S1(n_549), .A(I4[18]), .B(I5[18]), .C(I6[
		18]), .D(I7[18]), .Z(n_602));
	notech_mux4 i_53(.S0(n_548), .S1(n_549), .A(I4[17]), .B(I5[17]), .C(I6[
		17]), .D(I7[17]), .Z(n_601));
	notech_mux4 i_52(.S0(n_548), .S1(n_549), .A(I4[16]), .B(I5[16]), .C(I6[
		16]), .D(I7[16]), .Z(n_600));
	notech_mux4 i_51(.S0(n_54999), .S1(n_54988), .A(I4[15]), .B(I5[15]), .C(I6
		[15]), .D(I7[15]), .Z(n_599));
	notech_mux4 i_50(.S0(n_54999), .S1(n_54988), .A(I4[14]), .B(I5[14]), .C(I6
		[14]), .D(I7[14]), .Z(n_598));
	notech_mux4 i_49(.S0(n_54999), .S1(n_54988), .A(I4[13]), .B(I5[13]), .C(I6
		[13]), .D(I7[13]), .Z(n_597));
	notech_mux4 i_48(.S0(n_54999), .S1(n_54988), .A(I4[12]), .B(I5[12]), .C(I6
		[12]), .D(I7[12]), .Z(n_596));
	notech_mux4 i_47(.S0(n_54999), .S1(n_54988), .A(I4[11]), .B(I5[11]), .C(I6
		[11]), .D(I7[11]), .Z(n_595));
	notech_mux4 i_46(.S0(n_54999), .S1(n_54988), .A(I4[10]), .B(I5[10]), .C(I6
		[10]), .D(I7[10]), .Z(n_594));
	notech_mux4 i_45(.S0(n_54999), .S1(n_54988), .A(I4[9]), .B(I5[9]), .C(I6
		[9]), .D(I7[9]), .Z(n_593));
	notech_mux4 i_44(.S0(n_54999), .S1(n_54988), .A(I4[8]), .B(I5[8]), .C(I6
		[8]), .D(I7[8]), .Z(n_592));
	notech_mux4 i_43(.S0(n_54999), .S1(n_54988), .A(I4[7]), .B(I5[7]), .C(I6
		[7]), .D(I7[7]), .Z(n_591));
	notech_mux4 i_42(.S0(n_54999), .S1(n_54988), .A(I4[6]), .B(I5[6]), .C(I6
		[6]), .D(I7[6]), .Z(n_590));
	notech_mux4 i_41(.S0(n_54999), .S1(n_54988), .A(I4[5]), .B(I5[5]), .C(I6
		[5]), .D(I7[5]), .Z(n_589));
	notech_mux4 i_40(.S0(n_54999), .S1(n_54988), .A(I4[4]), .B(I5[4]), .C(I6
		[4]), .D(I7[4]), .Z(n_588));
	notech_mux4 i_39(.S0(n_54999), .S1(n_54988), .A(I4[3]), .B(I5[3]), .C(I6
		[3]), .D(I7[3]), .Z(n_587));
	notech_mux4 i_38(.S0(n_54999), .S1(n_54988), .A(I4[2]), .B(I5[2]), .C(I6
		[2]), .D(I7[2]), .Z(n_586));
	notech_mux4 i_37(.S0(n_54999), .S1(n_54988), .A(I4[1]), .B(I5[1]), .C(I6
		[1]), .D(I7[1]), .Z(n_585));
	notech_mux4 i_36(.S0(n_54999), .S1(n_54988), .A(I4[0]), .B(I5[0]), .C(I6
		[0]), .D(I7[0]), .Z(n_584));
	notech_mux4 i_33(.S0(n_55278), .S1(n_55267), .A(I0[31]), .B(I1[31]), .C(I2
		[31]), .D(I3[31]), .Z(n_581));
	notech_mux4 i_32(.S0(n_55278), .S1(n_55267), .A(I0[30]), .B(I1[30]), .C(I2
		[30]), .D(I3[30]), .Z(n_580));
	notech_mux4 i_31(.S0(n_55278), .S1(n_55267), .A(I0[29]), .B(I1[29]), .C(I2
		[29]), .D(I3[29]), .Z(n_579));
	notech_mux4 i_30(.S0(n_55278), .S1(n_55267), .A(I0[28]), .B(I1[28]), .C(I2
		[28]), .D(I3[28]), .Z(n_578));
	notech_mux4 i_29(.S0(n_55278), .S1(n_55267), .A(I0[27]), .B(I1[27]), .C(I2
		[27]), .D(I3[27]), .Z(n_577));
	notech_mux4 i_28(.S0(n_55278), .S1(n_55267), .A(I0[26]), .B(I1[26]), .C(I2
		[26]), .D(I3[26]), .Z(n_576));
	notech_mux4 i_27(.S0(n_55278), .S1(n_55267), .A(I0[25]), .B(I1[25]), .C(I2
		[25]), .D(I3[25]), .Z(n_575));
	notech_mux4 i_26(.S0(n_55278), .S1(n_55267), .A(I0[24]), .B(I1[24]), .C(I2
		[24]), .D(I3[24]), .Z(n_574));
	notech_mux4 i_25(.S0(n_55278), .S1(n_55267), .A(I0[23]), .B(I1[23]), .C(I2
		[23]), .D(I3[23]), .Z(n_573));
	notech_mux4 i_24(.S0(n_55278), .S1(n_55267), .A(I0[22]), .B(I1[22]), .C(I2
		[22]), .D(I3[22]), .Z(n_572));
	notech_mux4 i_23(.S0(n_55278), .S1(n_55267), .A(I0[21]), .B(I1[21]), .C(I2
		[21]), .D(I3[21]), .Z(n_571));
	notech_mux4 i_22(.S0(n_55278), .S1(n_55267), .A(I0[20]), .B(I1[20]), .C(I2
		[20]), .D(I3[20]), .Z(n_570));
	notech_mux4 i_21(.S0(n_55278), .S1(n_55267), .A(I0[19]), .B(I1[19]), .C(I2
		[19]), .D(I3[19]), .Z(n_569));
	notech_mux4 i_20(.S0(n_55278), .S1(n_55267), .A(I0[18]), .B(I1[18]), .C(I2
		[18]), .D(I3[18]), .Z(n_568));
	notech_mux4 i_19(.S0(n_55278), .S1(n_55267), .A(I0[17]), .B(I1[17]), .C(I2
		[17]), .D(I3[17]), .Z(n_567));
	notech_mux4 i_18(.S0(n_55278), .S1(n_55267), .A(I0[16]), .B(I1[16]), .C(I2
		[16]), .D(I3[16]), .Z(n_566));
	notech_mux4 i_17(.S0(n_55283), .S1(n_55272), .A(I0[15]), .B(I1[15]), .C(I2
		[15]), .D(I3[15]), .Z(n_565));
	notech_mux4 i_16(.S0(n_55283), .S1(n_55272), .A(I0[14]), .B(I1[14]), .C(I2
		[14]), .D(I3[14]), .Z(n_564));
	notech_mux4 i_15(.S0(n_55283), .S1(n_55272), .A(I0[13]), .B(I1[13]), .C(I2
		[13]), .D(I3[13]), .Z(n_563));
	notech_mux4 i_14(.S0(n_55283), .S1(n_55272), .A(I0[12]), .B(I1[12]), .C(I2
		[12]), .D(I3[12]), .Z(n_562));
	notech_mux4 i_13(.S0(n_55283), .S1(n_55272), .A(I0[11]), .B(I1[11]), .C(I2
		[11]), .D(I3[11]), .Z(n_561));
	notech_mux4 i_12(.S0(n_55283), .S1(n_55272), .A(I0[10]), .B(I1[10]), .C(I2
		[10]), .D(I3[10]), .Z(n_560));
	notech_mux4 i_11(.S0(n_55283), .S1(n_55272), .A(I0[9]), .B(I1[9]), .C(I2
		[9]), .D(I3[9]), .Z(n_559));
	notech_mux4 i_10(.S0(n_55283), .S1(n_55272), .A(I0[8]), .B(I1[8]), .C(I2
		[8]), .D(I3[8]), .Z(n_558));
	notech_mux4 i_9(.S0(n_55283), .S1(n_55272), .A(I0[7]), .B(I1[7]), .C(I2[
		7]), .D(I3[7]), .Z(n_557));
	notech_mux4 i_8(.S0(n_55283), .S1(n_55272), .A(I0[6]), .B(I1[6]), .C(I2[
		6]), .D(I3[6]), .Z(n_556));
	notech_mux4 i_7(.S0(n_55283), .S1(n_55272), .A(I0[5]), .B(I1[5]), .C(I2[
		5]), .D(I3[5]), .Z(n_555));
	notech_mux4 i_6(.S0(n_55283), .S1(n_55272), .A(I0[4]), .B(I1[4]), .C(I2[
		4]), .D(I3[4]), .Z(n_554));
	notech_mux4 i_5(.S0(n_55283), .S1(n_55272), .A(I0[3]), .B(I1[3]), .C(I2[
		3]), .D(I3[3]), .Z(n_553));
	notech_mux4 i_4(.S0(n_55283), .S1(n_55272), .A(I0[2]), .B(I1[2]), .C(I2[
		2]), .D(I3[2]), .Z(n_552));
	notech_mux4 i_3(.S0(n_55283), .S1(n_55272), .A(I0[1]), .B(I1[1]), .C(I2[
		1]), .D(I3[1]), .Z(n_551));
	notech_mux4 i_2(.S0(n_55283), .S1(n_55272), .A(I0[0]), .B(I1[0]), .C(I2[
		0]), .D(I3[0]), .Z(n_550));
	notech_inv i_173(.A(n_719), .Z(n_549));
	notech_inv i_172(.A(S[1]), .Z(n_719));
	notech_inv i_171(.A(n_718), .Z(n_548));
	notech_inv i_170(.A(S[0]), .Z(n_718));
	notech_nand2 i_28199(.A(n_18003), .B(n_18006), .Z(O0[0]));
	notech_nao3 i_28191(.A(n_55020), .B(n_584), .C(n_55012), .Z(n_18006));
	notech_nao3 i_28188(.A(n_550), .B(n_18765), .C(n_55012), .Z(n_18003));
	notech_nand2 i_5098337(.A(n_18027), .B(n_18030), .Z(O0[1]));
	notech_nao3 i_4298338(.A(n_55020), .B(n_585), .C(n_55012), .Z(n_18030)
		);
	notech_nao3 i_3998339(.A(n_551), .B(n_55021), .C(n_55012), .Z(n_18027)
		);
	notech_nand2 i_5098341(.A(n_18051), .B(n_18054), .Z(O0[2]));
	notech_nao3 i_4298342(.A(n_55020), .B(n_586), .C(n_55012), .Z(n_18054)
		);
	notech_nao3 i_3998343(.A(n_552), .B(n_18765), .C(n_55012), .Z(n_18051)
		);
	notech_nand2 i_5098345(.A(n_18075), .B(n_18078), .Z(O0[3]));
	notech_nao3 i_4298346(.A(n_55020), .B(n_587), .C(n_55012), .Z(n_18078)
		);
	notech_nao3 i_3998347(.A(n_553), .B(n_55021), .C(n_55012), .Z(n_18075)
		);
	notech_nand2 i_5098349(.A(n_18099), .B(n_18102), .Z(O0[4]));
	notech_nao3 i_4298350(.A(n_55020), .B(n_588), .C(n_55012), .Z(n_18102)
		);
	notech_nao3 i_3998351(.A(n_554), .B(n_18765), .C(n_55012), .Z(n_18099)
		);
	notech_nand2 i_5098353(.A(n_18123), .B(n_18126), .Z(O0[5]));
	notech_nao3 i_4298354(.A(n_684), .B(n_589), .C(n_55012), .Z(n_18126));
	notech_nao3 i_3998355(.A(n_555), .B(n_55021), .C(n_55012), .Z(n_18123)
		);
	notech_nand2 i_5098357(.A(n_18147), .B(n_18150), .Z(O0[6]));
	notech_nao3 i_4298358(.A(n_55020), .B(n_590), .C(n_55012), .Z(n_18150)
		);
	notech_nao3 i_3998359(.A(n_556), .B(n_18765), .C(n_55012), .Z(n_18147)
		);
	notech_nand2 i_5098361(.A(n_18171), .B(n_18174), .Z(O0[7]));
	notech_nao3 i_4298362(.A(n_55020), .B(n_591), .C(n_55012), .Z(n_18174)
		);
	notech_nao3 i_3998363(.A(n_557), .B(n_55021), .C(n_55012), .Z(n_18171)
		);
	notech_nand2 i_5098365(.A(n_18195), .B(n_18198), .Z(O0[8]));
	notech_nao3 i_4298366(.A(n_55020), .B(n_592), .C(n_55010), .Z(n_18198)
		);
	notech_nao3 i_3998367(.A(n_558), .B(n_18765), .C(n_55010), .Z(n_18195)
		);
	notech_nand2 i_5098369(.A(n_18219), .B(n_18222), .Z(O0[9]));
	notech_nao3 i_4298370(.A(n_55020), .B(n_593), .C(n_55010), .Z(n_18222)
		);
	notech_nao3 i_3998371(.A(n_559), .B(n_55021), .C(n_55010), .Z(n_18219)
		);
	notech_nand2 i_5098373(.A(n_18243), .B(n_18246), .Z(O0[10]));
	notech_nao3 i_4298374(.A(n_55020), .B(n_594), .C(n_55010), .Z(n_18246)
		);
	notech_nao3 i_3998375(.A(n_560), .B(n_18765), .C(n_55010), .Z(n_18243)
		);
	notech_nand2 i_5098377(.A(n_18267), .B(n_18270), .Z(O0[11]));
	notech_nao3 i_4298378(.A(n_55020), .B(n_595), .C(n_55010), .Z(n_18270)
		);
	notech_nao3 i_3998379(.A(n_561), .B(n_55021), .C(n_55010), .Z(n_18267)
		);
	notech_nand2 i_5098381(.A(n_18291), .B(n_18294), .Z(O0[12]));
	notech_nao3 i_4298382(.A(n_55020), .B(n_596), .C(n_55010), .Z(n_18294)
		);
	notech_nao3 i_3998383(.A(n_562), .B(n_18765), .C(n_55010), .Z(n_18291)
		);
	notech_nand2 i_5098385(.A(n_18315), .B(n_18318), .Z(O0[13]));
	notech_nao3 i_4298386(.A(n_55020), .B(n_597), .C(n_55010), .Z(n_18318)
		);
	notech_nao3 i_3998387(.A(n_563), .B(n_55021), .C(n_55010), .Z(n_18315)
		);
	notech_nand2 i_5098389(.A(n_18339), .B(n_18342), .Z(O0[14]));
	notech_nao3 i_4298390(.A(n_55020), .B(n_598), .C(n_55010), .Z(n_18342)
		);
	notech_nao3 i_3998391(.A(n_564), .B(n_18765), .C(n_55010), .Z(n_18339)
		);
	notech_nand2 i_5098393(.A(n_18363), .B(n_18366), .Z(O0[15]));
	notech_nao3 i_4298394(.A(n_55020), .B(n_599), .C(n_55010), .Z(n_18366)
		);
	notech_nao3 i_3998395(.A(n_565), .B(n_55021), .C(n_55010), .Z(n_18363)
		);
	notech_nand2 i_5098397(.A(n_18387), .B(n_18390), .Z(O0[16]));
	notech_nao3 i_4298398(.A(n_684), .B(n_600), .C(n_55017), .Z(n_18390));
	notech_nao3 i_3998399(.A(n_566), .B(n_18765), .C(n_55017), .Z(n_18387)
		);
	notech_nand2 i_5098401(.A(n_18411), .B(n_18414), .Z(O0[17]));
	notech_nao3 i_4298402(.A(n_684), .B(n_601), .C(n_55017), .Z(n_18414));
	notech_nao3 i_3998403(.A(n_567), .B(n_55021), .C(n_55017), .Z(n_18411)
		);
	notech_nand2 i_5098405(.A(n_18435), .B(n_18438), .Z(O0[18]));
	notech_nao3 i_4298406(.A(n_684), .B(n_602), .C(n_55017), .Z(n_18438));
	notech_nao3 i_3998407(.A(n_568), .B(n_18765), .C(n_55017), .Z(n_18435)
		);
	notech_nand2 i_5098409(.A(n_18459), .B(n_18462), .Z(O0[19]));
	notech_nao3 i_4298410(.A(n_684), .B(n_603), .C(n_55017), .Z(n_18462));
	notech_nao3 i_3998411(.A(n_569), .B(n_55021), .C(n_55017), .Z(n_18459)
		);
	notech_nand2 i_5098413(.A(n_18483), .B(n_18486), .Z(O0[20]));
	notech_nao3 i_4298414(.A(n_684), .B(n_604), .C(n_55017), .Z(n_18486));
	notech_nao3 i_3998415(.A(n_570), .B(n_18765), .C(n_55017), .Z(n_18483)
		);
	notech_nand2 i_5098417(.A(n_18507), .B(n_18510), .Z(O0[21]));
	notech_nao3 i_4298418(.A(n_684), .B(n_605), .C(n_55017), .Z(n_18510));
	notech_nao3 i_3998419(.A(n_571), .B(n_18765), .C(n_55017), .Z(n_18507)
		);
	notech_nand2 i_5098421(.A(n_18531), .B(n_18534), .Z(O0[22]));
	notech_nao3 i_4298422(.A(n_684), .B(n_606), .C(n_55017), .Z(n_18534));
	notech_nao3 i_3998423(.A(n_572), .B(n_18765), .C(n_55017), .Z(n_18531)
		);
	notech_nand2 i_5098425(.A(n_18555), .B(n_18558), .Z(O0[23]));
	notech_nao3 i_4298426(.A(n_684), .B(n_607), .C(n_55017), .Z(n_18558));
	notech_nao3 i_3998427(.A(n_573), .B(n_55021), .C(n_55017), .Z(n_18555)
		);
	notech_nand2 i_5098429(.A(n_18579), .B(n_18582), .Z(O0[24]));
	notech_nao3 i_4298430(.A(n_684), .B(n_608), .C(n_55015), .Z(n_18582));
	notech_nao3 i_3998431(.A(n_574), .B(n_18765), .C(n_55015), .Z(n_18579)
		);
	notech_nand2 i_5098433(.A(n_18603), .B(n_18606), .Z(O0[25]));
	notech_nao3 i_4298434(.A(n_684), .B(n_609), .C(n_55015), .Z(n_18606));
	notech_nao3 i_3998435(.A(n_575), .B(n_55021), .C(n_55015), .Z(n_18603)
		);
	notech_nand2 i_5098437(.A(n_18627), .B(n_18630), .Z(O0[26]));
	notech_nao3 i_4298438(.A(n_684), .B(n_610), .C(n_55015), .Z(n_18630));
	notech_nao3 i_3998439(.A(n_576), .B(n_18765), .C(n_55015), .Z(n_18627)
		);
	notech_nand2 i_5098441(.A(n_18651), .B(n_18654), .Z(O0[27]));
	notech_nao3 i_4298442(.A(n_684), .B(n_611), .C(n_55015), .Z(n_18654));
	notech_nao3 i_3998443(.A(n_577), .B(n_55021), .C(n_55015), .Z(n_18651)
		);
	notech_nand2 i_5098445(.A(n_18675), .B(n_18678), .Z(O0[28]));
	notech_nao3 i_4298446(.A(n_684), .B(n_612), .C(n_55015), .Z(n_18678));
	notech_nao3 i_3998447(.A(n_578), .B(n_18765), .C(n_55015), .Z(n_18675)
		);
	notech_nand2 i_5098449(.A(n_18699), .B(n_18702), .Z(O0[29]));
	notech_nao3 i_4298450(.A(n_684), .B(n_613), .C(n_55015), .Z(n_18702));
	notech_nao3 i_3998451(.A(n_579), .B(n_55021), .C(n_55015), .Z(n_18699)
		);
	notech_nand2 i_5098453(.A(n_18723), .B(n_18726), .Z(O0[30]));
	notech_nao3 i_4298454(.A(n_684), .B(n_614), .C(n_55015), .Z(n_18726));
	notech_nao3 i_3998455(.A(n_580), .B(n_18765), .C(n_55015), .Z(n_18723)
		);
	notech_inv i_398456(.A(n_684), .Z(n_18765));
	notech_nand2 i_5098457(.A(n_18747), .B(n_18750), .Z(O0[31]));
	notech_nao3 i_4298458(.A(n_684), .B(n_615), .C(n_55015), .Z(n_18750));
	notech_nao3 i_3998459(.A(n_581), .B(n_55021), .C(n_55015), .Z(n_18747)
		);
endmodule
module AWMUX_16_32_3(I0 , I1 , I2 , I3 , I4 , I5 , I6 , I7 , I8 , I9 , I10 , I11 , I12 , I13 , I14 , I15 , S , O0);
input  [31:0] I0;
input  [31:0] I1;
input  [31:0] I2;
input  [31:0] I3;
input  [31:0] I4;
input  [31:0] I5;
input  [31:0] I6;
input  [31:0] I7;
input  [31:0] I8;
input  [31:0] I9;
input  [31:0] I10;
input  [31:0] I11;
input  [31:0] I12;
input  [31:0] I13;
input  [31:0] I14;
input  [31:0] I15;
input  [3:0] S;
output  [31:0] O0;
reg [31:0] O0;

always @(I0 or I1 or I2 or I3 or I4 or I5 or I6 or I7 or I8 or I9 or I10 or I11 or I12 or I13 or I14 or I15 or S or O0)
begin
	case(S)
	4'h0 : O0 = I0;
	4'h1 : O0 = I1;
	4'h2 : O0 = I2;
	4'h3 : O0 = I3;
	4'h4 : O0 = I4;
	4'h5 : O0 = I5;
	4'h6 : O0 = I6;
	4'h7 : O0 = I7;
	4'h8 : O0 = I8;
	4'h9 : O0 = I9;
	4'ha : O0 = I10;
	4'hb : O0 = I11;
	4'hc : O0 = I12;
	4'hd : O0 = I13;
	4'he : O0 = I14;
	default : O0 = I15;
	endcase
end
endmodule

module AWMUX_16_32_4(I0 , I1 , I2 , I3 , I4 , I5 , I6 , I7 , I8 , I9 , I10 , I11 , I12 , I13 , I14 , I15 , S , O0);
input  [31:0] I0;
input  [31:0] I1;
input  [31:0] I2;
input  [31:0] I3;
input  [31:0] I4;
input  [31:0] I5;
input  [31:0] I6;
input  [31:0] I7;
input  [31:0] I8;
input  [31:0] I9;
input  [31:0] I10;
input  [31:0] I11;
input  [31:0] I12;
input  [31:0] I13;
input  [31:0] I14;
input  [31:0] I15;
input  [3:0] S;
output  [31:0] O0;
reg [31:0] O0;

always @(I0 or I1 or I2 or I3 or I4 or I5 or I6 or I7 or I8 or I9 or I10 or I11 or I12 or I13 or I14 or I15 or S or O0)
begin
	case(S)
	4'h0 : O0 = I0;
	4'h1 : O0 = I1;
	4'h2 : O0 = I2;
	4'h3 : O0 = I3;
	4'h4 : O0 = I4;
	4'h5 : O0 = I5;
	4'h6 : O0 = I6;
	4'h7 : O0 = I7;
	4'h8 : O0 = I8;
	4'h9 : O0 = I9;
	4'ha : O0 = I10;
	4'hb : O0 = I11;
	4'hc : O0 = I12;
	4'hd : O0 = I13;
	4'he : O0 = I14;
	default : O0 = I15;
	endcase
end
endmodule

module AWMUX_16_32_5(I0 , I1 , I2 , I3 , I4 , I5 , I6 , I7 , I8 , I9 , I10 , I11 , I12 , I13 , I14 , I15 , S , O0);
input  [31:0] I0;
input  [31:0] I1;
input  [31:0] I2;
input  [31:0] I3;
input  [31:0] I4;
input  [31:0] I5;
input  [31:0] I6;
input  [31:0] I7;
input  [31:0] I8;
input  [31:0] I9;
input  [31:0] I10;
input  [31:0] I11;
input  [31:0] I12;
input  [31:0] I13;
input  [31:0] I14;
input  [31:0] I15;
input  [3:0] S;
output  [31:0] O0;
reg [31:0] O0;

always @(I0 or I1 or I2 or I3 or I4 or I5 or I6 or I7 or I8 or I9 or I10 or I11 or I12 or I13 or I14 or I15 or S or O0)
begin
	case(S)
	4'h0 : O0 = I0;
	4'h1 : O0 = I1;
	4'h2 : O0 = I2;
	4'h3 : O0 = I3;
	4'h4 : O0 = I4;
	4'h5 : O0 = I5;
	4'h6 : O0 = I6;
	4'h7 : O0 = I7;
	4'h8 : O0 = I8;
	4'h9 : O0 = I9;
	4'ha : O0 = I10;
	4'hb : O0 = I11;
	4'hc : O0 = I12;
	4'hd : O0 = I13;
	4'he : O0 = I14;
	default : O0 = I15;
	endcase
end
endmodule

module AWMUX_16_32_6(I0 , I1 , I2 , I3 , I4 , I5 , I6 , I7 , I8 , I9 , I10 , I11 , I12 , I13 , I14 , I15 , S , O0);
input  [31:0] I0;
input  [31:0] I1;
input  [31:0] I2;
input  [31:0] I3;
input  [31:0] I4;
input  [31:0] I5;
input  [31:0] I6;
input  [31:0] I7;
input  [31:0] I8;
input  [31:0] I9;
input  [31:0] I10;
input  [31:0] I11;
input  [31:0] I12;
input  [31:0] I13;
input  [31:0] I14;
input  [31:0] I15;
input  [3:0] S;
output  [31:0] O0;
reg [31:0] O0;

always @(I0 or I1 or I2 or I3 or I4 or I5 or I6 or I7 or I8 or I9 or I10 or I11 or I12 or I13 or I14 or I15 or S or O0)
begin
	case(S)
	4'h0 : O0 = I0;
	4'h1 : O0 = I1;
	4'h2 : O0 = I2;
	4'h3 : O0 = I3;
	4'h4 : O0 = I4;
	4'h5 : O0 = I5;
	4'h6 : O0 = I6;
	4'h7 : O0 = I7;
	4'h8 : O0 = I8;
	4'h9 : O0 = I9;
	4'ha : O0 = I10;
	4'hb : O0 = I11;
	4'hc : O0 = I12;
	4'hd : O0 = I13;
	4'he : O0 = I14;
	default : O0 = I15;
	endcase
end
endmodule

module AWMUX_16_32_7(I0 , I1 , I2 , I3 , I4 , I5 , I6 , I7 , I8 , I9 , I10 , I11 , I12 , I13 , I14 , I15 , S , O0);
input  [31:0] I0;
input  [31:0] I1;
input  [31:0] I2;
input  [31:0] I3;
input  [31:0] I4;
input  [31:0] I5;
input  [31:0] I6;
input  [31:0] I7;
input  [31:0] I8;
input  [31:0] I9;
input  [31:0] I10;
input  [31:0] I11;
input  [31:0] I12;
input  [31:0] I13;
input  [31:0] I14;
input  [31:0] I15;
input  [3:0] S;
output  [31:0] O0;
reg [31:0] O0;

always @(I0 or I1 or I2 or I3 or I4 or I5 or I6 or I7 or I8 or I9 or I10 or I11 or I12 or I13 or I14 or I15 or S or O0)
begin
	case(S)
	4'h0 : O0 = I0;
	4'h1 : O0 = I1;
	4'h2 : O0 = I2;
	4'h3 : O0 = I3;
	4'h4 : O0 = I4;
	4'h5 : O0 = I5;
	4'h6 : O0 = I6;
	4'h7 : O0 = I7;
	4'h8 : O0 = I8;
	4'h9 : O0 = I9;
	4'ha : O0 = I10;
	4'hb : O0 = I11;
	4'hc : O0 = I12;
	4'hd : O0 = I13;
	4'he : O0 = I14;
	default : O0 = I15;
	endcase
end
endmodule

module vliw(clk, rstn, instrc, ie, readio_data, io_add, writeio_data, writeio_req
		, readio_req, writeio_ack, readio_ack, read_reqs, read_ack, read_data
		, over_seg, cr3, cr2, icr2, cr1, cr0, write_reqs, write_ack, write_data
		, Daddr, write_sz, read_sz, cs, add_src, from_acu, to_acu, seg_src
		, pg_en, ready_vliw, valid_op, imm, lenpc, pc_out, pc_req, opz, reps
		, adz, flush_tlb, flush_Dtlb, terminate, start_up, pg_fault, ipg_fault
		, wr_fault, pt_fault, repbytecache);

	input clk;
	input rstn;
	input [127:0] instrc;
	output ie;
	input [31:0] readio_data;
	output [31:0] io_add;
	output [31:0] writeio_data;
	output writeio_req;
	output readio_req;
	input writeio_ack;
	input readio_ack;
	output read_reqs;
	input read_ack;
	input [31:0] read_data;
	input [5:0] over_seg;
	output [31:0] cr3;
	input [31:0] cr2;
	input [31:0] icr2;
	output [31:0] cr1;
	output [31:0] cr0;
	output write_reqs;
	input write_ack;
	output [31:0] write_data;
	output [31:0] Daddr;
	output [1:0] write_sz;
	output [1:0] read_sz;
	output [31:0] cs;
	input [31:0] add_src;
	input [7:0] from_acu;
	output [63:0] to_acu;
	input [2:0] seg_src;
	output pg_en;
	output ready_vliw;
	input valid_op;
	input [63:0] imm;
	input [31:0] lenpc;
	output [31:0] pc_out;
	output pc_req;
	input [2:0] opz;
	input [2:0] reps;
	input adz;
	output flush_tlb;
	output flush_Dtlb;
	output terminate;
	input start_up;
	input pg_fault;
	input ipg_fault;
	input wr_fault;
	input pt_fault;
	output repbytecache;

	wire [4:0] fsm;
	wire [31:0] opa;
	wire [31:0] opb;
	wire [31:0] nbus_11271;
	wire [31:0] opc;
	wire [31:0] opd;
	wire [15:0] nbus_11273;
	wire [31:0] gs;
	wire [31:0] sav_ecx;
	wire [31:0] sav_edi;
	wire [31:0] sav_esi;
	wire [31:0] sav_esp;
	wire [31:0] temp_sp;
	wire [1:0] sav_cs;
	wire [31:0] cr2_reg;
	wire [31:0] nbus_14541;
	wire [4:0] vliw_pc;
	wire [31:0] temp_ss;
	wire [31:0] errco;
	wire [31:0] sav_epc;
	wire [2:0] mask8b;
	wire [1:0] pipe_mul;
	wire [4:0] fsmf;
	wire [31:0] Daddrgs;
	wire [63:0] to_acu101153;
	wire [31:0] nbus_11346;
	wire [31:0] nbus_11291;
	wire [31:0] nbus_11270;
	wire [31:0] Daddrs_8;
	wire [31:0] write_data_33;
	wire [31:0] write_data_32;
	wire [31:0] write_data_31;
	wire [31:0] write_data_30;
	wire [31:0] write_data_29;
	wire [31:0] write_data_28;
	wire [31:0] write_data_27;
	wire [31:0] write_data_26;
	wire [31:0] write_data_25;
	wire [31:0] opc_14;
	wire [31:0] opc_10;
	wire [31:0] Daddrs_3;
	wire [31:0] Daddrs_1;
	wire [63:0] divr_1;
	wire [31:0] regs_4_2;
	wire [31:0] opa_0;
	wire [31:0] resa_arithbox;
	wire [16:0] nbus_143;
	wire [32:0] nbus_142;
	wire [16:0] nbus_141;
	wire [32:0] nbus_140;
	wire [16:0] nbus_139;
	wire [32:0] nbus_138;
	wire [16:0] nbus_137;
	wire [32:0] nbus_136;
	wire [8:0] nbus_135;
	wire [16:0] nbus_134;
	wire [32:0] nbus_133;
	wire [63:0] mul64;
	wire [31:0] add_len_pc32;
	wire [31:0] resb_shift4box;
	wire [31:0] resa_shift4box;
	wire [31:0] resb_shiftbox;
	wire [31:0] resa_shiftbox;
	wire [3:0] calc_sz;
	wire [63:0] tsc;
	wire [3:0] all_cnt;
	wire [31:0] regs_14;
	wire [31:0] regs_12;
	wire [31:0] regs_11;
	wire [31:0] regs_10;
	wire [31:0] regs_8;
	wire [31:0] regs_7;
	wire [31:0] regs_6;
	wire [31:0] regs_5;
	wire [31:0] regs_4;
	wire [31:0] regs_3;
	wire [31:0] regs_2;
	wire [31:0] ecx;
	wire [63:0] divq;
	wire [63:0] divr;
	wire [31:0] regs_0;
	wire [31:0] ldtr;
	wire [31:0] gdtr;
	wire [31:0] idtr;
	wire [31:0] desc;



	notech_inv i_15650(.A(n_63817), .Z(n_63818));
	notech_inv i_15649(.A(\opcode[0] ), .Z(n_63817));
	notech_inv i_15632(.A(n_63799), .Z(n_63800));
	notech_inv i_15631(.A(\opcode[3] ), .Z(n_63799));
	notech_inv i_15628(.A(n_63795), .Z(n_63796));
	notech_inv i_15627(.A(n_63786), .Z(n_63795));
	notech_inv i_15626(.A(n_63793), .Z(n_63794));
	notech_inv i_15625(.A(n_63778), .Z(n_63793));
	notech_inv i_15624(.A(n_63791), .Z(n_63792));
	notech_inv i_15623(.A(n_63772), .Z(n_63791));
	notech_inv i_15622(.A(n_63789), .Z(n_63790));
	notech_inv i_15621(.A(n_63768), .Z(n_63789));
	notech_inv i_15620(.A(n_63787), .Z(n_63788));
	notech_inv i_15619(.A(n_63766), .Z(n_63787));
	notech_inv i_15618(.A(n_63785), .Z(n_63786));
	notech_inv i_15617(.A(n_63788), .Z(n_63785));
	notech_inv i_15616(.A(n_63783), .Z(n_63784));
	notech_inv i_15615(.A(n_63760), .Z(n_63783));
	notech_inv i_15614(.A(n_63781), .Z(n_63782));
	notech_inv i_15613(.A(n_63756), .Z(n_63781));
	notech_inv i_15612(.A(n_63779), .Z(n_63780));
	notech_inv i_15611(.A(n_63754), .Z(n_63779));
	notech_inv i_15610(.A(n_63777), .Z(n_63778));
	notech_inv i_15609(.A(n_63780), .Z(n_63777));
	notech_inv i_15608(.A(n_63775), .Z(n_63776));
	notech_inv i_15607(.A(n_63748), .Z(n_63775));
	notech_inv i_15606(.A(n_63773), .Z(n_63774));
	notech_inv i_15605(.A(n_63744), .Z(n_63773));
	notech_inv i_15604(.A(n_63771), .Z(n_63772));
	notech_inv i_15603(.A(n_63774), .Z(n_63771));
	notech_inv i_15602(.A(n_63769), .Z(n_63770));
	notech_inv i_15601(.A(n_63740), .Z(n_63769));
	notech_inv i_15600(.A(n_63767), .Z(n_63768));
	notech_inv i_15599(.A(n_63770), .Z(n_63767));
	notech_inv i_15598(.A(n_63765), .Z(n_63766));
	notech_inv i_15597(.A(n_63790), .Z(n_63765));
	notech_inv i_15596(.A(n_63763), .Z(n_63764));
	notech_inv i_15595(.A(n_63734), .Z(n_63763));
	notech_inv i_15594(.A(n_63761), .Z(n_63762));
	notech_inv i_15593(.A(n_63732), .Z(n_63761));
	notech_inv i_15592(.A(n_63759), .Z(n_63760));
	notech_inv i_15591(.A(n_63762), .Z(n_63759));
	notech_inv i_15590(.A(n_63757), .Z(n_63758));
	notech_inv i_15589(.A(n_63730), .Z(n_63757));
	notech_inv i_15588(.A(n_63755), .Z(n_63756));
	notech_inv i_15587(.A(n_63758), .Z(n_63755));
	notech_inv i_15586(.A(n_63753), .Z(n_63754));
	notech_inv i_15585(.A(n_63782), .Z(n_63753));
	notech_inv i_15584(.A(n_63751), .Z(n_63752));
	notech_inv i_15583(.A(n_63728), .Z(n_63751));
	notech_inv i_15580(.A(n_63747), .Z(n_63748));
	notech_inv i_15579(.A(n_63752), .Z(n_63747));
	notech_inv i_15576(.A(n_63743), .Z(n_63744));
	notech_inv i_15575(.A(n_63776), .Z(n_63743));
	notech_inv i_15572(.A(n_63739), .Z(n_63740));
	notech_inv i_15571(.A(n_63792), .Z(n_63739));
	notech_inv i_15568(.A(n_63735), .Z(n_63736));
	notech_inv i_15567(.A(\opcode[2] ), .Z(n_63735));
	notech_inv i_15566(.A(n_63733), .Z(n_63734));
	notech_inv i_15565(.A(n_63736), .Z(n_63733));
	notech_inv i_15564(.A(n_63731), .Z(n_63732));
	notech_inv i_15563(.A(n_63764), .Z(n_63731));
	notech_inv i_15562(.A(n_63729), .Z(n_63730));
	notech_inv i_15561(.A(n_63784), .Z(n_63729));
	notech_inv i_15560(.A(n_63727), .Z(n_63728));
	notech_inv i_15559(.A(n_63794), .Z(n_63727));
	notech_inv i_15552(.A(n_63719), .Z(n_63720));
	notech_inv i_15551(.A(n_63710), .Z(n_63719));
	notech_inv i_15550(.A(n_63717), .Z(n_63718));
	notech_inv i_15549(.A(n_63708), .Z(n_63717));
	notech_inv i_15548(.A(n_63715), .Z(n_63716));
	notech_inv i_15547(.A(n_63706), .Z(n_63715));
	notech_inv i_15544(.A(n_63711), .Z(n_63712));
	notech_inv i_15543(.A(n_63702), .Z(n_63711));
	notech_inv i_15542(.A(n_63709), .Z(n_63710));
	notech_inv i_15541(.A(n_63700), .Z(n_63709));
	notech_inv i_15540(.A(n_63707), .Z(n_63708));
	notech_inv i_15539(.A(n_63698), .Z(n_63707));
	notech_inv i_15538(.A(n_63705), .Z(n_63706));
	notech_inv i_15537(.A(n_63718), .Z(n_63705));
	notech_inv i_15534(.A(n_63701), .Z(n_63702));
	notech_inv i_15533(.A(\opcode[1] ), .Z(n_63701));
	notech_inv i_15532(.A(n_63699), .Z(n_63700));
	notech_inv i_15531(.A(n_63712), .Z(n_63699));
	notech_inv i_15530(.A(n_63697), .Z(n_63698));
	notech_inv i_15529(.A(n_63720), .Z(n_63697));
	notech_inv i_15526(.A(n_63693), .Z(n_63694));
	notech_inv i_15525(.A(n_63680), .Z(n_63693));
	notech_inv i_15524(.A(n_63691), .Z(n_63692));
	notech_inv i_15523(.A(n_63668), .Z(n_63691));
	notech_inv i_15522(.A(n_63689), .Z(n_63690));
	notech_inv i_15521(.A(n_63658), .Z(n_63689));
	notech_inv i_15520(.A(n_63687), .Z(n_63688));
	notech_inv i_15519(.A(n_63650), .Z(n_63687));
	notech_inv i_15518(.A(n_63685), .Z(n_63686));
	notech_inv i_15517(.A(n_63644), .Z(n_63685));
	notech_inv i_15516(.A(n_63683), .Z(n_63684));
	notech_inv i_15515(.A(n_63640), .Z(n_63683));
	notech_inv i_15514(.A(n_63681), .Z(n_63682));
	notech_inv i_15513(.A(n_63638), .Z(n_63681));
	notech_inv i_15512(.A(n_63679), .Z(n_63680));
	notech_inv i_15511(.A(n_63682), .Z(n_63679));
	notech_inv i_15508(.A(n_63675), .Z(n_63676));
	notech_inv i_15507(.A(n_63620), .Z(n_63675));
	notech_inv i_15506(.A(n_63673), .Z(n_63674));
	notech_inv i_15505(.A(n_63614), .Z(n_63673));
	notech_inv i_15504(.A(n_63671), .Z(n_63672));
	notech_inv i_15503(.A(n_63610), .Z(n_63671));
	notech_inv i_15502(.A(n_63669), .Z(n_63670));
	notech_inv i_15501(.A(n_63608), .Z(n_63669));
	notech_inv i_15500(.A(n_63667), .Z(n_63668));
	notech_inv i_15499(.A(n_63670), .Z(n_63667));
	notech_inv i_15498(.A(n_63665), .Z(n_63666));
	notech_inv i_15497(.A(n_63600), .Z(n_63665));
	notech_inv i_15496(.A(n_63663), .Z(n_63664));
	notech_inv i_15495(.A(n_63594), .Z(n_63663));
	notech_inv i_15494(.A(n_63661), .Z(n_63662));
	notech_inv i_15493(.A(n_63590), .Z(n_63661));
	notech_inv i_15492(.A(n_63659), .Z(n_63660));
	notech_inv i_15491(.A(n_63588), .Z(n_63659));
	notech_inv i_15490(.A(n_63657), .Z(n_63658));
	notech_inv i_15489(.A(n_63660), .Z(n_63657));
	notech_inv i_15488(.A(n_63655), .Z(n_63656));
	notech_inv i_15487(.A(n_63582), .Z(n_63655));
	notech_inv i_15486(.A(n_63653), .Z(n_63654));
	notech_inv i_15485(.A(n_63578), .Z(n_63653));
	notech_inv i_15484(.A(n_63651), .Z(n_63652));
	notech_inv i_15483(.A(n_63576), .Z(n_63651));
	notech_inv i_15482(.A(n_63649), .Z(n_63650));
	notech_inv i_15481(.A(n_63652), .Z(n_63649));
	notech_inv i_15480(.A(n_63647), .Z(n_63648));
	notech_inv i_15479(.A(n_63572), .Z(n_63647));
	notech_inv i_15478(.A(n_63645), .Z(n_63646));
	notech_inv i_15477(.A(n_63570), .Z(n_63645));
	notech_inv i_15476(.A(n_63643), .Z(n_63644));
	notech_inv i_15475(.A(n_63646), .Z(n_63643));
	notech_inv i_15474(.A(n_63641), .Z(n_63642));
	notech_inv i_15473(.A(n_63568), .Z(n_63641));
	notech_inv i_15472(.A(n_63639), .Z(n_63640));
	notech_inv i_15471(.A(n_63642), .Z(n_63639));
	notech_inv i_15470(.A(n_63637), .Z(n_63638));
	notech_inv i_15469(.A(n_63684), .Z(n_63637));
	notech_inv i_15458(.A(n_63625), .Z(n_63626));
	notech_inv i_15457(.A(n_63542), .Z(n_63625));
	notech_inv i_15456(.A(n_63623), .Z(n_63624));
	notech_inv i_15455(.A(n_63538), .Z(n_63623));
	notech_inv i_15454(.A(n_63621), .Z(n_63622));
	notech_inv i_15453(.A(n_63536), .Z(n_63621));
	notech_inv i_15452(.A(n_63619), .Z(n_63620));
	notech_inv i_15451(.A(n_63622), .Z(n_63619));
	notech_inv i_15450(.A(n_63617), .Z(n_63618));
	notech_inv i_15449(.A(n_63532), .Z(n_63617));
	notech_inv i_15448(.A(n_63615), .Z(n_63616));
	notech_inv i_15447(.A(n_63530), .Z(n_63615));
	notech_inv i_15446(.A(n_63613), .Z(n_63614));
	notech_inv i_15445(.A(n_63616), .Z(n_63613));
	notech_inv i_15444(.A(n_63611), .Z(n_63612));
	notech_inv i_15443(.A(n_63528), .Z(n_63611));
	notech_inv i_15442(.A(n_63609), .Z(n_63610));
	notech_inv i_15441(.A(n_63612), .Z(n_63609));
	notech_inv i_15440(.A(n_63607), .Z(n_63608));
	notech_inv i_15439(.A(n_63672), .Z(n_63607));
	notech_inv i_15438(.A(n_63605), .Z(n_63606));
	notech_inv i_15437(.A(n_63522), .Z(n_63605));
	notech_inv i_15436(.A(n_63603), .Z(n_63604));
	notech_inv i_15435(.A(n_63518), .Z(n_63603));
	notech_inv i_15434(.A(n_63601), .Z(n_63602));
	notech_inv i_15433(.A(n_63516), .Z(n_63601));
	notech_inv i_15432(.A(n_63599), .Z(n_63600));
	notech_inv i_15431(.A(n_63602), .Z(n_63599));
	notech_inv i_15430(.A(n_63597), .Z(n_63598));
	notech_inv i_15429(.A(n_63512), .Z(n_63597));
	notech_inv i_15428(.A(n_63595), .Z(n_63596));
	notech_inv i_15427(.A(n_63510), .Z(n_63595));
	notech_inv i_15426(.A(n_63593), .Z(n_63594));
	notech_inv i_15425(.A(n_63596), .Z(n_63593));
	notech_inv i_15424(.A(n_63591), .Z(n_63592));
	notech_inv i_15423(.A(n_63508), .Z(n_63591));
	notech_inv i_15422(.A(n_63589), .Z(n_63590));
	notech_inv i_15421(.A(n_63592), .Z(n_63589));
	notech_inv i_15420(.A(n_63587), .Z(n_63588));
	notech_inv i_15419(.A(n_63662), .Z(n_63587));
	notech_inv i_15418(.A(n_63585), .Z(n_63586));
	notech_inv i_15417(.A(n_63504), .Z(n_63585));
	notech_inv i_15416(.A(n_63583), .Z(n_63584));
	notech_inv i_15415(.A(n_63502), .Z(n_63583));
	notech_inv i_15414(.A(n_63581), .Z(n_63582));
	notech_inv i_15413(.A(n_63584), .Z(n_63581));
	notech_inv i_15412(.A(n_63579), .Z(n_63580));
	notech_inv i_15411(.A(n_63500), .Z(n_63579));
	notech_inv i_15410(.A(n_63577), .Z(n_63578));
	notech_inv i_15409(.A(n_63580), .Z(n_63577));
	notech_inv i_15408(.A(n_63575), .Z(n_63576));
	notech_inv i_15407(.A(n_63654), .Z(n_63575));
	notech_inv i_15406(.A(n_63573), .Z(n_63574));
	notech_inv i_15405(.A(n_63498), .Z(n_63573));
	notech_inv i_15404(.A(n_63571), .Z(n_63572));
	notech_inv i_15403(.A(n_63574), .Z(n_63571));
	notech_inv i_15402(.A(n_63569), .Z(n_63570));
	notech_inv i_15401(.A(n_63648), .Z(n_63569));
	notech_inv i_15400(.A(n_63567), .Z(n_63568));
	notech_inv i_15399(.A(n_63686), .Z(n_63567));
	notech_inv i_15398(.A(n_63565), .Z(n_63566));
	notech_inv i_15397(.A(n_63492), .Z(n_63565));
	notech_inv i_15378(.A(n_63545), .Z(n_63546));
	notech_inv i_15377(.A(n_63474), .Z(n_63545));
	notech_inv i_15376(.A(n_63543), .Z(n_63544));
	notech_inv i_15375(.A(n_63472), .Z(n_63543));
	notech_inv i_15374(.A(n_63541), .Z(n_63542));
	notech_inv i_15373(.A(n_63544), .Z(n_63541));
	notech_inv i_15372(.A(n_63539), .Z(n_63540));
	notech_inv i_15371(.A(n_63470), .Z(n_63539));
	notech_inv i_15370(.A(n_63537), .Z(n_63538));
	notech_inv i_15369(.A(n_63540), .Z(n_63537));
	notech_inv i_15368(.A(n_63535), .Z(n_63536));
	notech_inv i_15367(.A(n_63624), .Z(n_63535));
	notech_inv i_15366(.A(n_63533), .Z(n_63534));
	notech_inv i_15365(.A(n_63468), .Z(n_63533));
	notech_inv i_15364(.A(n_63531), .Z(n_63532));
	notech_inv i_15363(.A(n_63534), .Z(n_63531));
	notech_inv i_15362(.A(n_63529), .Z(n_63530));
	notech_inv i_15361(.A(n_63618), .Z(n_63529));
	notech_inv i_15360(.A(n_63527), .Z(n_63528));
	notech_inv i_15359(.A(n_63674), .Z(n_63527));
	notech_inv i_15358(.A(n_63525), .Z(n_63526));
	notech_inv i_15357(.A(n_63464), .Z(n_63525));
	notech_inv i_15356(.A(n_63523), .Z(n_63524));
	notech_inv i_15355(.A(n_63462), .Z(n_63523));
	notech_inv i_15354(.A(n_63521), .Z(n_63522));
	notech_inv i_15353(.A(n_63524), .Z(n_63521));
	notech_inv i_15352(.A(n_63519), .Z(n_63520));
	notech_inv i_15351(.A(n_63460), .Z(n_63519));
	notech_inv i_15350(.A(n_63517), .Z(n_63518));
	notech_inv i_15349(.A(n_63520), .Z(n_63517));
	notech_inv i_15348(.A(n_63515), .Z(n_63516));
	notech_inv i_15347(.A(n_63604), .Z(n_63515));
	notech_inv i_15346(.A(n_63513), .Z(n_63514));
	notech_inv i_15345(.A(n_63458), .Z(n_63513));
	notech_inv i_15344(.A(n_63511), .Z(n_63512));
	notech_inv i_15343(.A(n_63514), .Z(n_63511));
	notech_inv i_15342(.A(n_63509), .Z(n_63510));
	notech_inv i_15341(.A(n_63598), .Z(n_63509));
	notech_inv i_15340(.A(n_63507), .Z(n_63508));
	notech_inv i_15339(.A(n_63664), .Z(n_63507));
	notech_inv i_15338(.A(n_63505), .Z(n_63506));
	notech_inv i_15337(.A(n_63456), .Z(n_63505));
	notech_inv i_15336(.A(n_63503), .Z(n_63504));
	notech_inv i_15335(.A(n_63506), .Z(n_63503));
	notech_inv i_15334(.A(n_63501), .Z(n_63502));
	notech_inv i_15333(.A(n_63586), .Z(n_63501));
	notech_inv i_15332(.A(n_63499), .Z(n_63500));
	notech_inv i_15331(.A(n_63656), .Z(n_63499));
	notech_inv i_15330(.A(n_63497), .Z(n_63498));
	notech_inv i_15329(.A(n_63688), .Z(n_63497));
	notech_inv i_15328(.A(n_63495), .Z(n_63496));
	notech_inv i_15327(.A(n_63448), .Z(n_63495));
	notech_inv i_15326(.A(n_63493), .Z(n_63494));
	notech_inv i_15325(.A(n_63420), .Z(n_63493));
	notech_inv i_15324(.A(n_63491), .Z(n_63492));
	notech_inv i_15323(.A(n_63494), .Z(n_63491));
	notech_inv i_15308(.A(n_63475), .Z(n_63476));
	notech_inv i_15307(.A(n_63378), .Z(n_63475));
	notech_inv i_15306(.A(n_63473), .Z(n_63474));
	notech_inv i_15305(.A(n_63476), .Z(n_63473));
	notech_inv i_15304(.A(n_63471), .Z(n_63472));
	notech_inv i_15303(.A(n_63546), .Z(n_63471));
	notech_inv i_15302(.A(n_63469), .Z(n_63470));
	notech_inv i_15301(.A(n_63626), .Z(n_63469));
	notech_inv i_15300(.A(n_63467), .Z(n_63468));
	notech_inv i_15299(.A(n_63676), .Z(n_63467));
	notech_inv i_15298(.A(n_63465), .Z(n_63466));
	notech_inv i_15297(.A(n_63362), .Z(n_63465));
	notech_inv i_15296(.A(n_63463), .Z(n_63464));
	notech_inv i_15295(.A(n_63466), .Z(n_63463));
	notech_inv i_15294(.A(n_63461), .Z(n_63462));
	notech_inv i_15293(.A(n_63526), .Z(n_63461));
	notech_inv i_15292(.A(n_63459), .Z(n_63460));
	notech_inv i_15291(.A(n_63606), .Z(n_63459));
	notech_inv i_15290(.A(n_63457), .Z(n_63458));
	notech_inv i_15289(.A(n_63666), .Z(n_63457));
	notech_inv i_15288(.A(n_63455), .Z(n_63456));
	notech_inv i_15287(.A(n_63690), .Z(n_63455));
	notech_inv i_15280(.A(n_63447), .Z(n_63448));
	notech_inv i_15279(.A(clk), .Z(n_63447));
	notech_inv i_15252(.A(n_63419), .Z(n_63420));
	notech_inv i_15251(.A(n_63496), .Z(n_63419));
	notech_inv i_15210(.A(n_63377), .Z(n_63378));
	notech_inv i_15209(.A(n_63566), .Z(n_63377));
	notech_inv i_15194(.A(n_63361), .Z(n_63362));
	notech_inv i_15193(.A(n_63692), .Z(n_63361));
	notech_inv i_14336(.A(n_62348), .Z(n_62482));
	notech_inv i_14335(.A(n_62348), .Z(n_62481));
	notech_inv i_14334(.A(n_62348), .Z(n_62480));
	notech_inv i_14333(.A(n_62348), .Z(n_62479));
	notech_inv i_14331(.A(n_62348), .Z(n_62477));
	notech_inv i_14330(.A(n_62348), .Z(n_62476));
	notech_inv i_14329(.A(n_62348), .Z(n_62475));
	notech_inv i_14328(.A(n_62348), .Z(n_62474));
	notech_inv i_14325(.A(n_62348), .Z(n_62471));
	notech_inv i_14324(.A(n_62348), .Z(n_62470));
	notech_inv i_14323(.A(n_62348), .Z(n_62469));
	notech_inv i_14322(.A(n_62348), .Z(n_62468));
	notech_inv i_14320(.A(n_62348), .Z(n_62466));
	notech_inv i_14319(.A(n_62348), .Z(n_62465));
	notech_inv i_14318(.A(n_62348), .Z(n_62464));
	notech_inv i_14317(.A(n_62348), .Z(n_62463));
	notech_inv i_14314(.A(n_62451), .Z(n_62460));
	notech_inv i_14313(.A(n_62451), .Z(n_62459));
	notech_inv i_14312(.A(n_62451), .Z(n_62458));
	notech_inv i_14311(.A(n_62451), .Z(n_62457));
	notech_inv i_14309(.A(n_62451), .Z(n_62455));
	notech_inv i_14308(.A(n_62451), .Z(n_62454));
	notech_inv i_14307(.A(n_62451), .Z(n_62453));
	notech_inv i_14306(.A(n_62451), .Z(n_62452));
	notech_inv i_14305(.A(n_62468), .Z(n_62451));
	notech_inv i_14303(.A(n_62451), .Z(n_62449));
	notech_inv i_14302(.A(n_62451), .Z(n_62448));
	notech_inv i_14301(.A(n_62451), .Z(n_62447));
	notech_inv i_14300(.A(n_62451), .Z(n_62446));
	notech_inv i_14298(.A(n_62451), .Z(n_62444));
	notech_inv i_14297(.A(n_62451), .Z(n_62443));
	notech_inv i_14295(.A(n_62451), .Z(n_62441));
	notech_inv i_14291(.A(n_62428), .Z(n_62437));
	notech_inv i_14290(.A(n_62428), .Z(n_62436));
	notech_inv i_14288(.A(n_62428), .Z(n_62435));
	notech_inv i_14287(.A(n_62428), .Z(n_62434));
	notech_inv i_14285(.A(n_62428), .Z(n_62432));
	notech_inv i_14284(.A(n_62428), .Z(n_62431));
	notech_inv i_14283(.A(n_62428), .Z(n_62430));
	notech_inv i_14282(.A(n_62428), .Z(n_62429));
	notech_inv i_14280(.A(n_62474), .Z(n_62428));
	notech_inv i_14278(.A(n_62428), .Z(n_62426));
	notech_inv i_14277(.A(n_62428), .Z(n_62425));
	notech_inv i_14276(.A(n_62428), .Z(n_62424));
	notech_inv i_14275(.A(n_62428), .Z(n_62423));
	notech_inv i_14272(.A(n_62428), .Z(n_62421));
	notech_inv i_14271(.A(n_62428), .Z(n_62420));
	notech_inv i_14270(.A(n_62428), .Z(n_62419));
	notech_inv i_14269(.A(n_62428), .Z(n_62418));
	notech_inv i_14266(.A(n_62406), .Z(n_62415));
	notech_inv i_14264(.A(n_62406), .Z(n_62414));
	notech_inv i_14263(.A(n_62406), .Z(n_62413));
	notech_inv i_14262(.A(n_62406), .Z(n_62412));
	notech_inv i_14260(.A(n_62406), .Z(n_62410));
	notech_inv i_14259(.A(n_62406), .Z(n_62409));
	notech_inv i_14258(.A(n_62406), .Z(n_62408));
	notech_inv i_14256(.A(n_62406), .Z(n_62407));
	notech_inv i_14255(.A(n_62474), .Z(n_62406));
	notech_inv i_14253(.A(n_62406), .Z(n_62404));
	notech_inv i_14252(.A(n_62406), .Z(n_62403));
	notech_inv i_14251(.A(n_62406), .Z(n_62402));
	notech_inv i_14250(.A(n_62406), .Z(n_62401));
	notech_inv i_14247(.A(n_62406), .Z(n_62399));
	notech_inv i_14246(.A(n_62406), .Z(n_62398));
	notech_inv i_14245(.A(n_62406), .Z(n_62397));
	notech_inv i_14244(.A(n_62406), .Z(n_62396));
	notech_inv i_14239(.A(n_62383), .Z(n_62392));
	notech_inv i_14238(.A(n_62383), .Z(n_62391));
	notech_inv i_14237(.A(n_62383), .Z(n_62390));
	notech_inv i_14236(.A(n_62383), .Z(n_62389));
	notech_inv i_14234(.A(n_62383), .Z(n_62387));
	notech_inv i_14232(.A(n_62383), .Z(n_62386));
	notech_inv i_14231(.A(n_62383), .Z(n_62385));
	notech_inv i_14230(.A(n_62383), .Z(n_62384));
	notech_inv i_14229(.A(n_62468), .Z(n_62383));
	notech_inv i_14227(.A(n_62383), .Z(n_62381));
	notech_inv i_14226(.A(n_62383), .Z(n_62380));
	notech_inv i_14224(.A(n_62383), .Z(n_62379));
	notech_inv i_14223(.A(n_62383), .Z(n_62378));
	notech_inv i_14221(.A(n_62383), .Z(n_62376));
	notech_inv i_14220(.A(n_62383), .Z(n_62375));
	notech_inv i_14219(.A(n_62383), .Z(n_62374));
	notech_inv i_14218(.A(n_62383), .Z(n_62373));
	notech_inv i_14214(.A(n_62361), .Z(n_62370));
	notech_inv i_14213(.A(n_62361), .Z(n_62369));
	notech_inv i_14212(.A(n_62361), .Z(n_62368));
	notech_inv i_14211(.A(n_62361), .Z(n_62367));
	notech_inv i_14208(.A(n_62361), .Z(n_62365));
	notech_inv i_14207(.A(n_62361), .Z(n_62364));
	notech_inv i_14206(.A(n_62361), .Z(n_62363));
	notech_inv i_14205(.A(n_62361), .Z(n_62362));
	notech_inv i_14204(.A(n_62468), .Z(n_62361));
	notech_inv i_14202(.A(n_62361), .Z(n_62359));
	notech_inv i_14200(.A(n_62361), .Z(n_62358));
	notech_inv i_14199(.A(n_62361), .Z(n_62357));
	notech_inv i_14198(.A(n_62361), .Z(n_62356));
	notech_inv i_14196(.A(n_62361), .Z(n_62354));
	notech_inv i_14195(.A(n_62361), .Z(n_62353));
	notech_inv i_14194(.A(n_62361), .Z(n_62352));
	notech_inv i_14192(.A(n_62361), .Z(n_62351));
	notech_inv i_14189(.A(rstn), .Z(n_62348));
	notech_inv i_13820(.A(n_61963), .Z(n_61964));
	notech_inv i_13819(.A(instrc[121]), .Z(n_61963));
	notech_inv i_13815(.A(n_61952), .Z(n_61959));
	notech_inv i_13814(.A(n_61952), .Z(n_61958));
	notech_inv i_13808(.A(n_61952), .Z(n_61953));
	notech_inv i_13807(.A(n_2867), .Z(n_61952));
	notech_inv i_13799(.A(n_61943), .Z(n_61944));
	notech_inv i_13798(.A(instrc[122]), .Z(n_61943));
	notech_inv i_13796(.A(n_61922), .Z(n_61940));
	notech_inv i_13794(.A(n_61922), .Z(n_61938));
	notech_inv i_13790(.A(n_61922), .Z(n_61935));
	notech_inv i_13788(.A(n_61922), .Z(n_61933));
	notech_inv i_13784(.A(n_61922), .Z(n_61930));
	notech_inv i_13782(.A(n_61922), .Z(n_61928));
	notech_inv i_13778(.A(n_61922), .Z(n_61924));
	notech_inv i_13775(.A(n_1813), .Z(n_61922));
	notech_inv i_13771(.A(n_61906), .Z(n_61917));
	notech_inv i_13765(.A(n_61906), .Z(n_61912));
	notech_inv i_13759(.A(n_61906), .Z(n_61907));
	notech_inv i_13758(.A(fsm[1]), .Z(n_61906));
	notech_inv i_13756(.A(n_61895), .Z(n_61903));
	notech_inv i_13754(.A(n_61895), .Z(n_61901));
	notech_inv i_13750(.A(n_61895), .Z(n_61898));
	notech_inv i_13748(.A(n_61895), .Z(n_61896));
	notech_inv i_13747(.A(fsm[0]), .Z(n_61895));
	notech_inv i_13744(.A(n_61876), .Z(n_61892));
	notech_inv i_13742(.A(n_61876), .Z(n_61890));
	notech_inv i_13741(.A(n_61876), .Z(n_61889));
	notech_inv i_13736(.A(n_61876), .Z(n_61885));
	notech_inv i_13734(.A(n_61876), .Z(n_61883));
	notech_inv i_13731(.A(n_61876), .Z(n_61880));
	notech_inv i_13728(.A(n_61876), .Z(n_61878));
	notech_inv i_13727(.A(n_61876), .Z(n_61877));
	notech_inv i_13726(.A(n_316460792), .Z(n_61876));
	notech_inv i_13724(.A(n_61857), .Z(n_61873));
	notech_inv i_13722(.A(n_61857), .Z(n_61871));
	notech_inv i_13720(.A(n_61857), .Z(n_61870));
	notech_inv i_13716(.A(n_61857), .Z(n_61866));
	notech_inv i_13714(.A(n_61857), .Z(n_61864));
	notech_inv i_13710(.A(n_61857), .Z(n_61861));
	notech_inv i_13708(.A(n_61857), .Z(n_61859));
	notech_inv i_13707(.A(n_61857), .Z(n_61858));
	notech_inv i_13706(.A(pg_fault), .Z(n_61857));
	notech_inv i_13696(.A(n_61836), .Z(n_61846));
	notech_inv i_13695(.A(n_61836), .Z(n_61845));
	notech_inv i_13691(.A(n_61836), .Z(n_61841));
	notech_inv i_13687(.A(n_61836), .Z(n_61838));
	notech_inv i_13686(.A(n_61836), .Z(n_61837));
	notech_inv i_13685(.A(n_32789), .Z(n_61836));
	notech_inv i_13677(.A(n_61827), .Z(n_61828));
	notech_inv i_13676(.A(instrc[123]), .Z(n_61827));
	notech_inv i_13674(.A(n_61814), .Z(n_61824));
	notech_inv i_13672(.A(n_61814), .Z(n_61823));
	notech_inv i_13668(.A(n_61814), .Z(n_61819));
	notech_inv i_13663(.A(n_61814), .Z(n_61815));
	notech_inv i_13662(.A(n_32629), .Z(n_61814));
	notech_inv i_13654(.A(n_61805), .Z(n_61806));
	notech_inv i_13653(.A(n_2952), .Z(n_61805));
	notech_inv i_13645(.A(n_61796), .Z(n_61797));
	notech_inv i_13644(.A(n_32575), .Z(n_61796));
	notech_inv i_13634(.A(n_61785), .Z(n_61786));
	notech_inv i_13632(.A(instrc[120]), .Z(n_61785));
	notech_inv i_13622(.A(n_61774), .Z(n_61775));
	notech_inv i_13621(.A(n_32646), .Z(n_61774));
	notech_inv i_13613(.A(n_61765), .Z(n_61766));
	notech_inv i_13612(.A(n_32161), .Z(n_61765));
	notech_inv i_13604(.A(n_61756), .Z(n_61757));
	notech_inv i_13603(.A(n_32159), .Z(n_61756));
	notech_inv i_13595(.A(n_61747), .Z(n_61748));
	notech_inv i_13594(.A(n_309960727), .Z(n_61747));
	notech_inv i_13586(.A(n_61738), .Z(n_61739));
	notech_inv i_13584(.A(n_28008), .Z(n_61738));
	notech_inv i_13576(.A(n_61729), .Z(n_61730));
	notech_inv i_13575(.A(n_316260790), .Z(n_61729));
	notech_inv i_13572(.A(n_61730), .Z(n_61725));
	notech_inv i_13570(.A(n_61730), .Z(n_61723));
	notech_inv i_13564(.A(n_61730), .Z(n_61718));
	notech_inv i_13563(.A(n_61730), .Z(n_61717));
	notech_inv i_13556(.A(n_61730), .Z(n_61711));
	notech_inv i_13552(.A(n_61635), .Z(n_61707));
	notech_inv i_13551(.A(n_61635), .Z(n_61706));
	notech_inv i_13547(.A(n_61635), .Z(n_61702));
	notech_inv i_13542(.A(n_61635), .Z(n_61698));
	notech_inv i_13541(.A(n_61635), .Z(n_61697));
	notech_inv i_13536(.A(n_61635), .Z(n_61693));
	notech_inv i_13532(.A(n_61635), .Z(n_61689));
	notech_inv i_13531(.A(n_61635), .Z(n_61688));
	notech_inv i_13526(.A(n_61635), .Z(n_61684));
	notech_inv i_13522(.A(n_61635), .Z(n_61680));
	notech_inv i_13520(.A(n_61635), .Z(n_61679));
	notech_inv i_13516(.A(n_61635), .Z(n_61675));
	notech_inv i_13510(.A(n_61635), .Z(n_61670));
	notech_inv i_13509(.A(n_61635), .Z(n_61669));
	notech_inv i_13504(.A(n_61635), .Z(n_61665));
	notech_inv i_13500(.A(n_61635), .Z(n_61661));
	notech_inv i_13499(.A(n_61635), .Z(n_61660));
	notech_inv i_13494(.A(n_61635), .Z(n_61656));
	notech_inv i_13490(.A(n_61646), .Z(n_61652));
	notech_inv i_13488(.A(n_61646), .Z(n_61651));
	notech_inv i_13484(.A(n_61646), .Z(n_61647));
	notech_inv i_13483(.A(n_61660), .Z(n_61646));
	notech_inv i_13479(.A(n_61635), .Z(n_61643));
	notech_inv i_13478(.A(n_61635), .Z(n_61642));
	notech_inv i_13470(.A(n_1974696898), .Z(n_61635));
	notech_inv i_13468(.A(n_61606), .Z(n_61632));
	notech_inv i_13466(.A(n_61606), .Z(n_61630));
	notech_inv i_13463(.A(n_61606), .Z(n_61628));
	notech_inv i_13460(.A(n_61606), .Z(n_61625));
	notech_inv i_13458(.A(n_61606), .Z(n_61623));
	notech_inv i_13455(.A(n_61606), .Z(n_61621));
	notech_inv i_13452(.A(n_61606), .Z(n_61618));
	notech_inv i_13450(.A(n_61606), .Z(n_61616));
	notech_inv i_13447(.A(n_61606), .Z(n_61614));
	notech_inv i_13444(.A(n_61606), .Z(n_61611));
	notech_inv i_13442(.A(n_61606), .Z(n_61609));
	notech_inv i_13439(.A(n_61606), .Z(n_61607));
	notech_inv i_13438(.A(n_31365), .Z(n_61606));
	notech_inv i_13428(.A(n_61595), .Z(n_61596));
	notech_inv i_13427(.A(n_97990346), .Z(n_61595));
	notech_inv i_13386(.A(n_61446), .Z(n_61456));
	notech_inv i_13384(.A(n_61446), .Z(n_61455));
	notech_inv i_13380(.A(n_61446), .Z(n_61451));
	notech_inv i_13375(.A(n_61446), .Z(n_61447));
	notech_inv i_13374(.A(ipg_fault), .Z(n_61446));
	notech_inv i_13222(.A(n_61273), .Z(n_61286));
	notech_inv i_13220(.A(n_61273), .Z(n_61284));
	notech_inv i_13216(.A(n_61273), .Z(n_61281));
	notech_inv i_13214(.A(n_61273), .Z(n_61279));
	notech_inv i_13210(.A(n_61273), .Z(n_61275));
	notech_inv i_13208(.A(n_61273), .Z(cr0[0]));
	notech_inv i_13207(.A(\nbus_14546[0] ), .Z(n_61273));
	notech_inv i_13066(.A(n_61118), .Z(n_61119));
	notech_inv i_13065(.A(n_19698), .Z(n_61118));
	notech_inv i_13058(.A(n_61109), .Z(n_61110));
	notech_inv i_13057(.A(n_30712), .Z(n_61109));
	notech_inv i_13055(.A(n_61084), .Z(n_61106));
	notech_inv i_13053(.A(n_61084), .Z(n_61104));
	notech_inv i_13052(.A(n_61084), .Z(n_61103));
	notech_inv i_13048(.A(n_61084), .Z(n_61099));
	notech_inv i_13046(.A(n_61084), .Z(n_61097));
	notech_inv i_13043(.A(n_61084), .Z(n_61094));
	notech_inv i_13041(.A(n_61084), .Z(n_61092));
	notech_inv i_13040(.A(n_61084), .Z(n_61091));
	notech_inv i_13036(.A(n_61084), .Z(n_61087));
	notech_inv i_13034(.A(n_61084), .Z(n_61085));
	notech_inv i_13033(.A(n_33158), .Z(n_61084));
	notech_inv i_13026(.A(n_61075), .Z(n_61076));
	notech_inv i_13025(.A(n_314960777), .Z(n_61075));
	notech_inv i_13016(.A(n_61064), .Z(n_61065));
	notech_inv i_13015(.A(n_28098), .Z(n_61064));
	notech_inv i_13008(.A(n_61051), .Z(n_61056));
	notech_inv i_13004(.A(n_61051), .Z(n_61052));
	notech_inv i_13003(.A(n_32397), .Z(n_61051));
	notech_inv i_12996(.A(n_61042), .Z(n_61043));
	notech_inv i_12995(.A(n_113490501), .Z(n_61042));
	notech_inv i_12988(.A(n_61033), .Z(n_61034));
	notech_inv i_12987(.A(opa[15]), .Z(n_61033));
	notech_inv i_12980(.A(n_61024), .Z(n_61025));
	notech_inv i_12979(.A(opa[13]), .Z(n_61024));
	notech_inv i_12972(.A(n_61015), .Z(n_61016));
	notech_inv i_12971(.A(opa[12]), .Z(n_61015));
	notech_inv i_12964(.A(n_61006), .Z(n_61007));
	notech_inv i_12963(.A(opa[9]), .Z(n_61006));
	notech_inv i_12956(.A(n_60997), .Z(n_60998));
	notech_inv i_12955(.A(opa[7]), .Z(n_60997));
	notech_inv i_12948(.A(n_60988), .Z(n_60989));
	notech_inv i_12947(.A(opa[6]), .Z(n_60988));
	notech_inv i_12939(.A(n_60979), .Z(n_60980));
	notech_inv i_12938(.A(opa[5]), .Z(n_60979));
	notech_inv i_12930(.A(n_60970), .Z(n_60971));
	notech_inv i_12928(.A(opa[3]), .Z(n_60970));
	notech_inv i_12920(.A(n_60961), .Z(n_60962));
	notech_inv i_12919(.A(opa[2]), .Z(n_60961));
	notech_inv i_12911(.A(n_60952), .Z(n_60953));
	notech_inv i_12910(.A(opa[0]), .Z(n_60952));
	notech_inv i_12604(.A(n_60628), .Z(n_60629));
	notech_inv i_12603(.A(opb[31]), .Z(n_60628));
	notech_inv i_12595(.A(n_60619), .Z(n_60620));
	notech_inv i_12594(.A(nbus_11271[29]), .Z(n_60619));
	notech_inv i_12586(.A(n_60610), .Z(n_60611));
	notech_inv i_12585(.A(nbus_11271[30]), .Z(n_60610));
	notech_inv i_12582(.A(n_60599), .Z(n_60607));
	notech_inv i_12580(.A(n_60599), .Z(n_60605));
	notech_inv i_12577(.A(n_60599), .Z(n_60602));
	notech_inv i_12574(.A(n_60599), .Z(n_60600));
	notech_inv i_12573(.A(opc[31]), .Z(n_60599));
	notech_inv i_12565(.A(n_60590), .Z(n_60591));
	notech_inv i_12564(.A(nbus_11271[31]), .Z(n_60590));
	notech_inv i_12556(.A(n_60581), .Z(n_60582));
	notech_inv i_12555(.A(nbus_11271[26]), .Z(n_60581));
	notech_inv i_12547(.A(n_60572), .Z(n_60573));
	notech_inv i_12546(.A(nbus_11271[27]), .Z(n_60572));
	notech_inv i_12538(.A(n_60563), .Z(n_60564));
	notech_inv i_12537(.A(nbus_11271[28]), .Z(n_60563));
	notech_inv i_12529(.A(n_60554), .Z(n_60555));
	notech_inv i_12527(.A(nbus_11271[20]), .Z(n_60554));
	notech_inv i_12519(.A(n_60545), .Z(n_60546));
	notech_inv i_12518(.A(nbus_11271[21]), .Z(n_60545));
	notech_inv i_12510(.A(n_60536), .Z(n_60537));
	notech_inv i_12508(.A(nbus_11271[22]), .Z(n_60536));
	notech_inv i_12499(.A(n_60527), .Z(n_60528));
	notech_inv i_12498(.A(nbus_11271[23]), .Z(n_60527));
	notech_inv i_12490(.A(n_60518), .Z(n_60519));
	notech_inv i_12489(.A(nbus_11271[24]), .Z(n_60518));
	notech_inv i_12481(.A(n_60509), .Z(n_60510));
	notech_inv i_12480(.A(nbus_11271[25]), .Z(n_60509));
	notech_inv i_12472(.A(n_60500), .Z(n_60501));
	notech_inv i_12471(.A(nbus_11271[17]), .Z(n_60500));
	notech_inv i_12463(.A(n_60491), .Z(n_60492));
	notech_inv i_12461(.A(nbus_11271[18]), .Z(n_60491));
	notech_inv i_12453(.A(n_60482), .Z(n_60483));
	notech_inv i_12452(.A(nbus_11271[19]), .Z(n_60482));
	notech_inv i_12444(.A(n_60473), .Z(n_60474));
	notech_inv i_12443(.A(nbus_11271[16]), .Z(n_60473));
	notech_inv i_12437(.A(n_60466), .Z(n_60467));
	notech_inv i_12436(.A(opc[0]), .Z(n_60466));
	notech_inv i_12428(.A(n_60457), .Z(n_60458));
	notech_inv i_12427(.A(\nbus_11283[31] ), .Z(n_60457));
	notech_inv i_12425(.A(n_60448), .Z(n_60454));
	notech_inv i_12424(.A(n_60448), .Z(n_60453));
	notech_inv i_12419(.A(n_60448), .Z(n_60449));
	notech_inv i_12418(.A(n_32195), .Z(n_60448));
	notech_inv i_12410(.A(n_60439), .Z(n_60440));
	notech_inv i_12409(.A(instrc[113]), .Z(n_60439));
	notech_inv i_12401(.A(n_60430), .Z(n_60431));
	notech_inv i_12400(.A(instrc[114]), .Z(n_60430));
	notech_inv i_12392(.A(n_60421), .Z(n_60422));
	notech_inv i_12391(.A(instrc[112]), .Z(n_60421));
	notech_inv i_12168(.A(n_32583), .Z(n_60196));
	notech_inv i_12165(.A(n_32583), .Z(n_60194));
	notech_inv i_12160(.A(n_32583), .Z(n_60189));
	notech_inv i_12158(.A(n_32583), .Z(n_60188));
	notech_inv i_12152(.A(n_32583), .Z(n_60182));
	notech_inv i_12147(.A(n_60162), .Z(n_60177));
	notech_inv i_12145(.A(n_60162), .Z(n_60175));
	notech_inv i_12139(.A(n_60162), .Z(n_60170));
	notech_inv i_12138(.A(n_60162), .Z(n_60169));
	notech_inv i_12131(.A(n_60162), .Z(n_60163));
	notech_inv i_12130(.A(n_32401), .Z(n_60162));
	notech_inv i_12128(.A(n_32697), .Z(n_60159));
	notech_inv i_12125(.A(n_32697), .Z(n_60157));
	notech_inv i_12122(.A(n_32697), .Z(n_60154));
	notech_inv i_12120(.A(n_32697), .Z(n_60152));
	notech_inv i_11150(.A(n_59119), .Z(n_59120));
	notech_inv i_11149(.A(n_28534), .Z(n_59119));
	notech_inv i_11144(.A(n_59103), .Z(n_59115));
	notech_inv i_11143(.A(n_59103), .Z(n_59114));
	notech_inv i_11137(.A(n_59103), .Z(n_59109));
	notech_inv i_11132(.A(n_59103), .Z(n_59104));
	notech_inv i_11130(.A(n_2094), .Z(n_59103));
	notech_inv i_11128(.A(n_32548), .Z(n_59100));
	notech_inv i_11127(.A(n_32548), .Z(n_59099));
	notech_inv i_11122(.A(n_32548), .Z(n_59095));
	notech_inv i_11113(.A(n_59085), .Z(n_59086));
	notech_inv i_11112(.A(\nbus_11290[17] ), .Z(n_59085));
	notech_inv i_11104(.A(n_59076), .Z(n_59077));
	notech_inv i_11103(.A(\nbus_11290[18] ), .Z(n_59076));
	notech_inv i_11095(.A(n_59067), .Z(n_59068));
	notech_inv i_11094(.A(\nbus_11290[15] ), .Z(n_59067));
	notech_inv i_11086(.A(n_59058), .Z(n_59059));
	notech_inv i_11085(.A(\nbus_11290[16] ), .Z(n_59058));
	notech_inv i_11077(.A(n_59049), .Z(n_59050));
	notech_inv i_11076(.A(\nbus_11290[12] ), .Z(n_59049));
	notech_inv i_11068(.A(n_59040), .Z(n_59041));
	notech_inv i_11066(.A(\nbus_11290[14] ), .Z(n_59040));
	notech_inv i_11058(.A(n_59031), .Z(n_59032));
	notech_inv i_11057(.A(\nbus_11290[9] ), .Z(n_59031));
	notech_inv i_11049(.A(n_59022), .Z(n_59023));
	notech_inv i_11048(.A(\nbus_11290[10] ), .Z(n_59022));
	notech_inv i_11040(.A(n_59013), .Z(n_59014));
	notech_inv i_11039(.A(\nbus_11290[8] ), .Z(n_59013));
	notech_inv i_11031(.A(n_59000), .Z(n_59005));
	notech_inv i_11026(.A(n_59000), .Z(n_59001));
	notech_inv i_11025(.A(\nbus_11290[1] ), .Z(n_59000));
	notech_inv i_11017(.A(n_58991), .Z(n_58992));
	notech_inv i_11016(.A(\nbus_11290[30] ), .Z(n_58991));
	notech_inv i_11008(.A(n_58982), .Z(n_58983));
	notech_inv i_11007(.A(\nbus_11290[31] ), .Z(n_58982));
	notech_inv i_10999(.A(n_58973), .Z(n_58974));
	notech_inv i_10998(.A(\nbus_11290[11] ), .Z(n_58973));
	notech_inv i_10990(.A(n_58964), .Z(n_58965));
	notech_inv i_10989(.A(\nbus_11290[13] ), .Z(n_58964));
	notech_inv i_10981(.A(n_58955), .Z(n_58956));
	notech_inv i_10980(.A(\nbus_11290[0] ), .Z(n_58955));
	notech_inv i_10972(.A(n_58946), .Z(n_58947));
	notech_inv i_10970(.A(\nbus_11290[29] ), .Z(n_58946));
	notech_inv i_10962(.A(n_58937), .Z(n_58938));
	notech_inv i_10961(.A(\nbus_11290[27] ), .Z(n_58937));
	notech_inv i_10953(.A(n_58928), .Z(n_58929));
	notech_inv i_10952(.A(\nbus_11290[28] ), .Z(n_58928));
	notech_inv i_10944(.A(n_58919), .Z(n_58920));
	notech_inv i_10943(.A(\nbus_11290[25] ), .Z(n_58919));
	notech_inv i_10935(.A(n_58910), .Z(n_58911));
	notech_inv i_10934(.A(\nbus_11290[26] ), .Z(n_58910));
	notech_inv i_10926(.A(n_58901), .Z(n_58902));
	notech_inv i_10925(.A(\nbus_11290[23] ), .Z(n_58901));
	notech_inv i_10917(.A(n_58892), .Z(n_58893));
	notech_inv i_10916(.A(\nbus_11290[24] ), .Z(n_58892));
	notech_inv i_10908(.A(n_58883), .Z(n_58884));
	notech_inv i_10906(.A(\nbus_11290[21] ), .Z(n_58883));
	notech_inv i_10898(.A(n_58874), .Z(n_58875));
	notech_inv i_10897(.A(\nbus_11290[22] ), .Z(n_58874));
	notech_inv i_10889(.A(n_58865), .Z(n_58866));
	notech_inv i_10888(.A(\nbus_11290[19] ), .Z(n_58865));
	notech_inv i_10880(.A(n_58856), .Z(n_58857));
	notech_inv i_10879(.A(\nbus_11290[20] ), .Z(n_58856));
	notech_inv i_10871(.A(n_58847), .Z(n_58848));
	notech_inv i_10870(.A(n_391464445), .Z(n_58847));
	notech_inv i_10862(.A(n_58838), .Z(n_58839));
	notech_inv i_10861(.A(n_30367), .Z(n_58838));
	notech_inv i_10858(.A(n_58819), .Z(n_58835));
	notech_inv i_10856(.A(n_58819), .Z(n_58833));
	notech_inv i_10855(.A(n_58819), .Z(n_58832));
	notech_inv i_10849(.A(n_58819), .Z(n_58827));
	notech_inv i_10841(.A(n_58819), .Z(n_58820));
	notech_inv i_10840(.A(n_57675), .Z(n_58819));
	notech_inv i_10823(.A(n_58801), .Z(n_58802));
	notech_inv i_10822(.A(n_31474), .Z(n_58801));
	notech_inv i_10805(.A(n_58783), .Z(n_58784));
	notech_inv i_10804(.A(n_31476), .Z(n_58783));
	notech_inv i_10736(.A(n_58715), .Z(n_58716));
	notech_inv i_10735(.A(n_340461032), .Z(n_58715));
	notech_inv i_10727(.A(n_58706), .Z(n_58707));
	notech_inv i_10726(.A(n_2830), .Z(n_58706));
	notech_inv i_10722(.A(n_32342), .Z(n_58702));
	notech_inv i_10721(.A(n_32342), .Z(n_58701));
	notech_inv i_10716(.A(n_32342), .Z(n_58696));
	notech_inv i_10708(.A(n_32342), .Z(n_58691));
	notech_inv i_10699(.A(n_58681), .Z(n_58682));
	notech_inv i_10698(.A(n_336689251), .Z(n_58681));
	notech_inv i_10690(.A(n_58672), .Z(n_58673));
	notech_inv i_10688(.A(n_390164432), .Z(n_58672));
	notech_inv i_10680(.A(n_58663), .Z(n_58664));
	notech_inv i_10679(.A(n_25094), .Z(n_58663));
	notech_inv i_10671(.A(n_58654), .Z(n_58655));
	notech_inv i_10670(.A(n_4460), .Z(n_58654));
	notech_inv i_10662(.A(n_58645), .Z(n_58646));
	notech_inv i_10661(.A(n_1840), .Z(n_58645));
	notech_inv i_10653(.A(n_58636), .Z(n_58637));
	notech_inv i_10652(.A(n_4461), .Z(n_58636));
	notech_inv i_10644(.A(n_58627), .Z(n_58628));
	notech_inv i_10643(.A(n_30680), .Z(n_58627));
	notech_inv i_10635(.A(n_58618), .Z(n_58619));
	notech_inv i_10634(.A(n_348989371), .Z(n_58618));
	notech_inv i_10626(.A(n_58609), .Z(n_58610));
	notech_inv i_10624(.A(n_340561033), .Z(n_58609));
	notech_inv i_10616(.A(n_58600), .Z(n_58601));
	notech_inv i_10615(.A(n_32268), .Z(n_58600));
	notech_inv i_10613(.A(n_58601), .Z(n_58597));
	notech_inv i_10612(.A(n_58601), .Z(n_58596));
	notech_inv i_10607(.A(n_58601), .Z(n_58592));
	notech_inv i_10598(.A(n_58582), .Z(n_58583));
	notech_inv i_10597(.A(n_32275), .Z(n_58582));
	notech_inv i_10589(.A(n_58569), .Z(n_58574));
	notech_inv i_10584(.A(n_58569), .Z(n_58570));
	notech_inv i_10583(.A(n_30664), .Z(n_58569));
	notech_inv i_10581(.A(n_32249), .Z(n_58566));
	notech_inv i_10580(.A(n_32249), .Z(n_58565));
	notech_inv i_10575(.A(n_32249), .Z(n_58561));
	notech_inv i_10570(.A(n_32263), .Z(n_58555));
	notech_inv i_10564(.A(n_32263), .Z(n_58550));
	notech_inv i_10555(.A(n_58540), .Z(n_58541));
	notech_inv i_10554(.A(n_25467), .Z(n_58540));
	notech_inv i_10546(.A(n_58531), .Z(n_58532));
	notech_inv i_10544(.A(n_27843), .Z(n_58531));
	notech_inv i_10536(.A(n_58522), .Z(n_58523));
	notech_inv i_10535(.A(n_27919), .Z(n_58522));
	notech_inv i_10525(.A(n_58511), .Z(n_58512));
	notech_inv i_10524(.A(n_23345), .Z(n_58511));
	notech_inv i_10519(.A(n_58500), .Z(n_58506));
	notech_inv i_10514(.A(n_58500), .Z(n_58501));
	notech_inv i_10512(.A(n_318660814), .Z(n_58500));
	notech_inv i_10504(.A(n_58491), .Z(n_58492));
	notech_inv i_10503(.A(n_23353), .Z(n_58491));
	notech_inv i_10495(.A(n_58482), .Z(n_58483));
	notech_inv i_10494(.A(\nbus_11283[30] ), .Z(n_58482));
	notech_inv i_10486(.A(n_58473), .Z(n_58474));
	notech_inv i_10485(.A(\nbus_11283[29] ), .Z(n_58473));
	notech_inv i_10477(.A(n_58464), .Z(n_58465));
	notech_inv i_10476(.A(\nbus_11283[28] ), .Z(n_58464));
	notech_inv i_10468(.A(n_58455), .Z(n_58456));
	notech_inv i_10467(.A(\nbus_11283[27] ), .Z(n_58455));
	notech_inv i_10459(.A(n_58446), .Z(n_58447));
	notech_inv i_10458(.A(\nbus_11283[26] ), .Z(n_58446));
	notech_inv i_10450(.A(n_58437), .Z(n_58438));
	notech_inv i_10448(.A(\nbus_11283[25] ), .Z(n_58437));
	notech_inv i_10440(.A(n_58428), .Z(n_58429));
	notech_inv i_10439(.A(\nbus_11283[24] ), .Z(n_58428));
	notech_inv i_10431(.A(n_58419), .Z(n_58420));
	notech_inv i_10430(.A(\nbus_11283[23] ), .Z(n_58419));
	notech_inv i_10422(.A(n_58410), .Z(n_58411));
	notech_inv i_10421(.A(\nbus_11283[22] ), .Z(n_58410));
	notech_inv i_10413(.A(n_58401), .Z(n_58402));
	notech_inv i_10412(.A(\nbus_11283[21] ), .Z(n_58401));
	notech_inv i_10404(.A(n_58392), .Z(n_58393));
	notech_inv i_10403(.A(\nbus_11283[20] ), .Z(n_58392));
	notech_inv i_10395(.A(n_58383), .Z(n_58384));
	notech_inv i_10394(.A(\nbus_11283[19] ), .Z(n_58383));
	notech_inv i_10386(.A(n_58374), .Z(n_58375));
	notech_inv i_10385(.A(\nbus_11283[18] ), .Z(n_58374));
	notech_inv i_10377(.A(n_58365), .Z(n_58366));
	notech_inv i_10375(.A(\nbus_11283[17] ), .Z(n_58365));
	notech_inv i_10367(.A(n_58356), .Z(n_58357));
	notech_inv i_10366(.A(\nbus_11283[16] ), .Z(n_58356));
	notech_inv i_10358(.A(n_58347), .Z(n_58348));
	notech_inv i_10357(.A(nbus_11273[15]), .Z(n_58347));
	notech_inv i_10349(.A(n_58338), .Z(n_58339));
	notech_inv i_10348(.A(nbus_11273[14]), .Z(n_58338));
	notech_inv i_10340(.A(n_58329), .Z(n_58330));
	notech_inv i_10339(.A(nbus_11273[13]), .Z(n_58329));
	notech_inv i_10331(.A(n_58320), .Z(n_58321));
	notech_inv i_10330(.A(nbus_11273[12]), .Z(n_58320));
	notech_inv i_10322(.A(n_58311), .Z(n_58312));
	notech_inv i_10321(.A(nbus_11273[11]), .Z(n_58311));
	notech_inv i_10313(.A(n_58302), .Z(n_58303));
	notech_inv i_10310(.A(nbus_11273[10]), .Z(n_58302));
	notech_inv i_10302(.A(n_58293), .Z(n_58294));
	notech_inv i_10301(.A(nbus_11273[9]), .Z(n_58293));
	notech_inv i_10293(.A(n_58284), .Z(n_58285));
	notech_inv i_10292(.A(nbus_11273[8]), .Z(n_58284));
	notech_inv i_10281(.A(n_58273), .Z(n_58275));
	notech_inv i_10280(.A(nbus_11273[7]), .Z(n_58273));
	notech_inv i_10270(.A(n_58264), .Z(n_58265));
	notech_inv i_10269(.A(nbus_11273[6]), .Z(n_58264));
	notech_inv i_10261(.A(n_58255), .Z(n_58256));
	notech_inv i_10260(.A(nbus_11273[3]), .Z(n_58255));
	notech_inv i_10252(.A(n_58246), .Z(n_58247));
	notech_inv i_10251(.A(nbus_11273[2]), .Z(n_58246));
	notech_inv i_10243(.A(n_58237), .Z(n_58238));
	notech_inv i_10241(.A(nbus_11273[0]), .Z(n_58237));
	notech_inv i_10233(.A(n_58224), .Z(n_58229));
	notech_inv i_10229(.A(n_58224), .Z(n_58225));
	notech_inv i_10228(.A(nbus_11273[1]), .Z(n_58224));
	notech_inv i_10220(.A(n_58214), .Z(n_58215));
	notech_inv i_10219(.A(n_27814), .Z(n_58214));
	notech_inv i_10212(.A(n_33164), .Z(n_58206));
	notech_inv i_10211(.A(n_33164), .Z(n_58205));
	notech_inv i_10207(.A(n_33164), .Z(n_58202));
	notech_inv i_10206(.A(n_33164), .Z(n_58201));
	notech_inv i_10159(.A(n_58017), .Z(n_58018));
	notech_inv i_10158(.A(opd[31]), .Z(n_58017));
	notech_inv i_10148(.A(n_58006), .Z(n_58007));
	notech_inv i_10147(.A(n_23334), .Z(n_58006));
	notech_inv i_10139(.A(n_57997), .Z(n_57998));
	notech_inv i_10137(.A(n_23379), .Z(n_57997));
	notech_inv i_10127(.A(n_57986), .Z(n_57987));
	notech_inv i_10126(.A(n_30612), .Z(n_57986));
	notech_inv i_10118(.A(n_57973), .Z(n_57978));
	notech_inv i_10113(.A(n_57973), .Z(n_57974));
	notech_inv i_10112(.A(n_218373551), .Z(n_57973));
	notech_inv i_10104(.A(n_57964), .Z(n_57965));
	notech_inv i_10103(.A(opd[26]), .Z(n_57964));
	notech_inv i_10095(.A(n_57955), .Z(n_57956));
	notech_inv i_10094(.A(opd[27]), .Z(n_57955));
	notech_inv i_10086(.A(n_57945), .Z(n_57946));
	notech_inv i_10085(.A(opd[28]), .Z(n_57945));
	notech_inv i_10077(.A(n_57936), .Z(n_57937));
	notech_inv i_10076(.A(opd[29]), .Z(n_57936));
	notech_inv i_10067(.A(n_57927), .Z(n_57928));
	notech_inv i_10066(.A(n_301874370), .Z(n_57927));
	notech_inv i_10055(.A(n_57916), .Z(n_57917));
	notech_inv i_10054(.A(n_23373), .Z(n_57916));
	notech_inv i_10046(.A(n_57906), .Z(n_57907));
	notech_inv i_10045(.A(n_23371), .Z(n_57906));
	notech_inv i_10035(.A(n_57895), .Z(n_57896));
	notech_inv i_10034(.A(n_23367), .Z(n_57895));
	notech_inv i_10026(.A(n_57886), .Z(n_57887));
	notech_inv i_10024(.A(n_1826), .Z(n_57886));
	notech_inv i_10016(.A(n_57877), .Z(n_57878));
	notech_inv i_10015(.A(n_317751253), .Z(n_57877));
	notech_inv i_10005(.A(n_57866), .Z(n_57867));
	notech_inv i_10004(.A(n_1828), .Z(n_57866));
	notech_inv i_9894(.A(n_57744), .Z(n_57745));
	notech_inv i_9893(.A(n_1827), .Z(n_57744));
	notech_inv i_9867(.A(n_57713), .Z(n_57714));
	notech_inv i_9866(.A(instrc[119]), .Z(n_57713));
	notech_inv i_9858(.A(n_57704), .Z(n_57705));
	notech_inv i_9856(.A(instrc[118]), .Z(n_57704));
	notech_inv i_9848(.A(n_57695), .Z(n_57696));
	notech_inv i_9847(.A(instrc[117]), .Z(n_57695));
	notech_inv i_9839(.A(n_57685), .Z(n_57686));
	notech_inv i_9838(.A(n_33173), .Z(n_57685));
	notech_inv i_9834(.A(n_57671), .Z(n_57679));
	notech_inv i_9828(.A(n_57671), .Z(n_57672));
	notech_inv i_9827(.A(n_32319), .Z(n_57671));
	notech_inv i_9819(.A(n_57661), .Z(n_57662));
	notech_inv i_9818(.A(n_30698), .Z(n_57661));
	notech_inv i_9814(.A(n_57650), .Z(n_57657));
	notech_inv i_9813(.A(n_57650), .Z(n_57656));
	notech_inv i_9806(.A(n_57650), .Z(n_57651));
	notech_inv i_9805(.A(n_30678), .Z(n_57650));
	notech_inv i_9797(.A(n_57641), .Z(n_57642));
	notech_inv i_9796(.A(n_30737), .Z(n_57641));
	notech_inv i_9794(.A(n_32317), .Z(n_57638));
	notech_inv i_9793(.A(n_32317), .Z(n_57637));
	notech_inv i_9788(.A(n_32317), .Z(n_57633));
	notech_inv i_9782(.A(n_32252), .Z(n_57627));
	notech_inv i_9777(.A(n_32252), .Z(n_57622));
	notech_inv i_9771(.A(n_32227), .Z(n_57616));
	notech_inv i_9764(.A(n_32227), .Z(n_57609));
	notech_inv i_9757(.A(n_32227), .Z(n_57604));
	notech_inv i_9748(.A(n_57594), .Z(n_57595));
	notech_inv i_9747(.A(n_321860846), .Z(n_57594));
	notech_inv i_9739(.A(n_57585), .Z(n_57586));
	notech_inv i_9738(.A(n_30739), .Z(n_57585));
	notech_inv i_9728(.A(n_57574), .Z(n_57575));
	notech_inv i_9727(.A(n_157062602), .Z(n_57574));
	notech_inv i_9719(.A(n_57561), .Z(n_57566));
	notech_inv i_9714(.A(n_57561), .Z(n_57562));
	notech_inv i_9713(.A(n_32314), .Z(n_57561));
	notech_inv i_9705(.A(n_57552), .Z(n_57553));
	notech_inv i_9704(.A(n_30719), .Z(n_57552));
	notech_inv i_9696(.A(n_57543), .Z(n_57544));
	notech_inv i_9695(.A(n_116742608), .Z(n_57543));
	notech_inv i_9687(.A(n_57534), .Z(n_57535));
	notech_inv i_9685(.A(n_30309), .Z(n_57534));
	notech_inv i_9681(.A(n_32254), .Z(n_57529));
	notech_inv i_9675(.A(n_32254), .Z(n_57524));
	notech_inv i_9669(.A(n_32266), .Z(n_57517));
	notech_inv i_9664(.A(n_32266), .Z(n_57512));
	notech_inv i_9658(.A(n_32261), .Z(n_57506));
	notech_inv i_9652(.A(n_32261), .Z(n_57500));
	notech_inv i_9647(.A(n_32259), .Z(n_57494));
	notech_inv i_9641(.A(n_32259), .Z(n_57489));
	notech_inv i_9632(.A(n_57475), .Z(n_57480));
	notech_inv i_9627(.A(n_57475), .Z(n_57476));
	notech_inv i_9626(.A(n_30363), .Z(n_57475));
	notech_inv i_9624(.A(n_32244), .Z(n_57472));
	notech_inv i_9623(.A(n_32244), .Z(n_57471));
	notech_inv i_9618(.A(n_32244), .Z(n_57467));
	notech_inv i_9612(.A(n_32243), .Z(n_57461));
	notech_inv i_9607(.A(n_32243), .Z(n_57456));
	notech_inv i_9601(.A(n_32304), .Z(n_57449));
	notech_inv i_9595(.A(n_32304), .Z(n_57444));
	notech_inv i_9591(.A(n_32273), .Z(n_57436));
	notech_inv i_9589(.A(n_32273), .Z(n_57435));
	notech_inv i_9584(.A(n_32273), .Z(n_57429));
	notech_inv i_9578(.A(n_32273), .Z(n_57423));
	notech_inv i_9572(.A(n_32544), .Z(n_57417));
	notech_inv i_9567(.A(n_32544), .Z(n_57412));
	notech_inv i_9562(.A(n_32272), .Z(n_57407));
	notech_inv i_9561(.A(n_32272), .Z(n_57406));
	notech_inv i_9555(.A(n_32272), .Z(n_57401));
	notech_inv i_9552(.A(n_57375), .Z(n_57397));
	notech_inv i_9549(.A(n_57375), .Z(n_57395));
	notech_inv i_9548(.A(n_57375), .Z(n_57392));
	notech_inv i_9544(.A(n_57375), .Z(n_57386));
	notech_inv i_9541(.A(n_57375), .Z(n_57382));
	notech_inv i_9537(.A(n_57375), .Z(n_57378));
	notech_inv i_9533(.A(n_30729), .Z(n_57375));
	notech_inv i_9424(.A(n_57250), .Z(n_57256));
	notech_inv i_9419(.A(n_57250), .Z(n_57251));
	notech_inv i_9418(.A(n_444168025), .Z(n_57250));
	notech_inv i_9406(.A(n_57235), .Z(n_57236));
	notech_inv i_9405(.A(n_32203), .Z(n_57235));
	notech_inv i_9400(.A(n_57236), .Z(n_57230));
	notech_inv i_9394(.A(n_57236), .Z(n_57225));
	notech_inv i_9388(.A(n_32204), .Z(n_57218));
	notech_inv i_9382(.A(n_32204), .Z(n_57211));
	notech_inv i_9373(.A(n_57198), .Z(n_57199));
	notech_inv i_9372(.A(n_30679), .Z(n_57198));
	notech_inv i_9370(.A(n_32216), .Z(n_57195));
	notech_inv i_9367(.A(n_32216), .Z(n_57192));
	notech_inv i_9364(.A(n_32216), .Z(n_57189));
	notech_inv i_9362(.A(n_32216), .Z(n_57187));
	notech_inv i_9352(.A(n_57173), .Z(n_57178));
	notech_inv i_9348(.A(n_57173), .Z(n_57174));
	notech_inv i_9347(.A(n_30590), .Z(n_57173));
	notech_inv i_9344(.A(n_32220), .Z(n_57170));
	notech_inv i_9342(.A(n_32220), .Z(n_57168));
	notech_inv i_9338(.A(n_32220), .Z(n_57164));
	notech_inv i_9336(.A(n_32220), .Z(n_57163));
	notech_inv i_9332(.A(n_32223), .Z(n_57158));
	notech_inv i_9331(.A(n_32223), .Z(n_57157));
	notech_inv i_9325(.A(n_32223), .Z(n_57152));
	notech_inv i_9319(.A(n_32223), .Z(n_57147));
	notech_inv i_9314(.A(n_32224), .Z(n_57141));
	notech_inv i_9308(.A(n_32224), .Z(n_57136));
	notech_inv i_9302(.A(n_32224), .Z(n_57130));
	notech_inv i_9296(.A(n_125342694), .Z(n_57122));
	notech_inv i_9291(.A(n_125342694), .Z(n_57117));
	notech_inv i_9285(.A(n_125342694), .Z(n_57112));
	notech_inv i_9279(.A(n_32311), .Z(n_57103));
	notech_inv i_9274(.A(n_32311), .Z(n_57097));
	notech_inv i_9268(.A(n_32208), .Z(n_57091));
	notech_inv i_9262(.A(n_32208), .Z(n_57086));
	notech_inv i_9256(.A(n_32208), .Z(n_57081));
	notech_inv i_9247(.A(n_57067), .Z(n_57072));
	notech_inv i_9243(.A(n_57067), .Z(n_57068));
	notech_inv i_9242(.A(n_30473), .Z(n_57067));
	notech_inv i_9239(.A(n_32211), .Z(n_57064));
	notech_inv i_9237(.A(n_32211), .Z(n_57062));
	notech_inv i_9234(.A(n_32211), .Z(n_57059));
	notech_inv i_9231(.A(n_32211), .Z(n_57057));
	notech_inv i_9219(.A(n_57044), .Z(n_57045));
	notech_inv i_9218(.A(n_30448), .Z(n_57044));
	notech_inv i_9210(.A(n_57033), .Z(n_57034));
	notech_inv i_9208(.A(n_318871159), .Z(n_57033));
	notech_inv i_9200(.A(n_57018), .Z(n_57024));
	notech_inv i_9195(.A(n_57018), .Z(n_57020));
	notech_inv i_9194(.A(n_4347), .Z(n_57018));
	notech_inv i_9189(.A(n_57000), .Z(n_57012));
	notech_inv i_9184(.A(n_57000), .Z(n_57006));
	notech_inv i_9178(.A(n_57000), .Z(n_57001));
	notech_inv i_9177(.A(n_32196), .Z(n_57000));
	notech_inv i_9169(.A(n_56991), .Z(n_56992));
	notech_inv i_9168(.A(n_318971160), .Z(n_56991));
	notech_inv i_9160(.A(n_56982), .Z(n_56983));
	notech_inv i_9158(.A(n_31478), .Z(n_56982));
	notech_inv i_9150(.A(n_56973), .Z(n_56974));
	notech_inv i_9149(.A(n_31477), .Z(n_56973));
	notech_inv i_9141(.A(n_56964), .Z(n_56965));
	notech_inv i_9140(.A(n_31472), .Z(n_56964));
	notech_inv i_9132(.A(n_56955), .Z(n_56956));
	notech_inv i_9131(.A(n_31473), .Z(n_56955));
	notech_inv i_9129(.A(n_56946), .Z(n_56952));
	notech_inv i_9128(.A(n_56946), .Z(n_56951));
	notech_inv i_9123(.A(n_56946), .Z(n_56947));
	notech_inv i_9122(.A(gs[2]), .Z(n_56946));
	notech_inv i_9112(.A(n_56935), .Z(n_56936));
	notech_inv i_9110(.A(n_98190348), .Z(n_56935));
	notech_inv i_9106(.A(n_56922), .Z(n_56929));
	notech_inv i_9100(.A(n_56922), .Z(n_56923));
	notech_inv i_9099(.A(n_25428), .Z(n_56922));
	notech_inv i_9091(.A(n_56913), .Z(n_56914));
	notech_inv i_9090(.A(n_60316478), .Z(n_56913));
	notech_inv i_9082(.A(n_56903), .Z(n_56904));
	notech_inv i_9081(.A(n_4437), .Z(n_56903));
	notech_inv i_9070(.A(n_56890), .Z(n_56891));
	notech_inv i_9069(.A(n_60516480), .Z(n_56890));
	notech_inv i_9059(.A(n_56879), .Z(n_56880));
	notech_inv i_9058(.A(n_60216477), .Z(n_56879));
	notech_inv i_9050(.A(n_56870), .Z(n_56871));
	notech_inv i_9049(.A(n_59316468), .Z(n_56870));
	notech_inv i_9041(.A(n_56860), .Z(n_56861));
	notech_inv i_9040(.A(n_60916484), .Z(n_56860));
	notech_inv i_9029(.A(n_56849), .Z(n_56850));
	notech_inv i_9028(.A(n_61016485), .Z(n_56849));
	notech_inv i_9020(.A(n_56840), .Z(n_56841));
	notech_inv i_9019(.A(n_4438), .Z(n_56840));
	notech_inv i_9011(.A(n_56831), .Z(n_56832));
	notech_inv i_9010(.A(n_4436), .Z(n_56831));
	notech_inv i_9002(.A(n_56822), .Z(n_56823));
	notech_inv i_9001(.A(n_61716492), .Z(n_56822));
	notech_inv i_8976(.A(n_56791), .Z(n_56792));
	notech_inv i_8974(.A(n_2382), .Z(n_56791));
	notech_inv i_8966(.A(n_56782), .Z(n_56783));
	notech_inv i_8965(.A(n_245877510), .Z(n_56782));
	notech_inv i_8957(.A(n_56773), .Z(n_56774));
	notech_inv i_8956(.A(n_24134), .Z(n_56773));
	notech_inv i_8945(.A(n_56761), .Z(n_56762));
	notech_inv i_8944(.A(n_4447), .Z(n_56761));
	notech_inv i_8933(.A(n_56749), .Z(n_56750));
	notech_inv i_8932(.A(n_24127), .Z(n_56749));
	notech_inv i_8922(.A(n_56737), .Z(n_56738));
	notech_inv i_8921(.A(n_24144), .Z(n_56737));
	notech_inv i_8913(.A(n_56727), .Z(n_56728));
	notech_inv i_8912(.A(n_24138), .Z(n_56727));
	notech_inv i_8904(.A(n_56717), .Z(n_56718));
	notech_inv i_8903(.A(n_24142), .Z(n_56717));
	notech_inv i_8892(.A(n_56706), .Z(n_56707));
	notech_inv i_8891(.A(n_24141), .Z(n_56706));
	notech_inv i_8635(.A(\nbus_11334[0] ), .Z(n_56442));
	notech_inv i_8633(.A(\nbus_11334[0] ), .Z(n_56440));
	notech_inv i_8630(.A(\nbus_11334[0] ), .Z(n_56437));
	notech_inv i_8627(.A(\nbus_11334[0] ), .Z(n_56435));
	notech_inv i_8622(.A(n_56415), .Z(n_56429));
	notech_inv i_8620(.A(n_56415), .Z(n_56428));
	notech_inv i_8614(.A(n_56415), .Z(n_56422));
	notech_inv i_8607(.A(n_56415), .Z(n_56416));
	notech_inv i_8606(.A(n_220280703), .Z(n_56415));
	notech_inv i_8603(.A(n_56402), .Z(n_56412));
	notech_inv i_8602(.A(n_56402), .Z(n_56411));
	notech_inv i_8598(.A(n_56402), .Z(n_56407));
	notech_inv i_8594(.A(n_56402), .Z(n_56404));
	notech_inv i_8593(.A(n_56402), .Z(n_56403));
	notech_inv i_8592(.A(n_315992478), .Z(n_56402));
	notech_inv i_8590(.A(\nbus_11277[0] ), .Z(n_56399));
	notech_inv i_8587(.A(\nbus_11277[0] ), .Z(n_56397));
	notech_inv i_8584(.A(\nbus_11277[0] ), .Z(n_56394));
	notech_inv i_8582(.A(\nbus_11277[0] ), .Z(n_56392));
	notech_inv i_8578(.A(n_56378), .Z(n_56388));
	notech_inv i_8577(.A(n_56378), .Z(n_56387));
	notech_inv i_8572(.A(n_56378), .Z(n_56383));
	notech_inv i_8569(.A(n_56378), .Z(n_56380));
	notech_inv i_8568(.A(n_56378), .Z(n_56379));
	notech_inv i_8567(.A(n_2140), .Z(n_56378));
	notech_inv i_8556(.A(n_56367), .Z(n_56368));
	notech_inv i_8555(.A(n_309892426), .Z(n_56367));
	notech_inv i_8547(.A(n_56358), .Z(n_56359));
	notech_inv i_8546(.A(n_4353), .Z(n_56358));
	notech_inv i_8538(.A(n_56349), .Z(n_56350));
	notech_inv i_8537(.A(n_4352), .Z(n_56349));
	notech_inv i_8529(.A(n_56340), .Z(n_56341));
	notech_inv i_8528(.A(n_4350), .Z(n_56340));
	notech_inv i_8517(.A(n_56329), .Z(n_56330));
	notech_inv i_8515(.A(n_4349), .Z(n_56329));
	notech_inv i_8507(.A(n_56320), .Z(n_56321));
	notech_inv i_8506(.A(n_4424), .Z(n_56320));
	notech_inv i_8467(.A(n_56278), .Z(n_56279));
	notech_inv i_8466(.A(\nbus_11353[0] ), .Z(n_56278));
	notech_inv i_8456(.A(n_56267), .Z(n_56268));
	notech_inv i_8455(.A(n_212333654), .Z(n_56267));
	notech_inv i_8444(.A(n_56256), .Z(n_56257));
	notech_inv i_8441(.A(n_209388005), .Z(n_56256));
	notech_inv i_8430(.A(n_56245), .Z(n_56246));
	notech_inv i_8429(.A(n_30682), .Z(n_56245));
	notech_inv i_8419(.A(n_56234), .Z(n_56235));
	notech_inv i_8418(.A(n_208687999), .Z(n_56234));
	notech_inv i_8410(.A(n_56225), .Z(n_56226));
	notech_inv i_8408(.A(n_207687990), .Z(n_56225));
	notech_inv i_8398(.A(n_56214), .Z(n_56215));
	notech_inv i_8397(.A(n_208587998), .Z(n_56214));
	notech_inv i_8389(.A(n_56205), .Z(n_56206));
	notech_inv i_8388(.A(n_167287599), .Z(n_56205));
	notech_inv i_8380(.A(n_56196), .Z(n_56197));
	notech_inv i_8379(.A(n_207887992), .Z(n_56196));
	notech_inv i_8371(.A(n_56187), .Z(n_56188));
	notech_inv i_8370(.A(n_30683), .Z(n_56187));
	notech_inv i_8258(.A(n_56062), .Z(n_56063));
	notech_inv i_8256(.A(n_98090347), .Z(n_56062));
	notech_inv i_8236(.A(n_56040), .Z(n_56041));
	notech_inv i_8235(.A(n_4456), .Z(n_56040));
	notech_inv i_8231(.A(n_56029), .Z(n_56036));
	notech_inv i_8230(.A(n_56029), .Z(n_56035));
	notech_inv i_8224(.A(n_56029), .Z(n_56030));
	notech_inv i_8223(.A(n_385164382), .Z(n_56029));
	notech_inv i_8213(.A(n_56018), .Z(n_56019));
	notech_inv i_8212(.A(\nbus_11305[0] ), .Z(n_56018));
	notech_inv i_8202(.A(n_56007), .Z(n_56008));
	notech_inv i_8200(.A(n_159362625), .Z(n_56007));
	notech_inv i_8197(.A(n_30788), .Z(n_56003));
	notech_inv i_8196(.A(n_30788), .Z(n_56002));
	notech_inv i_8190(.A(n_30788), .Z(n_55997));
	notech_inv i_8179(.A(n_55985), .Z(n_55986));
	notech_inv i_8178(.A(n_445582455), .Z(n_55985));
	notech_inv i_8167(.A(n_55974), .Z(n_55975));
	notech_inv i_8166(.A(n_126126588), .Z(n_55974));
	notech_inv i_8158(.A(n_55965), .Z(n_55966));
	notech_inv i_8157(.A(n_125926586), .Z(n_55965));
	notech_inv i_8147(.A(n_55954), .Z(n_55955));
	notech_inv i_8146(.A(n_26585), .Z(n_55954));
	notech_inv i_8138(.A(n_55945), .Z(n_55946));
	notech_inv i_8136(.A(n_26600), .Z(n_55945));
	notech_inv i_8126(.A(n_55934), .Z(n_55935));
	notech_inv i_8125(.A(n_164362675), .Z(n_55934));
	notech_inv i_8115(.A(n_55923), .Z(n_55924));
	notech_inv i_8114(.A(n_30961), .Z(n_55923));
	notech_inv i_8103(.A(n_55912), .Z(n_55913));
	notech_inv i_8102(.A(n_330460932), .Z(n_55912));
	notech_inv i_8094(.A(n_55903), .Z(n_55904));
	notech_inv i_8093(.A(n_164196010), .Z(n_55903));
	notech_inv i_8083(.A(n_55892), .Z(n_55893));
	notech_inv i_8082(.A(n_30918), .Z(n_55892));
	notech_inv i_8074(.A(n_55883), .Z(n_55884));
	notech_inv i_8072(.A(n_333360961), .Z(n_55883));
	notech_inv i_8062(.A(n_55872), .Z(n_55873));
	notech_inv i_8061(.A(n_389964430), .Z(n_55872));
	notech_inv i_8051(.A(n_55861), .Z(n_55862));
	notech_inv i_8050(.A(n_442068004), .Z(n_55861));
	notech_inv i_8039(.A(n_55850), .Z(n_55851));
	notech_inv i_8038(.A(n_176766199), .Z(n_55850));
	notech_inv i_8028(.A(n_55839), .Z(n_55840));
	notech_inv i_8027(.A(n_212880631), .Z(n_55839));
	notech_inv i_8019(.A(n_55830), .Z(n_55831));
	notech_inv i_8018(.A(n_323660864), .Z(n_55830));
	notech_inv i_8007(.A(n_55819), .Z(n_55820));
	notech_inv i_8006(.A(n_173966175), .Z(n_55819));
	notech_inv i_7998(.A(n_55810), .Z(n_55811));
	notech_inv i_7997(.A(\nbus_11278[0] ), .Z(n_55810));
	notech_inv i_7989(.A(n_55801), .Z(n_55802));
	notech_inv i_7988(.A(n_5774), .Z(n_55801));
	notech_inv i_7980(.A(n_55792), .Z(n_55793));
	notech_inv i_7979(.A(n_330560933), .Z(n_55792));
	notech_inv i_7959(.A(n_55770), .Z(n_55771));
	notech_inv i_7958(.A(n_30894), .Z(n_55770));
	notech_inv i_7902(.A(n_55656), .Z(n_55657));
	notech_inv i_7901(.A(n_98390350), .Z(n_55656));
	notech_inv i_7891(.A(n_55645), .Z(n_55646));
	notech_inv i_7890(.A(n_98490351), .Z(n_55645));
	notech_inv i_7882(.A(n_55636), .Z(n_55637));
	notech_inv i_7880(.A(n_30738), .Z(n_55636));
	notech_inv i_7872(.A(n_55627), .Z(n_55628));
	notech_inv i_7871(.A(n_447268056), .Z(n_55627));
	notech_inv i_7863(.A(n_55618), .Z(n_55619));
	notech_inv i_7862(.A(n_30744), .Z(n_55618));
	notech_inv i_7854(.A(n_55609), .Z(n_55610));
	notech_inv i_7853(.A(n_447368057), .Z(n_55609));
	notech_inv i_7843(.A(n_55598), .Z(n_55599));
	notech_inv i_7842(.A(\nbus_11320[0] ), .Z(n_55598));
	notech_inv i_7831(.A(n_55587), .Z(n_55588));
	notech_inv i_7830(.A(n_249536174), .Z(n_55587));
	notech_inv i_7822(.A(n_55578), .Z(n_55579));
	notech_inv i_7821(.A(n_194891308), .Z(n_55578));
	notech_inv i_7811(.A(n_55567), .Z(n_55568));
	notech_inv i_7810(.A(n_348389365), .Z(n_55567));
	notech_inv i_7782(.A(n_55494), .Z(n_55495));
	notech_inv i_7781(.A(n_98290349), .Z(n_55494));
	notech_inv i_7701(.A(n_55288), .Z(n_55289));
	notech_inv i_7700(.A(n_31326), .Z(n_55288));
	notech_inv i_7673(.A(n_55257), .Z(n_55258));
	notech_inv i_7671(.A(n_28747367), .Z(n_55257));
	notech_inv i_7661(.A(n_55246), .Z(n_55247));
	notech_inv i_7660(.A(n_29047370), .Z(n_55246));
	notech_inv i_7652(.A(n_55237), .Z(n_55238));
	notech_inv i_7651(.A(n_29347373), .Z(n_55237));
	notech_inv i_7641(.A(n_55226), .Z(n_55227));
	notech_inv i_7639(.A(n_292192264), .Z(n_55226));
	notech_inv i_7631(.A(n_55217), .Z(n_55218));
	notech_inv i_7630(.A(n_292292265), .Z(n_55217));
	notech_inv i_7620(.A(n_55206), .Z(n_55207));
	notech_inv i_7619(.A(n_293792280), .Z(n_55206));
	notech_inv i_7611(.A(n_55197), .Z(n_55198));
	notech_inv i_7610(.A(n_30753), .Z(n_55197));
	notech_inv i_7599(.A(n_55186), .Z(n_55187));
	notech_inv i_7598(.A(n_20898), .Z(n_55186));
	notech_inv i_7590(.A(n_55177), .Z(n_55178));
	notech_inv i_7589(.A(n_20897), .Z(n_55177));
	notech_inv i_7581(.A(n_55168), .Z(n_55169));
	notech_inv i_7580(.A(n_149493977), .Z(n_55168));
	notech_inv i_7570(.A(n_55157), .Z(n_55158));
	notech_inv i_7569(.A(n_149093973), .Z(n_55157));
	notech_inv i_7461(.A(n_55038), .Z(n_55039));
	notech_inv i_7460(.A(n_148793970), .Z(n_55038));
	notech_inv i_7406(.A(n_54978), .Z(n_54979));
	notech_inv i_7405(.A(n_309595536), .Z(n_54978));
	notech_inv i_7395(.A(n_54967), .Z(n_54968));
	notech_inv i_7394(.A(n_309095532), .Z(n_54967));
	notech_inv i_7286(.A(n_54848), .Z(n_54849));
	notech_inv i_7285(.A(n_308695529), .Z(n_54848));
	notech_inv i_7277(.A(n_54839), .Z(n_54840));
	notech_inv i_7276(.A(n_319295608), .Z(n_54839));
	notech_inv i_7266(.A(n_54828), .Z(n_54829));
	notech_inv i_7265(.A(n_318895605), .Z(n_54828));
	notech_inv i_7257(.A(n_54819), .Z(n_54820));
	notech_inv i_7254(.A(n_318295602), .Z(n_54819));
	notech_inv i_7146(.A(n_54700), .Z(n_54701));
	notech_inv i_7145(.A(n_30741), .Z(n_54700));
	notech_inv i_7037(.A(n_54581), .Z(n_54582));
	notech_inv i_7036(.A(n_156394046), .Z(n_54581));
	notech_inv i_7028(.A(n_54572), .Z(n_54573));
	notech_inv i_7027(.A(n_156094043), .Z(n_54572));
	notech_inv i_7018(.A(n_54563), .Z(n_54564));
	notech_inv i_7017(.A(n_163794120), .Z(n_54563));
	notech_inv i_7007(.A(n_54552), .Z(n_54553));
	notech_inv i_7006(.A(n_163394116), .Z(n_54552));
	notech_inv i_6998(.A(n_54543), .Z(n_54544));
	notech_inv i_6996(.A(n_30742), .Z(n_54543));
	notech_inv i_6886(.A(n_54422), .Z(n_54423));
	notech_inv i_6884(.A(n_31293), .Z(n_54422));
	notech_inv i_6874(.A(n_54411), .Z(n_54412));
	notech_inv i_6873(.A(n_125190618), .Z(n_54411));
	notech_inv i_6872(.A(n_54406), .Z(n_54409));
	notech_inv i_6871(.A(n_54406), .Z(n_54408));
	notech_inv i_6870(.A(n_54406), .Z(n_54407));
	notech_inv i_6868(.A(n_279195265), .Z(n_54406));
	notech_inv i_6867(.A(n_54402), .Z(n_54405));
	notech_inv i_6866(.A(n_54402), .Z(n_54404));
	notech_inv i_6865(.A(n_54402), .Z(n_54403));
	notech_inv i_6864(.A(n_279195265), .Z(n_54402));
	notech_inv i_6863(.A(n_54397), .Z(n_54400));
	notech_inv i_6862(.A(n_54397), .Z(n_54399));
	notech_inv i_6860(.A(n_54397), .Z(n_54398));
	notech_inv i_6859(.A(n_30749), .Z(n_54397));
	notech_inv i_6858(.A(n_54393), .Z(n_54396));
	notech_inv i_6857(.A(n_54393), .Z(n_54395));
	notech_inv i_6856(.A(n_54393), .Z(n_54394));
	notech_inv i_6855(.A(n_30749), .Z(n_54393));
	notech_inv i_6854(.A(n_54387), .Z(n_54391));
	notech_inv i_6852(.A(n_54387), .Z(n_54390));
	notech_inv i_6851(.A(n_54387), .Z(n_54389));
	notech_inv i_6850(.A(n_54387), .Z(n_54388));
	notech_inv i_6849(.A(n_280395276), .Z(n_54387));
	notech_inv i_6848(.A(n_54382), .Z(n_54386));
	notech_inv i_6847(.A(n_54382), .Z(n_54385));
	notech_inv i_6846(.A(n_54382), .Z(n_54384));
	notech_inv i_6844(.A(n_54382), .Z(n_54383));
	notech_inv i_6843(.A(n_280395276), .Z(n_54382));
	notech_inv i_6842(.A(n_54377), .Z(n_54380));
	notech_inv i_6841(.A(n_54377), .Z(n_54379));
	notech_inv i_6840(.A(n_54377), .Z(n_54378));
	notech_inv i_6839(.A(n_280295275), .Z(n_54377));
	notech_inv i_6838(.A(n_54373), .Z(n_54376));
	notech_inv i_6836(.A(n_54373), .Z(n_54375));
	notech_inv i_6835(.A(n_54373), .Z(n_54374));
	notech_inv i_6834(.A(n_280295275), .Z(n_54373));
	notech_inv i_6833(.A(n_54367), .Z(n_54371));
	notech_inv i_6832(.A(n_54367), .Z(n_54370));
	notech_inv i_6831(.A(n_54367), .Z(n_54369));
	notech_inv i_6830(.A(n_54367), .Z(n_54368));
	notech_inv i_6828(.A(n_279895271), .Z(n_54367));
	notech_inv i_6827(.A(n_54362), .Z(n_54366));
	notech_inv i_6826(.A(n_54362), .Z(n_54365));
	notech_inv i_6825(.A(n_54362), .Z(n_54364));
	notech_inv i_6824(.A(n_54362), .Z(n_54363));
	notech_inv i_6823(.A(n_279895271), .Z(n_54362));
	notech_inv i_6822(.A(n_54357), .Z(n_54360));
	notech_inv i_6820(.A(n_54357), .Z(n_54359));
	notech_inv i_6819(.A(n_54357), .Z(n_54358));
	notech_inv i_6818(.A(n_279795270), .Z(n_54357));
	notech_inv i_6817(.A(n_54353), .Z(n_54356));
	notech_inv i_6816(.A(n_54353), .Z(n_54355));
	notech_inv i_6815(.A(n_54353), .Z(n_54354));
	notech_inv i_6814(.A(n_279795270), .Z(n_54353));
	notech_inv i_6812(.A(n_54347), .Z(n_54351));
	notech_inv i_6811(.A(n_54347), .Z(n_54350));
	notech_inv i_6810(.A(n_54347), .Z(n_54349));
	notech_inv i_6809(.A(n_54347), .Z(n_54348));
	notech_inv i_6808(.A(n_279395267), .Z(n_54347));
	notech_inv i_6807(.A(n_54342), .Z(n_54346));
	notech_inv i_6806(.A(n_54342), .Z(n_54345));
	notech_inv i_6804(.A(n_54342), .Z(n_54344));
	notech_inv i_6803(.A(n_54342), .Z(n_54343));
	notech_inv i_6802(.A(n_279395267), .Z(n_54342));
	notech_inv i_6801(.A(n_54337), .Z(n_54340));
	notech_inv i_6800(.A(n_54337), .Z(n_54339));
	notech_inv i_6799(.A(n_54337), .Z(n_54338));
	notech_inv i_6798(.A(n_278895262), .Z(n_54337));
	notech_inv i_6796(.A(n_54333), .Z(n_54336));
	notech_inv i_6795(.A(n_54333), .Z(n_54335));
	notech_inv i_6794(.A(n_54333), .Z(n_54334));
	notech_inv i_6793(.A(n_278895262), .Z(n_54333));
	notech_inv i_6792(.A(n_54328), .Z(n_54331));
	notech_inv i_6791(.A(n_54328), .Z(n_54330));
	notech_inv i_6790(.A(n_54328), .Z(n_54329));
	notech_inv i_6788(.A(n_114590512), .Z(n_54328));
	notech_inv i_6787(.A(n_54324), .Z(n_54327));
	notech_inv i_6786(.A(n_54324), .Z(n_54326));
	notech_inv i_6785(.A(n_54324), .Z(n_54325));
	notech_inv i_6784(.A(n_114590512), .Z(n_54324));
	notech_inv i_6783(.A(n_54319), .Z(n_54322));
	notech_inv i_6782(.A(n_54319), .Z(n_54321));
	notech_inv i_6780(.A(n_54319), .Z(n_54320));
	notech_inv i_6779(.A(n_30724), .Z(n_54319));
	notech_inv i_6778(.A(n_54315), .Z(n_54318));
	notech_inv i_6777(.A(n_54315), .Z(n_54317));
	notech_inv i_6776(.A(n_54315), .Z(n_54316));
	notech_inv i_6775(.A(n_30724), .Z(n_54315));
	notech_inv i_6774(.A(n_54309), .Z(n_54313));
	notech_inv i_6772(.A(n_54309), .Z(n_54312));
	notech_inv i_6771(.A(n_54309), .Z(n_54311));
	notech_inv i_6770(.A(n_54309), .Z(n_54310));
	notech_inv i_6769(.A(n_115190518), .Z(n_54309));
	notech_inv i_6768(.A(n_54304), .Z(n_54308));
	notech_inv i_6767(.A(n_54304), .Z(n_54307));
	notech_inv i_6766(.A(n_54304), .Z(n_54306));
	notech_inv i_6764(.A(n_54304), .Z(n_54305));
	notech_inv i_6763(.A(n_115190518), .Z(n_54304));
	notech_inv i_6762(.A(n_54299), .Z(n_54302));
	notech_inv i_6761(.A(n_54299), .Z(n_54301));
	notech_inv i_6760(.A(n_54299), .Z(n_54300));
	notech_inv i_6759(.A(n_115090517), .Z(n_54299));
	notech_inv i_6758(.A(n_54295), .Z(n_54298));
	notech_inv i_6756(.A(n_54295), .Z(n_54297));
	notech_inv i_6755(.A(n_54295), .Z(n_54296));
	notech_inv i_6754(.A(n_115090517), .Z(n_54295));
	notech_inv i_6753(.A(n_54289), .Z(n_54293));
	notech_inv i_6752(.A(n_54289), .Z(n_54292));
	notech_inv i_6751(.A(n_54289), .Z(n_54291));
	notech_inv i_6750(.A(n_54289), .Z(n_54290));
	notech_inv i_6748(.A(n_114990516), .Z(n_54289));
	notech_inv i_6747(.A(n_54284), .Z(n_54288));
	notech_inv i_6746(.A(n_54284), .Z(n_54287));
	notech_inv i_6745(.A(n_54284), .Z(n_54286));
	notech_inv i_6744(.A(n_54284), .Z(n_54285));
	notech_inv i_6743(.A(n_114990516), .Z(n_54284));
	notech_inv i_6742(.A(n_54279), .Z(n_54282));
	notech_inv i_6740(.A(n_54279), .Z(n_54281));
	notech_inv i_6739(.A(n_54279), .Z(n_54280));
	notech_inv i_6738(.A(n_114790514), .Z(n_54279));
	notech_inv i_6737(.A(n_54275), .Z(n_54278));
	notech_inv i_6736(.A(n_54275), .Z(n_54277));
	notech_inv i_6735(.A(n_54275), .Z(n_54276));
	notech_inv i_6734(.A(n_114790514), .Z(n_54275));
	notech_inv i_6732(.A(n_54269), .Z(n_54273));
	notech_inv i_6731(.A(n_54269), .Z(n_54272));
	notech_inv i_6730(.A(n_54269), .Z(n_54271));
	notech_inv i_6729(.A(n_54269), .Z(n_54270));
	notech_inv i_6728(.A(n_114290509), .Z(n_54269));
	notech_inv i_6727(.A(n_54264), .Z(n_54268));
	notech_inv i_6726(.A(n_54264), .Z(n_54267));
	notech_inv i_6724(.A(n_54264), .Z(n_54266));
	notech_inv i_6723(.A(n_54264), .Z(n_54265));
	notech_inv i_6722(.A(n_114290509), .Z(n_54264));
	notech_inv i_6721(.A(n_54151), .Z(n_54154));
	notech_inv i_6720(.A(n_54151), .Z(n_54153));
	notech_inv i_6719(.A(n_54151), .Z(n_54152));
	notech_inv i_6718(.A(n_114090507), .Z(n_54151));
	notech_inv i_6716(.A(n_54147), .Z(n_54150));
	notech_inv i_6715(.A(n_54147), .Z(n_54149));
	notech_inv i_6714(.A(n_54147), .Z(n_54148));
	notech_inv i_6713(.A(n_114090507), .Z(n_54147));
	notech_nao3 i_188387608(.A(n_347671363), .B(n_30336), .C(n_349371378), .Z
		(n_349971384));
	notech_nao3 i_206687607(.A(n_63818), .B(n_61823), .C(n_32575), .Z(n_544)
		);
	notech_ao4 i_148187604(.A(n_60157), .B(n_30305), .C(n_60194), .D(n_3452)
		, .Z(n_349871383));
	notech_and4 i_51761(.A(fsm[4]), .B(fsm[2]), .C(fsm[3]), .D(n_316260790),
		 .Z(n_349671381));
	notech_and4 i_51763(.A(fsm[4]), .B(fsm[2]), .C(fsm[3]), .D(n_32520), .Z(n_59560
		));
	notech_and2 i_182987602(.A(n_349871383), .B(n_341771329), .Z(n_349571380
		));
	notech_ao4 i_116587601(.A(n_60175), .B(n_30305), .C(n_32394), .D(n_315360781
		), .Z(n_57340));
	notech_or2 i_51758(.A(n_301560644), .B(n_316160789), .Z(n_349471379));
	notech_nand2 i_26899(.A(n_349471379), .B(n_347271361), .Z(n_349371378)
		);
	notech_and2 i_137787599(.A(n_32628), .B(n_32391), .Z(n_349271377));
	notech_or4 i_194987598(.A(n_32576), .B(n_32397), .C(n_32184), .D(n_32391
		), .Z(n_349171376));
	notech_or4 i_156087597(.A(n_32396), .B(n_28534), .C(n_61935), .D(n_61959
		), .Z(n_349071375));
	notech_or4 i_104587594(.A(n_32391), .B(n_309960727), .C(n_314960777), .D
		(n_61056), .Z(n_348771372));
	notech_or2 i_157387593(.A(n_32484), .B(n_30712), .Z(n_348571371));
	notech_nao3 i_178687592(.A(n_30681), .B(n_30382), .C(n_349971384), .Z(n_348471370
		));
	notech_and2 i_75287591(.A(n_348771372), .B(n_23326), .Z(n_348271368));
	notech_and2 i_148487590(.A(n_349171376), .B(n_1847), .Z(n_348171367));
	notech_and2 i_137287589(.A(n_349071375), .B(n_57283), .Z(n_348071366));
	notech_nand2 i_169687588(.A(n_32514), .B(n_32506), .Z(n_347971365));
	notech_nand3 i_26900(.A(n_349471379), .B(n_347271361), .C(n_30336), .Z(n_347771364
		));
	notech_nao3 i_51760(.A(n_61917), .B(n_61901), .C(n_316160789), .Z(n_347671363
		));
	notech_nao3 i_178487587(.A(n_32646), .B(n_61823), .C(n_32575), .Z(n_347471362
		));
	notech_nao3 i_145837488(.A(n_315760785), .B(n_30650), .C(n_301560644), .Z
		(n_2036));
	notech_or2 i_51757(.A(n_316160789), .B(n_30304), .Z(n_347271361));
	notech_nao3 i_161887585(.A(n_32646), .B(n_63800), .C(n_49651676), .Z(n_49351679
		));
	notech_or2 i_192437456(.A(n_312671105), .B(n_30670), .Z(n_2004));
	notech_or4 i_205637477(.A(n_59114), .B(n_19725), .C(n_30330), .D(n_61870
		), .Z(n_2025));
	notech_ao4 i_152437484(.A(n_2091), .B(n_30383), .C(n_30374), .D(n_2081),
		 .Z(n_2032));
	notech_nand2 i_61537533(.A(n_32506), .B(n_30650), .Z(n_2081));
	notech_or2 i_41937545(.A(n_19707), .B(n_61688), .Z(n_2094));
	notech_nand2 i_3120701(.A(n_341071324), .B(n_340571319), .Z(n_20074));
	notech_or4 i_169437559(.A(n_32589), .B(n_28534), .C(n_63700), .D(n_63794
		), .Z(n_2111));
	notech_or4 i_168937560(.A(n_32589), .B(n_28008), .C(\opcode[1] ), .D(\opcode[2] 
		), .Z(n_2112));
	notech_nao3 i_122237561(.A(n_3368), .B(n_323071195), .C(n_323171196), .Z
		(n_2113));
	notech_and4 i_80437590(.A(n_3326), .B(n_2032), .C(n_57016), .D(n_56582),
		 .Z(n_57681));
	notech_nor2 i_37013(.A(n_56867), .B(n_53445), .Z(n_2130));
	notech_ao4 i_183437470(.A(n_3456), .B(n_33321), .C(n_61845), .D(n_57019)
		, .Z(n_2018));
	notech_nand3 i_180737471(.A(n_323771202), .B(n_315171127), .C(n_323871203
		), .Z(n_2019));
	notech_or4 i_79637591(.A(n_2091), .B(n_347671363), .C(n_347971365), .D(n_347771364
		), .Z(n_57688));
	notech_or2 i_203637592(.A(n_311371095), .B(n_30307), .Z(n_56603));
	notech_and2 i_56137541(.A(n_316471137), .B(n_30560), .Z(n_2090));
	notech_ao4 i_152337593(.A(n_2091), .B(n_347271361), .C(n_30636), .D(n_2081
		), .Z(n_57016));
	notech_and2 i_56537594(.A(n_48030), .B(n_315271128), .Z(n_57915));
	notech_nand2 i_47863(.A(n_316571138), .B(n_57724), .Z(n_10054));
	notech_or4 i_31400(.A(n_61935), .B(n_61959), .C(n_61870), .D(n_61625), .Z
		(n_2152));
	notech_and4 i_162837478(.A(n_61959), .B(n_61935), .C(n_61099), .D(n_61688
		), .Z(n_2026));
	notech_or2 i_100137640(.A(n_311171093), .B(n_57449), .Z(n_57501));
	notech_and4 i_12137644(.A(instrc[119]), .B(instrc[118]), .C(n_33152), .D
		(instrc[117]), .Z(n_58274));
	notech_and2 i_176037645(.A(n_33152), .B(instrc[117]), .Z(n_56820));
	notech_and4 i_170437650(.A(n_30636), .B(n_30374), .C(n_19629), .D(n_30377
		), .Z(n_56867));
	notech_nand2 i_140737491(.A(n_30374), .B(n_30636), .Z(n_2039));
	notech_or4 i_27034(.A(n_49651676), .B(n_32383), .C(\opcode[2] ), .D(n_61959
		), .Z(n_2178));
	notech_and3 i_68237653(.A(n_32386), .B(n_3457), .C(n_1850), .Z(n_57799)
		);
	notech_or4 i_204987581(.A(n_32575), .B(n_60175), .C(n_32646), .D(\opcode[3] 
		), .Z(n_347071359));
	notech_or4 i_196237654(.A(n_32575), .B(n_32628), .C(n_60175), .D(n_31407
		), .Z(n_56663));
	notech_nao3 i_55937542(.A(n_32481), .B(n_61625), .C(n_32484), .Z(n_2091)
		);
	notech_ao4 i_152237485(.A(n_329571252), .B(n_329671253), .C(n_32573), .D
		(n_60157), .Z(n_2033));
	notech_nao3 i_206037656(.A(n_63212389), .B(\opcode[0] ), .C(n_329571252)
		, .Z(n_59515));
	notech_or4 i_50337(.A(n_61889), .B(n_59515), .C(n_61723), .D(n_61870), .Z
		(n_59599));
	notech_or4 i_206237698(.A(n_61889), .B(n_30304), .C(n_316260790), .D(n_61870
		), .Z(n_56582));
	notech_or4 i_9209(.A(n_311371095), .B(n_61723), .C(n_301960648), .D(n_19725
		), .Z(n_50148));
	notech_or4 i_81037699(.A(n_60175), .B(n_61845), .C(n_544), .D(n_31407), 
		.Z(n_57675));
	notech_or4 i_80737700(.A(n_30323), .B(n_2091), .C(n_322771192), .D(n_30324
		), .Z(n_57678));
	notech_or4 i_146187580(.A(n_32391), .B(n_309960727), .C(n_314960777), .D
		(n_60175), .Z(n_3469));
	notech_or4 i_76537701(.A(n_314960777), .B(n_28098), .C(n_76712523), .D(n_60175
		), .Z(n_57717));
	notech_and3 i_97737706(.A(n_321871184), .B(n_321971185), .C(n_60157), .Z
		(n_57521));
	notech_mux2 i_3111677(.S(n_61284), .A(regs_14[30]), .B(add_len_pc32[30])
		, .Z(\add_len_pc[30] ));
	notech_nao3 i_31837709(.A(n_32186), .B(n_339871312), .C(n_2004), .Z(n_5680
		));
	notech_and4 i_145329822(.A(n_3395), .B(n_339471310), .C(n_3390), .D(n_3393
		), .Z(n_5750));
	notech_or4 i_11327(.A(n_60194), .B(n_32576), .C(n_32184), .D(n_32391), .Z
		(n_48030));
	notech_or4 i_5878(.A(n_61889), .B(n_57749), .C(n_61723), .D(n_61870), .Z
		(n_53429));
	notech_and2 i_151937732(.A(n_57799), .B(n_314971125), .Z(n_57019));
	notech_ao3 i_5862(.A(n_61099), .B(n_61688), .C(n_57099), .Z(n_53445));
	notech_and3 i_141437733(.A(n_30560), .B(n_316471137), .C(n_316271135), .Z
		(n_57099));
	notech_nand3 i_184337748(.A(n_61901), .B(n_61917), .C(n_315760785), .Z(n_56755
		));
	notech_or4 i_149437754(.A(n_61889), .B(n_57340), .C(n_61723), .D(n_61870
		), .Z(n_57041));
	notech_or4 i_179137755(.A(n_32383), .B(n_309960727), .C(n_314960777), .D
		(n_60157), .Z(n_56794));
	notech_nao3 i_205537761(.A(n_32646), .B(n_63212389), .C(n_329571252), .Z
		(n_59516));
	notech_or4 i_75737774(.A(n_311071092), .B(n_19548), .C(n_313471111), .D(n_2113
		), .Z(n_57724));
	notech_nand3 i_50458(.A(n_331971276), .B(n_330171258), .C(n_3381), .Z(\nbus_11314[0] 
		));
	notech_nand2 i_130640117(.A(nbus_11271[0]), .B(nbus_11271[1]), .Z(n_57206
		));
	notech_and2 i_129040118(.A(opc[0]), .B(opc[1]), .Z(n_57222));
	notech_nand3 i_139440079(.A(opc[0]), .B(opc[1]), .C(opc[2]), .Z(n_317051260
		));
	notech_nand2 i_207540139(.A(rep_en2), .B(n_30937), .Z(n_56572));
	notech_or4 i_196540140(.A(rep_en3), .B(rep_en2), .C(rep_en1), .D(rep_en4
		), .Z(n_56661));
	notech_or4 i_162740142(.A(rep_en3), .B(rep_en2), .C(rep_en1), .D(n_30938
		), .Z(n_56930));
	notech_nao3 i_116940145(.A(rep_en3), .B(n_30937), .C(rep_en2), .Z(n_57336
		));
	notech_nand2 i_141043282(.A(n_31604), .B(n_31605), .Z(n_320851229));
	notech_and4 i_94229174(.A(n_308971072), .B(n_308871071), .C(n_308371067)
		, .D(n_308771070), .Z(n_5243));
	notech_and4 i_93829170(.A(n_307471058), .B(n_307371057), .C(n_306971053)
		, .D(n_307271056), .Z(n_5711));
	notech_and4 i_93729169(.A(n_305971044), .B(n_305871043), .C(n_305471039)
		, .D(n_305771042), .Z(n_5720));
	notech_and4 i_93029163(.A(n_299870988), .B(n_299670987), .C(n_299270983)
		, .D(n_299570986), .Z(n_5356));
	notech_and4 i_92929162(.A(n_298370974), .B(n_298270973), .C(n_297870969)
		, .D(n_298170972), .Z(n_5436));
	notech_and4 i_92829161(.A(n_296970960), .B(n_296870959), .C(n_296470955)
		, .D(n_296770958), .Z(n_5397));
	notech_and4 i_92743349(.A(n_295570946), .B(n_295470945), .C(n_295070941)
		, .D(n_295370944), .Z(n_5444));
	notech_and4 i_91943355(.A(n_294170932), .B(n_294070931), .C(n_293670927)
		, .D(n_293970930), .Z(n_5269));
	notech_and4 i_94129173(.A(n_292670917), .B(n_292570916), .C(n_292170912)
		, .D(n_292470915), .Z(n_5758));
	notech_nand3 i_8948(.A(n_31604), .B(n_31605), .C(opz[2]), .Z(n_50409));
	notech_nand2 i_119543369(.A(n_50409), .B(n_272170713), .Z(n_59558));
	notech_and4 i_145429833(.A(n_263670631), .B(n_263570630), .C(n_263170626
		), .D(n_263470629), .Z(n_300822033));
	notech_nao3 i_45346425(.A(n_321271180), .B(n_311471096), .C(n_321371181)
		, .Z(n_300322028));
	notech_and2 i_126646414(.A(n_309671079), .B(n_251470509), .Z(n_299222017
		));
	notech_and2 i_110946416(.A(n_310171083), .B(n_262270617), .Z(n_299422019
		));
	notech_nand2 i_120671(.A(n_272070712), .B(n_271570707), .Z(n_19894));
	notech_nand2 i_220672(.A(n_270970702), .B(n_270370696), .Z(n_19900));
	notech_nand2 i_920679(.A(n_269770690), .B(n_267770670), .Z(n_19942));
	notech_nand2 i_1520685(.A(n_266770660), .B(n_266270655), .Z(n_19978));
	notech_nand2 i_3220702(.A(n_264870643), .B(n_264370638), .Z(n_20080));
	notech_and4 i_143146429(.A(n_268970682), .B(n_268870681), .C(n_268470677
		), .D(n_268770680), .Z(n_300722032));
	notech_mux2 i_3211678(.S(n_61284), .A(regs_14[31]), .B(add_len_pc32[31])
		, .Z(\add_len_pc[31] ));
	notech_mux2 i_1511661(.S(n_61284), .A(n_532), .B(add_len_pc32[14]), .Z(\add_len_pc[14] 
		));
	notech_mux2 i_911655(.S(n_61284), .A(n_526), .B(add_len_pc32[8]), .Z(\add_len_pc[8] 
		));
	notech_mux2 i_211648(.S(n_61284), .A(n_519), .B(add_len_pc32[1]), .Z(\add_len_pc[1] 
		));
	notech_mux2 i_111647(.S(n_61284), .A(n_518), .B(add_len_pc32[0]), .Z(\add_len_pc[0] 
		));
	notech_and4 i_144229700(.A(n_234070336), .B(n_233970335), .C(n_233570331
		), .D(n_233870334), .Z(n_319725273));
	notech_ao3 i_43846448(.A(n_309871081), .B(n_311471096), .C(n_321371181),
		 .Z(n_58042));
	notech_and2 i_106446450(.A(n_310271084), .B(n_262270617), .Z(n_57441));
	notech_and4 i_416994(.A(n_248770482), .B(n_248670481), .C(n_249770492), 
		.D(n_248570480), .Z(n_11953));
	notech_nand2 i_1717007(.A(n_248170476), .B(n_247670471), .Z(n_12031));
	notech_nand2 i_1917009(.A(n_247170466), .B(n_246670461), .Z(n_12043));
	notech_nand2 i_720677(.A(n_245970455), .B(n_245270448), .Z(n_19930));
	notech_nand2 i_820678(.A(n_244570441), .B(n_243870434), .Z(n_19936));
	notech_nand2 i_1720687(.A(n_242770423), .B(n_242270418), .Z(n_19990));
	notech_nand2 i_1820688(.A(n_240270398), .B(n_239770393), .Z(n_19996));
	notech_nand2 i_1920689(.A(n_237770373), .B(n_237270368), .Z(n_20002));
	notech_nand2 i_2020690(.A(n_235270348), .B(n_234770343), .Z(n_20008));
	notech_and4 i_144129691(.A(n_236570361), .B(n_236470360), .C(n_236070356
		), .D(n_236370359), .Z(n_319825274));
	notech_and4 i_144029680(.A(n_239070386), .B(n_238970385), .C(n_238570381
		), .D(n_238870384), .Z(n_319951172));
	notech_and4 i_143929669(.A(n_241570411), .B(n_241470410), .C(n_241070406
		), .D(n_241370409), .Z(n_320051171));
	notech_mux2 i_2011666(.S(n_61284), .A(regs_14[19]), .B(add_len_pc32[19])
		, .Z(\add_len_pc[19] ));
	notech_mux2 i_1911665(.S(n_61284), .A(regs_14[18]), .B(add_len_pc32[18])
		, .Z(\add_len_pc[18] ));
	notech_mux2 i_1811664(.S(n_61284), .A(regs_14[17]), .B(add_len_pc32[17])
		, .Z(\add_len_pc[17] ));
	notech_mux2 i_1711663(.S(n_61281), .A(regs_14[16]), .B(add_len_pc32[16])
		, .Z(\add_len_pc[16] ));
	notech_mux2 i_811654(.S(n_61281), .A(n_525), .B(add_len_pc32[7]), .Z(\add_len_pc[7] 
		));
	notech_mux2 i_711653(.S(n_61281), .A(n_524), .B(add_len_pc32[6]), .Z(\add_len_pc[6] 
		));
	notech_and4 i_93329166(.A(n_304471030), .B(n_304371029), .C(n_303971025)
		, .D(n_304271028), .Z(n_59464));
	notech_and4 i_93229165(.A(n_302971016), .B(n_302871015), .C(n_302471011)
		, .D(n_302771014), .Z(n_59465));
	notech_and4 i_93129164(.A(n_301271002), .B(n_301171001), .C(n_300770997)
		, .D(n_301071000), .Z(n_59466));
	notech_and4 i_144329711(.A(n_208570097), .B(n_208470096), .C(n_207970092
		), .D(n_208370095), .Z(n_346771358));
	notech_and4 i_144429722(.A(n_206070073), .B(n_205970072), .C(n_205570068
		), .D(n_205870071), .Z(n_3466));
	notech_and4 i_144529734(.A(n_203170049), .B(n_203070048), .C(n_202470044
		), .D(n_202970047), .Z(n_3464));
	notech_or4 i_20667(.A(n_2383), .B(n_32159), .C(n_32161), .D(n_33157), .Z
		(n_38705));
	notech_mux2 i_2611672(.S(n_61281), .A(regs_14[25]), .B(add_len_pc32[25])
		, .Z(n_3463));
	notech_mux2 i_2511671(.S(n_61281), .A(regs_14[24]), .B(add_len_pc32[24])
		, .Z(n_3462));
	notech_mux2 i_2411670(.S(n_61281), .A(regs_14[23]), .B(add_len_pc32[23])
		, .Z(n_3461));
	notech_mux2 i_2311669(.S(n_61281), .A(regs_14[22]), .B(add_len_pc32[22])
		, .Z(n_3460));
	notech_mux2 i_2211668(.S(n_61281), .A(regs_14[21]), .B(add_len_pc32[21])
		, .Z(n_3459));
	notech_mux2 i_2111667(.S(n_61281), .A(regs_14[20]), .B(add_len_pc32[20])
		, .Z(n_3458));
	notech_and4 i_145029791(.A(n_173869774), .B(n_173769773), .C(n_173369769
		), .D(n_173669772), .Z(n_284131522));
	notech_and4 i_144929780(.A(n_176369799), .B(n_176269798), .C(n_175869794
		), .D(n_176169797), .Z(n_284231523));
	notech_nand2 i_2717017(.A(n_182269856), .B(n_181669851), .Z(n_12091));
	notech_nand2 i_2817018(.A(n_181169846), .B(n_180669841), .Z(n_12097));
	notech_nand2 i_3017020(.A(n_180169836), .B(n_179569831), .Z(n_12109));
	notech_and4 i_721349(.A(n_178169817), .B(n_178069816), .C(n_179069826), 
		.D(n_177969815), .Z(n_20420));
	notech_nand2 i_2720697(.A(n_177569811), .B(n_177069806), .Z(n_20050));
	notech_nand2 i_2820698(.A(n_175069786), .B(n_174569781), .Z(n_20056));
	notech_nand2 i_2920699(.A(n_172569761), .B(n_171869756), .Z(n_20062));
	notech_nand2 i_3020700(.A(n_171369751), .B(n_170869746), .Z(n_20068));
	notech_or4 i_19088(.A(opa[7]), .B(n_30270), .C(n_27835), .D(n_156269600)
		, .Z(n_40282));
	notech_mux2 i_3011676(.S(n_61281), .A(regs_14[29]), .B(add_len_pc32[29])
		, .Z(\add_len_pc[29] ));
	notech_mux2 i_2911675(.S(n_61286), .A(regs_14[28]), .B(add_len_pc32[28])
		, .Z(\add_len_pc[28] ));
	notech_mux2 i_2811674(.S(n_61286), .A(regs_14[27]), .B(add_len_pc32[27])
		, .Z(\add_len_pc[27] ));
	notech_mux2 i_2711673(.S(n_61286), .A(regs_14[26]), .B(add_len_pc32[26])
		, .Z(\add_len_pc[26] ));
	notech_ao4 i_165355966(.A(n_27835), .B(n_57657), .C(n_30368), .D(n_57679
		), .Z(n_56908));
	notech_nand2 i_3117021(.A(n_156069598), .B(n_155569593), .Z(n_12115));
	notech_and4 i_721893(.A(n_154569583), .B(n_154469582), .C(n_154369581), 
		.D(n_154969587), .Z(n_12328));
	notech_and3 i_105460718(.A(n_116742608), .B(n_58218), .C(n_180276862), .Z
		(n_57450));
	notech_and2 i_106760767(.A(n_324078249), .B(n_57450), .Z(n_57438));
	notech_and2 i_43560772(.A(n_58083), .B(n_151169549), .Z(n_5783));
	notech_or4 i_42560774(.A(n_61723), .B(n_61889), .C(n_383264363), .D(n_61870
		), .Z(n_58055));
	notech_or4 i_38660780(.A(n_61912), .B(n_61901), .C(n_61889), .D(n_383264363
		), .Z(n_5774));
	notech_nand2 i_717573(.A(n_150869546), .B(n_150269540), .Z(n_11602));
	notech_and4 i_216992(.A(n_148669524), .B(n_148569523), .C(n_149569533), 
		.D(n_148469522), .Z(n_11941));
	notech_and4 i_716997(.A(n_147069508), .B(n_146969507), .C(n_148069518), 
		.D(n_146869506), .Z(n_11971));
	notech_and4 i_1517005(.A(n_146069498), .B(n_145969497), .C(n_145869496),
		 .D(n_146369501), .Z(n_12019));
	notech_nand2 i_721829(.A(n_145069488), .B(n_144469482), .Z(n_12680));
	notech_and4 i_721765(.A(n_134869386), .B(n_134769385), .C(n_134269380), 
		.D(n_134669384), .Z(n_15206));
	notech_and4 i_721509(.A(n_132869366), .B(n_132769365), .C(n_133269370), 
		.D(n_132669364), .Z(n_15558));
	notech_and4 i_721317(.A(n_131369351), .B(n_131269350), .C(n_131869356), 
		.D(n_131169349), .Z(n_15910));
	notech_nand2 i_721061(.A(n_130469342), .B(n_129869336), .Z(n_16259));
	notech_nand2 i_720997(.A(n_129269330), .B(n_128669324), .Z(n_18560));
	notech_or4 i_196671995(.A(n_49651676), .B(n_32383), .C(n_61056), .D(reps
		[2]), .Z(n_3457));
	notech_or4 i_69171997(.A(n_348471370), .B(n_59560), .C(n_2091), .D(n_30364
		), .Z(n_3456));
	notech_and2 i_49387572(.A(n_1817), .B(n_59502), .Z(n_3455));
	notech_nao3 i_20887569(.A(n_63818), .B(\opcode[3] ), .C(n_49651676), .Z(n_3452
		));
	notech_or4 i_52987568(.A(n_32663), .B(n_309860726), .C(n_312460752), .D(n_2952
		), .Z(n_49651676));
	notech_or4 i_41387566(.A(ecx[16]), .B(ecx[17]), .C(ecx[19]), .D(ecx[18])
		, .Z(n_3450));
	notech_or4 i_41287563(.A(ecx[21]), .B(ecx[23]), .C(ecx[20]), .D(ecx[22])
		, .Z(n_344671355));
	notech_or4 i_41187559(.A(ecx[25]), .B(ecx[24]), .C(ecx[27]), .D(ecx[26])
		, .Z(n_344271352));
	notech_or4 i_41087556(.A(ecx[29]), .B(ecx[28]), .C(ecx[30]), .D(ecx[31])
		, .Z(n_3439));
	notech_or4 i_39987552(.A(ecx[1]), .B(ecx[0]), .C(ecx[3]), .D(ecx[2]), .Z
		(n_343471345));
	notech_or4 i_39887549(.A(ecx[7]), .B(ecx[5]), .C(ecx[4]), .D(ecx[6]), .Z
		(n_343171342));
	notech_or4 i_40087546(.A(ecx[9]), .B(ecx[8]), .C(n_342471336), .D(n_342371335
		), .Z(n_342771339));
	notech_nand2 i_39087543(.A(n_31419), .B(n_31418), .Z(n_342471336));
	notech_or4 i_39687542(.A(ecx[13]), .B(ecx[12]), .C(ecx[15]), .D(ecx[14])
		, .Z(n_342371335));
	notech_and2 i_140887537(.A(n_349471379), .B(n_30681), .Z(n_57105));
	notech_or4 i_2205(.A(n_49651676), .B(n_32397), .C(n_32646), .D(n_61823),
		 .Z(n_59502));
	notech_ao3 i_131987536(.A(n_30287), .B(n_1850), .C(n_1854), .Z(n_57194)
		);
	notech_and3 i_73287535(.A(n_57340), .B(n_349571380), .C(n_341871330), .Z
		(n_57749));
	notech_or4 i_46287534(.A(n_49651676), .B(n_32397), .C(\opcode[0] ), .D(n_61823
		), .Z(n_341871330));
	notech_or4 i_46087533(.A(n_49651676), .B(n_60194), .C(\opcode[0] ), .D(n_61823
		), .Z(n_341771329));
	notech_or4 i_15856(.A(n_49651676), .B(n_32383), .C(\opcode[1] ), .D(n_61935
		), .Z(n_3415));
	notech_or4 i_2687531(.A(n_3450), .B(n_344671355), .C(n_3439), .D(n_344271352
		), .Z(n_341471327));
	notech_and2 i_41687530(.A(n_61286), .B(n_341471327), .Z(n_341271326));
	notech_ao4 i_122987529(.A(n_315460782), .B(n_60175), .C(n_27924), .D(n_32397
		), .Z(n_57283));
	notech_or4 i_587527(.A(n_343171342), .B(n_343471345), .C(n_342771339), .D
		(n_341271326), .Z(n_57385));
	notech_and4 i_90936719(.A(n_340871322), .B(n_340671320), .C(n_317571148)
		, .D(n_317871151), .Z(n_341071324));
	notech_ao4 i_90436723(.A(n_5758), .B(n_311871099), .C(n_33194), .D(n_311771098
		), .Z(n_340871322));
	notech_ao4 i_90736721(.A(n_30326), .B(n_33322), .C(n_311471096), .D(n_31506
		), .Z(n_340671320));
	notech_and4 i_91436714(.A(n_340371317), .B(n_340171315), .C(n_318371154)
		, .D(n_318671157), .Z(n_340571319));
	notech_ao4 i_91036718(.A(n_319071161), .B(nbus_11271[30]), .C(n_310671088
		), .D(\nbus_11290[30] ), .Z(n_340371317));
	notech_ao4 i_91236716(.A(n_318871159), .B(n_33323), .C(n_318771158), .D(n_311271094
		), .Z(n_340171315));
	notech_ao4 i_104136602(.A(n_19655), .B(n_60453), .C(n_61845), .D(n_312571104
		), .Z(n_339871312));
	notech_ao4 i_104336600(.A(n_59099), .B(n_31929), .C(n_57103), .D(n_31602
		), .Z(n_3395));
	notech_ao4 i_104436599(.A(n_57122), .B(n_31801), .C(n_57616), .D(n_33320
		), .Z(n_339471310));
	notech_and2 i_105036595(.A(n_3392), .B(n_3391), .Z(n_3393));
	notech_ao4 i_104636597(.A(n_57141), .B(n_31769), .C(n_57157), .D(n_33319
		), .Z(n_3392));
	notech_ao4 i_104736596(.A(n_57168), .B(n_31865), .C(n_30590), .D(n_32026
		), .Z(n_3391));
	notech_and4 i_105836588(.A(n_3388), .B(n_3387), .C(n_338571309), .D(n_3384
		), .Z(n_3390));
	notech_ao4 i_105236594(.A(n_57192), .B(n_31737), .C(n_57062), .D(n_31705
		), .Z(n_3388));
	notech_ao4 i_105336593(.A(n_30473), .B(n_31833), .C(n_57091), .D(n_31897
		), .Z(n_3387));
	notech_ao4 i_105536591(.A(n_57218), .B(n_31438), .C(n_57230), .D(n_31673
		), .Z(n_338571309));
	notech_ao4 i_105636590(.A(n_30679), .B(n_31962), .C(n_58701), .D(n_31994
		), .Z(n_3384));
	notech_and2 i_108136568(.A(instrc[119]), .B(instrc[118]), .Z(n_3382));
	notech_and4 i_110136548(.A(n_3373), .B(n_61099), .C(n_3377), .D(n_348571371
		), .Z(n_3381));
	notech_and3 i_109436555(.A(n_58832), .B(n_57678), .C(n_57717), .Z(n_3377
		));
	notech_and4 i_110036549(.A(n_57681), .B(n_2130), .C(n_3372), .D(n_57688)
		, .Z(n_3373));
	notech_ao3 i_109736552(.A(n_56603), .B(n_50148), .C(n_10054), .Z(n_3372)
		);
	notech_ao4 i_112036532(.A(n_57336), .B(n_317171144), .C(n_316971142), .D
		(n_30345), .Z(n_3368));
	notech_and4 i_112636526(.A(nbus_11271[29]), .B(nbus_11271[30]), .C(nbus_11271
		[31]), .D(n_336071306), .Z(n_336671308));
	notech_and3 i_112536527(.A(nbus_11271[26]), .B(nbus_11271[27]), .C(nbus_11271
		[28]), .Z(n_336071306));
	notech_and4 i_113136521(.A(nbus_11271[20]), .B(nbus_11271[21]), .C(nbus_11271
		[22]), .D(n_335771304), .Z(n_335871305));
	notech_and3 i_112836524(.A(nbus_11271[23]), .B(nbus_11271[24]), .C(nbus_11271
		[25]), .Z(n_335771304));
	notech_and4 i_113736515(.A(nbus_11271[17]), .B(nbus_11271[18]), .C(nbus_11271
		[19]), .D(n_3349), .Z(n_335271300));
	notech_and3 i_113636516(.A(nbus_11271[14]), .B(nbus_11271[15]), .C(nbus_11271
		[16]), .Z(n_3349));
	notech_and4 i_114236510(.A(nbus_11271[11]), .B(nbus_11271[12]), .C(nbus_11271
		[13]), .D(n_334271294), .Z(n_334771297));
	notech_ao3 i_114136511(.A(nbus_11271[8]), .B(nbus_11271[10]), .C(opc[9])
		, .Z(n_334271294));
	notech_xor2 i_115236502(.A(n_59558), .B(opc[3]), .Z(n_333271287));
	notech_ao4 i_73837520(.A(n_2091), .B(n_57105), .C(n_19603), .D(n_2081), 
		.Z(n_3326));
	notech_ao3 i_110636544(.A(n_331471271), .B(n_331071267), .C(n_331771274)
		, .Z(n_331971276));
	notech_nand3 i_79837514(.A(n_53429), .B(n_2025), .C(n_323671201), .Z(n_331771274
		));
	notech_ao4 i_73537522(.A(n_61845), .B(n_59515), .C(n_331271269), .D(n_2081
		), .Z(n_331471271));
	notech_or4 i_195837454(.A(n_19637), .B(n_19645), .C(n_30358), .D(n_19629
		), .Z(n_331271269));
	notech_ao3 i_110436545(.A(n_2018), .B(n_2036), .C(n_2019), .Z(n_331071267
		));
	notech_and4 i_117436481(.A(n_349171376), .B(n_1847), .C(n_348071366), .D
		(n_56794), .Z(n_330471261));
	notech_and4 i_111236539(.A(n_329971256), .B(n_322671191), .C(n_325071215
		), .D(n_322271188), .Z(n_330171258));
	notech_ao4 i_110836543(.A(n_61845), .B(n_313971115), .C(n_2152), .D(n_313771114
		), .Z(n_329971256));
	notech_and3 i_117936476(.A(n_2033), .B(n_348271368), .C(n_2111), .Z(n_329871255
		));
	notech_nand2 i_118236473(.A(n_32646), .B(n_63212389), .Z(n_329671253));
	notech_or2 i_118336472(.A(n_32663), .B(n_2952), .Z(n_329571252));
	notech_and4 i_120036456(.A(n_328971246), .B(n_328671243), .C(n_328271239
		), .D(n_327671236), .Z(n_329171248));
	notech_and4 i_118736468(.A(\nbus_11290[30] ), .B(\nbus_11290[31] ), .C(\nbus_11290[11] 
		), .D(\nbus_11290[13] ), .Z(n_328971246));
	notech_and4 i_119036465(.A(\nbus_11290[0] ), .B(\nbus_11290[29] ), .C(\nbus_11290[27] 
		), .D(\nbus_11290[28] ), .Z(n_328671243));
	notech_and4 i_119536461(.A(\nbus_11290[25] ), .B(\nbus_11290[26] ), .C(\nbus_11290[23] 
		), .D(\nbus_11290[24] ), .Z(n_328271239));
	notech_and4 i_119836458(.A(\nbus_11290[21] ), .B(\nbus_11290[22] ), .C(\nbus_11290[19] 
		), .D(\nbus_11290[20] ), .Z(n_327671236));
	notech_and4 i_120336453(.A(\nbus_11290[17] ), .B(\nbus_11290[18] ), .C(\nbus_11290[15] 
		), .D(\nbus_11290[16] ), .Z(n_326871231));
	notech_and4 i_120836450(.A(\nbus_11290[12] ), .B(\nbus_11290[14] ), .C(\nbus_11290[9] 
		), .D(\nbus_11290[10] ), .Z(n_326571228));
	notech_and4 i_121636442(.A(\nbus_11290[5] ), .B(\nbus_11290[6] ), .C(n_325971223
		), .D(n_325771221), .Z(n_326271225));
	notech_and2 i_121036448(.A(\nbus_11290[7] ), .B(\nbus_11290[8] ), .Z(n_325971223
		));
	notech_and4 i_121536443(.A(\nbus_11290[3] ), .B(\nbus_11290[4] ), .C(\nbus_11290[1] 
		), .D(\nbus_11290[2] ), .Z(n_325771221));
	notech_ao4 i_122087524(.A(n_314271118), .B(n_49651676), .C(n_32575), .D(n_349271377
		), .Z(n_325471218));
	notech_mux2 i_122187523(.S(nZF), .A(n_32391), .B(n_32628), .Z(n_325371217
		));
	notech_ao4 i_111036541(.A(n_313571112), .B(n_2091), .C(n_324971214), .D(n_30346
		), .Z(n_325071215));
	notech_or4 i_122436439(.A(n_348471370), .B(n_59560), .C(n_2091), .D(n_19548
		), .Z(n_324971214));
	notech_or4 i_208637441(.A(n_19637), .B(n_19645), .C(n_19620), .D(n_19629
		), .Z(n_324671211));
	notech_or2 i_52837039(.A(n_2112), .B(n_314571121), .Z(n_324171206));
	notech_or4 i_52737040(.A(n_314960777), .B(n_32627), .C(n_60157), .D(n_314471120
		), .Z(n_324071205));
	notech_or4 i_52537041(.A(n_49651676), .B(n_32628), .C(n_60194), .D(n_57385
		), .Z(n_323971204));
	notech_or4 i_53637033(.A(n_61889), .B(n_315071126), .C(n_61723), .D(n_61870
		), .Z(n_323871203));
	notech_or4 i_53537034(.A(n_301560644), .B(n_301760646), .C(n_324671211),
		 .D(n_2081), .Z(n_323771202));
	notech_or4 i_53937030(.A(n_32484), .B(n_30343), .C(n_61684), .D(n_30618)
		, .Z(n_323671201));
	notech_nor2 i_55837013(.A(n_50409), .B(opc[4]), .Z(n_323571200));
	notech_and2 i_56637012(.A(opc[4]), .B(n_50409), .Z(n_323271197));
	notech_ao4 i_55237019(.A(n_1839), .B(n_57206), .C(n_30342), .D(n_317271145
		), .Z(n_323171196));
	notech_nao3 i_55137020(.A(n_316671139), .B(n_30425), .C(opa[0]), .Z(n_323071195
		));
	notech_nor2 i_57137011(.A(readio_ack), .B(writeio_ack), .Z(n_322771192)
		);
	notech_or4 i_51337052(.A(n_61845), .B(n_313671113), .C(\opcode[1] ), .D(\opcode[2] 
		), .Z(n_322671191));
	notech_or2 i_51637049(.A(n_32484), .B(n_309271075), .Z(n_322271188));
	notech_nao3 i_49437067(.A(n_61959), .B(n_63780), .C(n_58274), .Z(n_321971185
		));
	notech_or2 i_102337772(.A(n_311171093), .B(n_32304), .Z(n_321871184));
	notech_and4 i_15853(.A(n_32310), .B(n_61099), .C(n_32321), .D(n_32311), 
		.Z(n_321371181));
	notech_or2 i_50037779(.A(n_32292), .B(n_57103), .Z(n_321271180));
	notech_nao3 i_27115(.A(n_58274), .B(n_63780), .C(n_310571087), .Z(n_319071161
		));
	notech_nao3 i_27204(.A(n_19655), .B(n_30524), .C(n_57012), .Z(n_318971160
		));
	notech_or4 i_27206(.A(n_61845), .B(\opcode[1] ), .C(\opcode[2] ), .D(n_30305
		), .Z(n_318871159));
	notech_nand2 i_27222(.A(opc_10[30]), .B(n_63780), .Z(n_318771158));
	notech_nao3 i_38337172(.A(n_19655), .B(read_data[30]), .C(n_60453), .Z(n_318671157
		));
	notech_or2 i_38637169(.A(n_309971082), .B(\nbus_11283[30] ), .Z(n_318371154
		));
	notech_or2 i_38937166(.A(n_5750), .B(n_311571097), .Z(n_317871151));
	notech_nand2 i_39237163(.A(sav_epc[30]), .B(n_61871), .Z(n_317571148));
	notech_ao3 i_55537016(.A(rep_en5), .B(\nbus_11283[31] ), .C(n_56661), .Z
		(n_317271145));
	notech_and4 i_15037350(.A(n_336671308), .B(n_335871305), .C(n_335271300)
		, .D(n_334771297), .Z(n_317171144));
	notech_or4 i_14837352(.A(opc[6]), .B(opc[7]), .C(opc[5]), .D(n_316871141
		), .Z(n_317071143));
	notech_and2 i_14737353(.A(n_57336), .B(n_30937), .Z(n_316971142));
	notech_or4 i_14637354(.A(opc[3]), .B(opc[2]), .C(opc[4]), .D(n_57206), .Z
		(n_316871141));
	notech_or4 i_14937351(.A(n_317051260), .B(n_323271197), .C(n_323571200),
		 .D(n_333271287), .Z(n_316671139));
	notech_or4 i_55037021(.A(n_32575), .B(n_32391), .C(n_60175), .D(n_61845)
		, .Z(n_316571138));
	notech_or4 i_54937022(.A(n_32383), .B(n_63736), .C(n_61959), .D(n_32394)
		, .Z(n_316471137));
	notech_nao3 i_11237386(.A(n_338861016), .B(n_391464445), .C(n_30367), .Z
		(n_316371136));
	notech_nand2 i_54837023(.A(nZF), .B(n_316371136), .Z(n_316271135));
	notech_or4 i_53837031(.A(n_32576), .B(n_32184), .C(n_32383), .D(n_60157)
		, .Z(n_315271128));
	notech_or4 i_53737032(.A(n_314960777), .B(n_28008), .C(n_61841), .D(n_60157
		), .Z(n_315171127));
	notech_and4 i_19937327(.A(n_48030), .B(n_315271128), .C(n_30341), .D(n_330471261
		), .Z(n_315071126));
	notech_or2 i_53237035(.A(n_1817), .B(cond_1), .Z(n_314971125));
	notech_and4 i_10937389(.A(n_326871231), .B(n_326571228), .C(n_326271225)
		, .D(n_329171248), .Z(n_314571121));
	notech_and2 i_10837390(.A(n_59099), .B(n_38705), .Z(n_314471120));
	notech_or2 i_52337042(.A(n_349271377), .B(n_57385), .Z(n_314371119));
	notech_and2 i_10637392(.A(n_314371119), .B(n_325371217), .Z(n_314271118)
		);
	notech_and4 i_10737391(.A(n_324071205), .B(n_324171206), .C(n_329871255)
		, .D(n_323971204), .Z(n_313971115));
	notech_and2 i_10537393(.A(n_28533), .B(n_325471218), .Z(n_313771114));
	notech_ao4 i_10437394(.A(n_32575), .B(n_349271377), .C(n_49351679), .D(n_30313
		), .Z(n_313671113));
	notech_and2 i_10237396(.A(n_56755), .B(n_19655), .Z(n_313571112));
	notech_nao3 i_10337395(.A(n_61901), .B(n_32536), .C(n_61917), .Z(n_313471111
		));
	notech_and3 i_43937121(.A(n_61099), .B(n_61684), .C(n_30651), .Z(n_312671105
		));
	notech_and4 i_11337385(.A(n_32386), .B(n_3455), .C(n_1850), .D(n_3415), 
		.Z(n_312571104));
	notech_nand3 i_42237137(.A(n_310271084), .B(n_310171083), .C(n_310971091
		), .Z(n_311971100));
	notech_and3 i_114837712(.A(n_310871090), .B(n_310771089), .C(n_309671079
		), .Z(n_311871099));
	notech_and3 i_114737711(.A(n_310471086), .B(n_310371085), .C(n_309771080
		), .Z(n_311771098));
	notech_ao3 i_37937710(.A(n_321271180), .B(n_309871081), .C(n_321371181),
		 .Z(n_311571097));
	notech_ao4 i_24037708(.A(n_61841), .B(n_32181), .C(n_32308), .D(n_57103)
		, .Z(n_311471096));
	notech_nao3 i_148037486(.A(n_61099), .B(n_61625), .C(n_19734), .Z(n_311371095
		));
	notech_nand3 i_136637495(.A(n_56820), .B(n_3382), .C(n_311971100), .Z(n_311271094
		));
	notech_ao4 i_84037511(.A(n_63752), .B(n_61958), .C(n_61056), .D(n_58274)
		, .Z(n_311171093));
	notech_nao3 i_61837532(.A(n_30383), .B(n_30650), .C(n_348471370), .Z(n_311071092
		));
	notech_ao4 i_28537549(.A(n_2848), .B(n_30698), .C(n_32290), .D(n_32311),
		 .Z(n_310971091));
	notech_or2 i_15846(.A(n_310971091), .B(n_57501), .Z(n_310871090));
	notech_or2 i_150137764(.A(n_310271084), .B(n_57501), .Z(n_310771089));
	notech_or2 i_129637639(.A(n_310571087), .B(n_57501), .Z(n_310671088));
	notech_ao4 i_29337769(.A(n_57638), .B(n_2848), .C(n_32308), .D(n_32311),
		 .Z(n_310571087));
	notech_or2 i_15848(.A(n_57521), .B(n_310971091), .Z(n_310471086));
	notech_or2 i_150837762(.A(n_57521), .B(n_310271084), .Z(n_310371085));
	notech_ao4 i_28937641(.A(n_57679), .B(n_2848), .C(n_32288), .D(n_32311),
		 .Z(n_310271084));
	notech_ao4 i_29737642(.A(n_2848), .B(n_57657), .C(n_32292), .D(n_32311),
		 .Z(n_310171083));
	notech_or2 i_130237643(.A(n_310571087), .B(n_57521), .Z(n_309971082));
	notech_or2 i_50637659(.A(n_32288), .B(n_57103), .Z(n_309871081));
	notech_or2 i_147737766(.A(n_57521), .B(n_310171083), .Z(n_309771080));
	notech_or2 i_146637767(.A(n_310171083), .B(n_57501), .Z(n_309671079));
	notech_nand3 i_187640064(.A(n_315760785), .B(n_316260790), .C(n_30712), 
		.Z(n_309271075));
	notech_ao4 i_172141633(.A(n_58596), .B(n_32027), .C(n_58566), .D(n_31995
		), .Z(n_308971072));
	notech_ao4 i_172241632(.A(n_31439), .B(n_30664), .C(n_57529), .D(n_33318
		), .Z(n_308871071));
	notech_and2 i_172641628(.A(n_308671069), .B(n_308571068), .Z(n_308771070
		));
	notech_ao4 i_172441630(.A(n_57449), .B(n_31603), .C(n_57435), .D(n_31963
		), .Z(n_308671069));
	notech_ao4 i_172541629(.A(n_57417), .B(n_31930), .C(n_57407), .D(n_31898
		), .Z(n_308571068));
	notech_and4 i_173441620(.A(n_308171065), .B(n_308071064), .C(n_307871062
		), .D(n_307771061), .Z(n_308371067));
	notech_ao4 i_172841626(.A(n_57517), .B(n_31866), .C(n_58555), .D(n_31834
		), .Z(n_308171065));
	notech_ao4 i_172941625(.A(n_57506), .B(n_31802), .C(n_57494), .D(n_31770
		), .Z(n_308071064));
	notech_ao4 i_173141623(.A(n_57627), .B(n_33317), .C(n_30363), .D(n_31738
		), .Z(n_307871062));
	notech_ao4 i_173241622(.A(n_57471), .B(n_31706), .C(n_57461), .D(n_31674
		), .Z(n_307771061));
	notech_ao4 i_176341591(.A(n_58596), .B(n_32023), .C(n_58565), .D(n_31991
		), .Z(n_307471058));
	notech_ao4 i_176541590(.A(n_31435), .B(n_58574), .C(n_57529), .D(n_33278
		), .Z(n_307371057));
	notech_and2 i_177041586(.A(n_307171055), .B(n_307071054), .Z(n_307271056
		));
	notech_ao4 i_176741588(.A(n_57449), .B(n_31599), .C(n_57435), .D(n_31959
		), .Z(n_307171055));
	notech_ao4 i_176841587(.A(n_57417), .B(n_31926), .C(n_57407), .D(n_31894
		), .Z(n_307071054));
	notech_and4 i_177941578(.A(n_306671051), .B(n_306571050), .C(n_306371048
		), .D(n_306271047), .Z(n_306971053));
	notech_ao4 i_177241584(.A(n_57517), .B(n_31862), .C(n_58555), .D(n_31830
		), .Z(n_306671051));
	notech_ao4 i_177441583(.A(n_57506), .B(n_31798), .C(n_57494), .D(n_31766
		), .Z(n_306571050));
	notech_ao4 i_177641581(.A(n_57627), .B(n_33277), .C(n_57480), .D(n_31734
		), .Z(n_306371048));
	notech_ao4 i_177741580(.A(n_57471), .B(n_31702), .C(n_57461), .D(n_31670
		), .Z(n_306271047));
	notech_ao4 i_178041577(.A(n_58597), .B(n_32022), .C(n_58566), .D(n_31990
		), .Z(n_305971044));
	notech_ao4 i_178141576(.A(n_31434), .B(n_30664), .C(n_57529), .D(n_33276
		), .Z(n_305871043));
	notech_and2 i_178641572(.A(n_305671041), .B(n_305571040), .Z(n_305771042
		));
	notech_ao4 i_178441574(.A(n_57449), .B(n_31598), .C(n_57435), .D(n_31958
		), .Z(n_305671041));
	notech_ao4 i_178541573(.A(n_57417), .B(n_31925), .C(n_57407), .D(n_31893
		), .Z(n_305571040));
	notech_and4 i_179641564(.A(n_305271037), .B(n_305071036), .C(n_304871034
		), .D(n_304771033), .Z(n_305471039));
	notech_ao4 i_178941570(.A(n_57517), .B(n_31861), .C(n_58555), .D(n_31829
		), .Z(n_305271037));
	notech_ao4 i_179041569(.A(n_57506), .B(n_31797), .C(n_57494), .D(n_31765
		), .Z(n_305071036));
	notech_ao4 i_179241567(.A(n_57627), .B(n_33275), .C(n_30363), .D(n_31733
		), .Z(n_304871034));
	notech_ao4 i_179441566(.A(n_57472), .B(n_31701), .C(n_57461), .D(n_31669
		), .Z(n_304771033));
	notech_ao4 i_184641521(.A(n_58597), .B(n_32018), .C(n_58566), .D(n_31986
		), .Z(n_304471030));
	notech_ao4 i_184741520(.A(n_30664), .B(n_31430), .C(n_57529), .D(n_33283
		), .Z(n_304371029));
	notech_and2 i_185141516(.A(n_304171027), .B(n_304071026), .Z(n_304271028
		));
	notech_ao4 i_184941518(.A(n_57449), .B(n_31594), .C(n_57435), .D(n_31954
		), .Z(n_304171027));
	notech_ao4 i_185041517(.A(n_57417), .B(n_31921), .C(n_57407), .D(n_31889
		), .Z(n_304071026));
	notech_and4 i_185941508(.A(n_303771023), .B(n_303671022), .C(n_303371020
		), .D(n_303271019), .Z(n_303971025));
	notech_ao4 i_185341514(.A(n_57517), .B(n_31857), .C(n_58555), .D(n_31825
		), .Z(n_303771023));
	notech_ao4 i_185441513(.A(n_57506), .B(n_31793), .C(n_57494), .D(n_31761
		), .Z(n_303671022));
	notech_ao4 i_185641511(.A(n_57627), .B(n_33282), .C(n_30363), .D(n_31729
		), .Z(n_303371020));
	notech_ao4 i_185741510(.A(n_57472), .B(n_31697), .C(n_57461), .D(n_31665
		), .Z(n_303271019));
	notech_ao4 i_186041507(.A(n_58597), .B(n_32017), .C(n_58566), .D(n_31985
		), .Z(n_302971016));
	notech_ao4 i_186241506(.A(n_30664), .B(n_31429), .C(n_57529), .D(n_33287
		), .Z(n_302871015));
	notech_and2 i_186641502(.A(n_302671013), .B(n_302571012), .Z(n_302771014
		));
	notech_ao4 i_186441504(.A(n_57449), .B(n_31593), .C(n_57435), .D(n_31953
		), .Z(n_302671013));
	notech_ao4 i_186541503(.A(n_57417), .B(n_31920), .C(n_57407), .D(n_31888
		), .Z(n_302571012));
	notech_and4 i_187441494(.A(n_302271009), .B(n_302171008), .C(n_301971006
		), .D(n_301671005), .Z(n_302471011));
	notech_ao4 i_186841500(.A(n_57517), .B(n_31856), .C(n_58555), .D(n_31824
		), .Z(n_302271009));
	notech_ao4 i_186941499(.A(n_57506), .B(n_31792), .C(n_57494), .D(n_31760
		), .Z(n_302171008));
	notech_ao4 i_187141497(.A(n_57627), .B(n_33286), .C(n_30363), .D(n_31728
		), .Z(n_301971006));
	notech_ao4 i_187241496(.A(n_57472), .B(n_31696), .C(n_57461), .D(n_31664
		), .Z(n_301671005));
	notech_ao4 i_187541493(.A(n_58596), .B(n_32016), .C(n_58565), .D(n_31984
		), .Z(n_301271002));
	notech_ao4 i_187641492(.A(n_58574), .B(n_31428), .C(n_33291), .D(n_57529
		), .Z(n_301171001));
	notech_and2 i_188041488(.A(n_300970999), .B(n_300870998), .Z(n_301071000
		));
	notech_ao4 i_187841490(.A(n_57449), .B(n_31592), .C(n_57435), .D(n_31952
		), .Z(n_300970999));
	notech_ao4 i_187941489(.A(n_57417), .B(n_31919), .C(n_57407), .D(n_31887
		), .Z(n_300870998));
	notech_and4 i_188841480(.A(n_300570995), .B(n_300470994), .C(n_300270992
		), .D(n_300170991), .Z(n_300770997));
	notech_ao4 i_188241486(.A(n_57517), .B(n_31855), .C(n_58555), .D(n_31823
		), .Z(n_300570995));
	notech_ao4 i_188341485(.A(n_57506), .B(n_31791), .C(n_57494), .D(n_31759
		), .Z(n_300470994));
	notech_ao4 i_188541483(.A(n_57627), .B(n_33290), .C(n_57480), .D(n_31727
		), .Z(n_300270992));
	notech_ao4 i_188641482(.A(n_57471), .B(n_31695), .C(n_57461), .D(n_31663
		), .Z(n_300170991));
	notech_ao4 i_189041479(.A(n_58596), .B(n_32015), .C(n_58565), .D(n_31983
		), .Z(n_299870988));
	notech_ao4 i_189141478(.A(n_31427), .B(n_58574), .C(n_57529), .D(n_33309
		), .Z(n_299670987));
	notech_and2 i_189641474(.A(n_299470985), .B(n_299370984), .Z(n_299570986
		));
	notech_ao4 i_189341476(.A(n_57449), .B(n_31591), .C(n_57435), .D(n_31951
		), .Z(n_299470985));
	notech_ao4 i_189441475(.A(n_57417), .B(n_31918), .C(n_57406), .D(n_31886
		), .Z(n_299370984));
	notech_and4 i_190741466(.A(n_299070981), .B(n_298970980), .C(n_298770978
		), .D(n_298670977), .Z(n_299270983));
	notech_ao4 i_189841472(.A(n_57517), .B(n_31854), .C(n_58555), .D(n_31822
		), .Z(n_299070981));
	notech_ao4 i_189941471(.A(n_57506), .B(n_31790), .C(n_57494), .D(n_31758
		), .Z(n_298970980));
	notech_ao4 i_190341469(.A(n_57627), .B(n_33308), .C(n_57480), .D(n_31726
		), .Z(n_298770978));
	notech_ao4 i_190441468(.A(n_57471), .B(n_31694), .C(n_57461), .D(n_31662
		), .Z(n_298670977));
	notech_ao4 i_190841465(.A(n_58596), .B(n_32014), .C(n_58565), .D(n_31982
		), .Z(n_298370974));
	notech_ao4 i_190941464(.A(n_31426), .B(n_58574), .C(n_57529), .D(n_33307
		), .Z(n_298270973));
	notech_and2 i_191341460(.A(n_298070971), .B(n_297970970), .Z(n_298170972
		));
	notech_ao4 i_191141462(.A(n_57449), .B(n_31590), .C(n_57435), .D(n_31950
		), .Z(n_298070971));
	notech_ao4 i_191241461(.A(n_57417), .B(n_31917), .C(n_57406), .D(n_31885
		), .Z(n_297970970));
	notech_and4 i_192241452(.A(n_297670967), .B(n_297570966), .C(n_297370964
		), .D(n_297270963), .Z(n_297870969));
	notech_ao4 i_191541458(.A(n_57517), .B(n_31853), .C(n_58555), .D(n_31821
		), .Z(n_297670967));
	notech_ao4 i_191641457(.A(n_57506), .B(n_31789), .C(n_57494), .D(n_31757
		), .Z(n_297570966));
	notech_ao4 i_191941455(.A(n_57627), .B(n_33306), .C(n_57480), .D(n_31725
		), .Z(n_297370964));
	notech_ao4 i_192041454(.A(n_57471), .B(n_31693), .C(n_57461), .D(n_31661
		), .Z(n_297270963));
	notech_ao4 i_192341451(.A(n_58596), .B(n_32013), .C(n_58565), .D(n_31981
		), .Z(n_296970960));
	notech_ao4 i_192441450(.A(n_31425), .B(n_58574), .C(n_57529), .D(n_33305
		), .Z(n_296870959));
	notech_and2 i_192841446(.A(n_296670957), .B(n_296570956), .Z(n_296770958
		));
	notech_ao4 i_192641448(.A(n_57449), .B(n_31589), .C(n_57435), .D(n_31949
		), .Z(n_296670957));
	notech_ao4 i_192741447(.A(n_57417), .B(n_31916), .C(n_57406), .D(n_31884
		), .Z(n_296570956));
	notech_and4 i_193641438(.A(n_296270953), .B(n_296170952), .C(n_295970950
		), .D(n_295870949), .Z(n_296470955));
	notech_ao4 i_193041444(.A(n_57517), .B(n_31852), .C(n_58555), .D(n_31820
		), .Z(n_296270953));
	notech_ao4 i_193141443(.A(n_57506), .B(n_31788), .C(n_57494), .D(n_31756
		), .Z(n_296170952));
	notech_ao4 i_193341441(.A(n_57627), .B(n_33304), .C(n_57480), .D(n_31724
		), .Z(n_295970950));
	notech_ao4 i_193441440(.A(n_57471), .B(n_31692), .C(n_57461), .D(n_31660
		), .Z(n_295870949));
	notech_ao4 i_193741437(.A(n_58596), .B(n_32012), .C(n_58565), .D(n_31980
		), .Z(n_295570946));
	notech_ao4 i_193841436(.A(n_31424), .B(n_58574), .C(n_57529), .D(n_33303
		), .Z(n_295470945));
	notech_and2 i_194341432(.A(n_295270943), .B(n_295170942), .Z(n_295370944
		));
	notech_ao4 i_194041434(.A(n_57449), .B(n_31588), .C(n_57435), .D(n_31948
		), .Z(n_295270943));
	notech_ao4 i_194241433(.A(n_57417), .B(n_31915), .C(n_57406), .D(n_31883
		), .Z(n_295170942));
	notech_and4 i_195141424(.A(n_294870939), .B(n_294770938), .C(n_294570936
		), .D(n_294470935), .Z(n_295070941));
	notech_ao4 i_194541430(.A(n_57517), .B(n_31851), .C(n_58555), .D(n_31819
		), .Z(n_294870939));
	notech_ao4 i_194641429(.A(n_57506), .B(n_31787), .C(n_57494), .D(n_31755
		), .Z(n_294770938));
	notech_ao4 i_194841427(.A(n_57627), .B(n_33302), .C(n_57480), .D(n_31723
		), .Z(n_294570936));
	notech_ao4 i_194941426(.A(n_57471), .B(n_31691), .C(n_57461), .D(n_31659
		), .Z(n_294470935));
	notech_ao4 i_202541353(.A(n_58597), .B(n_32004), .C(n_58566), .D(n_31972
		), .Z(n_294170932));
	notech_ao4 i_202741352(.A(n_31416), .B(n_58574), .C(n_57529), .D(n_33315
		), .Z(n_294070931));
	notech_and2 i_203141348(.A(n_293870929), .B(n_293770928), .Z(n_293970930
		));
	notech_ao4 i_202941350(.A(n_57449), .B(n_31580), .C(n_57435), .D(n_31939
		), .Z(n_293870929));
	notech_ao4 i_203041349(.A(n_57417), .B(n_31907), .C(n_57406), .D(n_31875
		), .Z(n_293770928));
	notech_and4 i_203941340(.A(n_293470925), .B(n_293370924), .C(n_293170922
		), .D(n_293070921), .Z(n_293670927));
	notech_ao4 i_203341346(.A(n_57517), .B(n_31843), .C(n_58555), .D(n_31811
		), .Z(n_293470925));
	notech_ao4 i_203441345(.A(n_57506), .B(n_31779), .C(n_57494), .D(n_31747
		), .Z(n_293370924));
	notech_ao4 i_203641343(.A(n_57627), .B(n_33314), .C(n_57480), .D(n_31715
		), .Z(n_293170922));
	notech_ao4 i_203741342(.A(n_57472), .B(n_31683), .C(n_57461), .D(n_31651
		), .Z(n_293070921));
	notech_ao4 i_219041190(.A(n_32026), .B(n_58597), .C(n_58566), .D(n_31994
		), .Z(n_292670917));
	notech_ao4 i_219141189(.A(n_31438), .B(n_30664), .C(n_57529), .D(n_33319
		), .Z(n_292570916));
	notech_and2 i_219541185(.A(n_292370914), .B(n_292270913), .Z(n_292470915
		));
	notech_ao4 i_219341187(.A(n_57449), .B(n_31602), .C(n_57435), .D(n_31962
		), .Z(n_292370914));
	notech_ao4 i_219441186(.A(n_57417), .B(n_31929), .C(n_57407), .D(n_31897
		), .Z(n_292270913));
	notech_and4 i_220341177(.A(n_291970910), .B(n_291870909), .C(n_291670907
		), .D(n_291570906), .Z(n_292170912));
	notech_ao4 i_219741183(.A(n_57517), .B(n_31865), .C(n_58555), .D(n_31833
		), .Z(n_291970910));
	notech_ao4 i_219841182(.A(n_57506), .B(n_31801), .C(n_31769), .D(n_57494
		), .Z(n_291870909));
	notech_ao4 i_220041180(.A(n_57627), .B(n_33320), .C(n_30363), .D(n_31737
		), .Z(n_291670907));
	notech_ao4 i_220141179(.A(n_57472), .B(n_31705), .C(n_57461), .D(n_31673
		), .Z(n_291570906));
	notech_nand3 i_113642204(.A(opz[1]), .B(n_31606), .C(n_31604), .Z(n_272170713
		));
	notech_and4 i_175444759(.A(n_271870710), .B(n_253070525), .C(n_271670708
		), .D(n_252770522), .Z(n_272070712));
	notech_ao4 i_175044763(.A(n_318871159), .B(n_33310), .C(n_309771080), .D
		(n_33169), .Z(n_271870710));
	notech_or4 i_76768524(.A(n_379164322), .B(n_324660874), .C(n_33173), .D(n_30733
		), .Z(n_134672731));
	notech_or2 i_77468517(.A(n_54741988), .B(n_31480), .Z(n_135372738));
	notech_nand3 i_820966(.A(n_137972764), .B(n_137072755), .C(n_137872763),
		 .Z(n_18914));
	notech_nao3 i_79168500(.A(n_63752), .B(opc_10[6]), .C(n_376664297), .Z(n_135872743
		));
	notech_or2 i_79868493(.A(n_54741988), .B(n_31479), .Z(n_136572750));
	notech_nand3 i_720965(.A(n_139072775), .B(n_138172766), .C(n_138972774),
		 .Z(n_18908));
	notech_ao4 i_78868503(.A(n_29681), .B(n_324760875), .C(n_29680), .D(n_324260870
		), .Z(n_137072755));
	notech_ao4 i_78068511(.A(n_376564296), .B(n_324160869), .C(n_376764298),
		 .D(n_324560873), .Z(n_137172756));
	notech_ao4 i_78168510(.A(n_376864299), .B(n_100242443), .C(n_94542386), 
		.D(n_324060868), .Z(n_137272757));
	notech_ao4 i_78268509(.A(n_323760865), .B(n_57136), .C(n_376964300), .D(n_33165
		), .Z(n_137472759));
	notech_and3 i_78368508(.A(n_324860876), .B(n_134672731), .C(n_135372738)
		, .Z(n_137672761));
	notech_and4 i_78668505(.A(n_137472759), .B(n_137272757), .C(n_137172756)
		, .D(n_137672761), .Z(n_137872763));
	notech_ao4 i_78768504(.A(n_29678), .B(n_324460872), .C(n_324360871), .D(n_29677
		), .Z(n_137972764));
	notech_ao4 i_81368479(.A(n_29681), .B(n_325460882), .C(n_29680), .D(n_325660884
		), .Z(n_138172766));
	notech_ao4 i_80468487(.A(n_324960877), .B(n_376564296), .C(n_325360881),
		 .D(n_376764298), .Z(n_138272767));
	notech_ao4 i_80568486(.A(n_100542446), .B(n_376864299), .C(n_94542386), 
		.D(n_325160879), .Z(n_138372768));
	notech_ao4 i_80668485(.A(n_57136), .B(n_325060878), .C(n_376964300), .D(n_33166
		), .Z(n_138572770));
	notech_and3 i_80768484(.A(n_135872743), .B(n_325860886), .C(n_136572750)
		, .Z(n_138772772));
	notech_and4 i_81068481(.A(n_138572770), .B(n_138372768), .C(n_138272767)
		, .D(n_138772772), .Z(n_138972774));
	notech_ao4 i_81168480(.A(n_325760885), .B(n_29678), .C(n_325560883), .D(n_29677
		), .Z(n_139072775));
	notech_or2 i_15566002(.A(n_31071), .B(n_26275), .Z(n_139972784));
	notech_or2 i_15066007(.A(n_334660974), .B(n_332460952), .Z(n_140472789)
		);
	notech_ao3 i_14566012(.A(n_19612), .B(read_data[4]), .C(n_35412112), .Z(n_140972794
		));
	notech_or2 i_17365984(.A(n_31122), .B(n_26275), .Z(n_141772802));
	notech_or2 i_16865989(.A(n_334860976), .B(n_332460952), .Z(n_142272807)
		);
	notech_ao3 i_16365994(.A(n_19612), .B(read_data[5]), .C(n_35412112), .Z(n_142772812
		));
	notech_ao4 i_113565044(.A(n_331160939), .B(\nbus_11290[5] ), .C(n_61099)
		, .D(n_30782), .Z(n_142872813));
	notech_ao4 i_113465045(.A(n_334960977), .B(n_26603), .C(n_331460942), .D
		(n_31478), .Z(n_143072815));
	notech_ao3 i_113765042(.A(n_142872813), .B(n_143072815), .C(n_142772812)
		, .Z(n_143172816));
	notech_ao4 i_113165048(.A(n_332260950), .B(n_33135), .C(n_31098), .D(n_332160949
		), .Z(n_143272817));
	notech_ao4 i_113065049(.A(n_31118), .B(n_26268), .C(n_31099), .D(n_26278
		), .Z(n_143472819));
	notech_and4 i_113865041(.A(n_143272817), .B(n_143472819), .C(n_142272807
		), .D(n_143172816), .Z(n_143672821));
	notech_ao4 i_112465053(.A(n_31125), .B(n_26277), .C(n_31119), .D(n_26271
		), .Z(n_143772822));
	notech_ao4 i_112365054(.A(n_31126), .B(n_26272), .C(n_31123), .D(n_26276
		), .Z(n_143972824));
	notech_and3 i_112865051(.A(n_143772822), .B(n_143972824), .C(n_141772802
		), .Z(n_144072825));
	notech_ao4 i_112165056(.A(n_126126588), .B(n_32064), .C(n_125926586), .D
		(n_33327), .Z(n_144172826));
	notech_ao4 i_112065057(.A(n_28240), .B(nbus_11273[5]), .C(n_26585), .D(n_30977
		), .Z(n_144272827));
	notech_ao4 i_111665061(.A(n_331160939), .B(\nbus_11290[4] ), .C(n_61099)
		, .D(n_30781), .Z(n_144572830));
	notech_ao4 i_111565062(.A(n_334760975), .B(n_26603), .C(n_331460942), .D
		(n_31477), .Z(n_144772832));
	notech_ao3 i_111865059(.A(n_144572830), .B(n_144772832), .C(n_140972794)
		, .Z(n_144872833));
	notech_ao4 i_111265065(.A(n_332260950), .B(n_33104), .C(n_31047), .D(n_332160949
		), .Z(n_144972834));
	notech_ao4 i_111165066(.A(n_31067), .B(n_26268), .C(n_31048), .D(n_26278
		), .Z(n_145172836));
	notech_and4 i_111965058(.A(n_144972834), .B(n_145172836), .C(n_140472789
		), .D(n_144872833), .Z(n_145372838));
	notech_ao4 i_110765070(.A(n_31074), .B(n_26277), .C(n_31068), .D(n_26271
		), .Z(n_145472839));
	notech_ao4 i_110665071(.A(n_31075), .B(n_26272), .C(n_31072), .D(n_26276
		), .Z(n_145672841));
	notech_and3 i_110965068(.A(n_145472839), .B(n_145672841), .C(n_139972784
		), .Z(n_145772842));
	notech_ao4 i_110065073(.A(n_126126588), .B(n_32063), .C(n_125926586), .D
		(n_33326), .Z(n_145872843));
	notech_ao4 i_109965074(.A(n_28240), .B(nbus_11273[4]), .C(n_26585), .D(n_30975
		), .Z(n_145972844));
	notech_nor2 i_54252538(.A(n_363450925), .B(n_442968013), .Z(n_146672851)
		);
	notech_ao3 i_54352537(.A(n_63752), .B(opc_10[23]), .C(n_442768011), .Z(n_147372858
		));
	notech_or4 i_2420758(.A(n_77826105), .B(n_185473225), .C(n_147372858), .D
		(n_146672851), .Z(n_19706));
	notech_nor2 i_58952492(.A(n_3466), .B(n_442968013), .Z(n_147872863));
	notech_ao3 i_59052491(.A(opc_10[21]), .B(n_63754), .C(n_442768011), .Z(n_148572870
		));
	notech_or4 i_2220756(.A(n_75626083), .B(n_186773235), .C(n_148572870), .D
		(n_147872863), .Z(n_19694));
	notech_or4 i_61252469(.A(n_339561023), .B(n_2829), .C(n_444168025), .D(n_346771358
		), .Z(n_149072875));
	notech_nao3 i_61352468(.A(opc_10[20]), .B(n_63736), .C(n_442768011), .Z(n_149772882
		));
	notech_nand3 i_2120755(.A(n_187873246), .B(n_149772882), .C(n_149072875)
		, .Z(n_19688));
	notech_nor2 i_64452437(.A(n_363450925), .B(n_443468018), .Z(n_149872883)
		);
	notech_ao3 i_64552436(.A(n_63752), .B(opc_10[23]), .C(n_443568019), .Z(n_150572890
		));
	notech_or4 i_2420854(.A(n_77826105), .B(n_188473252), .C(n_150572890), .D
		(n_149872883), .Z(n_19358));
	notech_or4 i_66052421(.A(n_32217), .B(n_2829), .C(n_57256), .D(n_3464), 
		.Z(n_150672891));
	notech_nao3 i_66152420(.A(opc_10[22]), .B(n_63736), .C(n_443568019), .Z(n_151372898
		));
	notech_nand3 i_2320853(.A(n_189273260), .B(n_150672891), .C(n_151372898)
		, .Z(n_19352));
	notech_nor2 i_67652405(.A(n_3466), .B(n_443468018), .Z(n_151472899));
	notech_ao3 i_67752404(.A(opc_10[21]), .B(n_63736), .C(n_443568019), .Z(n_152172906
		));
	notech_or4 i_2220852(.A(n_75626083), .B(n_189873266), .C(n_152172906), .D
		(n_151472899), .Z(n_19346));
	notech_or4 i_69252389(.A(n_2829), .B(n_444168025), .C(n_346771358), .D(n_32217
		), .Z(n_152272907));
	notech_nao3 i_69352388(.A(opc_10[20]), .B(n_63736), .C(n_443568019), .Z(n_152972914
		));
	notech_nand3 i_2120851(.A(n_190673274), .B(n_152272907), .C(n_152972914)
		, .Z(n_19340));
	notech_nor2 i_74052341(.A(n_363450925), .B(n_443968023), .Z(n_153072915)
		);
	notech_ao3 i_74152340(.A(n_63752), .B(opc_10[23]), .C(n_444068024), .Z(n_153772922
		));
	notech_or4 i_2420982(.A(n_77826105), .B(n_191273280), .C(n_153772922), .D
		(n_153072915), .Z(n_19010));
	notech_nor2 i_77252309(.A(n_3466), .B(n_443968023), .Z(n_153872923));
	notech_ao3 i_77352308(.A(opc_10[21]), .B(n_63736), .C(n_444068024), .Z(n_154572930
		));
	notech_or4 i_2220980(.A(n_75626083), .B(n_191973287), .C(n_154572930), .D
		(n_153872923), .Z(n_18998));
	notech_or4 i_79052293(.A(n_339561023), .B(n_444168025), .C(n_346771358),
		 .D(n_340461032), .Z(n_154672931));
	notech_nao3 i_79152292(.A(opc_10[20]), .B(n_63782), .C(n_444068024), .Z(n_155372938
		));
	notech_nand3 i_2120979(.A(n_192773295), .B(n_154672931), .C(n_155372938)
		, .Z(n_18992));
	notech_or4 i_84052245(.A(n_340461032), .B(n_32217), .C(n_444168025), .D(n_363450925
		), .Z(n_155472939));
	notech_nao3 i_84152244(.A(n_63752), .B(opc_10[23]), .C(n_299122016), .Z(n_156172946
		));
	notech_nand3 i_2421014(.A(n_193473302), .B(n_156172946), .C(n_155472939)
		, .Z(n_18662));
	notech_or4 i_87252213(.A(n_340461032), .B(n_32217), .C(n_57256), .D(n_3466
		), .Z(n_156272947));
	notech_nao3 i_87352212(.A(opc_10[21]), .B(n_63736), .C(n_299122016), .Z(n_156972954
		));
	notech_nand3 i_2221012(.A(n_194173309), .B(n_156972954), .C(n_156272947)
		, .Z(n_18650));
	notech_or2 i_88852197(.A(n_346771358), .B(n_303822063), .Z(n_157072955)
		);
	notech_nao3 i_88952196(.A(opc_10[20]), .B(n_63736), .C(n_299122016), .Z(n_157772962
		));
	notech_nand3 i_2121011(.A(n_194873316), .B(n_157772962), .C(n_157072955)
		, .Z(n_18644));
	notech_nor2 i_93652149(.A(n_363450925), .B(n_325325323), .Z(n_157872963)
		);
	notech_ao3 i_93752148(.A(n_63776), .B(opc_10[23]), .C(n_315725234), .Z(n_158572970
		));
	notech_or4 i_2421078(.A(n_77826105), .B(n_195473322), .C(n_158572970), .D
		(n_157872963), .Z(n_16361));
	notech_nor2 i_96852117(.A(n_3466), .B(n_325325323), .Z(n_158672971));
	notech_ao3 i_96952116(.A(opc_10[21]), .B(n_63736), .C(n_315725234), .Z(n_159372978
		));
	notech_or4 i_2221076(.A(n_75626083), .B(n_196173329), .C(n_159372978), .D
		(n_158672971), .Z(n_16349));
	notech_or4 i_98452101(.A(n_340361031), .B(n_57256), .C(n_346771358), .D(n_339561023
		), .Z(n_159472979));
	notech_nao3 i_98552100(.A(opc_10[20]), .B(n_63736), .C(n_315725234), .Z(n_160172986
		));
	notech_nand3 i_2121075(.A(n_196973337), .B(n_159472979), .C(n_160172986)
		, .Z(n_16343));
	notech_nor2 i_117251916(.A(n_3464), .B(n_122226549), .Z(n_160272987));
	notech_ao3 i_117351915(.A(opc_10[22]), .B(n_63736), .C(n_337461002), .Z(n_161372998
		));
	notech_or4 i_2321333(.A(n_161372998), .B(n_197873346), .C(n_197373341), 
		.D(n_160272987), .Z(n_16006));
	notech_nor2 i_119751893(.A(n_3466), .B(n_122226549), .Z(n_161472999));
	notech_ao3 i_119851892(.A(opc_10[21]), .B(n_63736), .C(n_337461002), .Z(n_162573010
		));
	notech_or4 i_2221332(.A(n_162573010), .B(n_198873356), .C(n_198373351), 
		.D(n_161472999), .Z(n_16000));
	notech_nor2 i_122051870(.A(n_346771358), .B(n_122226549), .Z(n_162673011
		));
	notech_ao3 i_122151869(.A(opc_10[20]), .B(n_63736), .C(n_337461002), .Z(n_163773022
		));
	notech_or4 i_2121331(.A(n_163773022), .B(n_199873366), .C(n_199373361), 
		.D(n_162673011), .Z(n_15994));
	notech_nor2 i_134551745(.A(n_124126568), .B(n_363350926), .Z(n_163873023
		));
	notech_ao3 i_134651744(.A(n_63776), .B(opc_10[25]), .C(n_337661004), .Z(n_164973034
		));
	notech_or4 i_2621528(.A(n_164973034), .B(n_200873376), .C(n_200373371), 
		.D(n_163873023), .Z(n_15672));
	notech_nor2 i_139151699(.A(n_363450925), .B(n_124126568), .Z(n_165073035
		));
	notech_ao3 i_139251698(.A(n_63776), .B(opc_10[23]), .C(n_337661004), .Z(n_166173046
		));
	notech_or4 i_2421526(.A(n_166173046), .B(n_201873386), .C(n_201373381), 
		.D(n_165073035), .Z(n_15660));
	notech_nor2 i_141451676(.A(n_3464), .B(n_124126568), .Z(n_166273047));
	notech_ao3 i_141551675(.A(opc_10[22]), .B(n_63736), .C(n_337661004), .Z(n_167273057
		));
	notech_or4 i_2321525(.A(n_167273057), .B(n_202873396), .C(n_202373391), 
		.D(n_166273047), .Z(n_15654));
	notech_nor2 i_143751653(.A(n_3466), .B(n_124126568), .Z(n_167373058));
	notech_ao3 i_143851652(.A(opc_10[21]), .B(n_63736), .C(n_337661004), .Z(n_168373068
		));
	notech_or4 i_2221524(.A(n_168373068), .B(n_203873406), .C(n_203373401), 
		.D(n_167373058), .Z(n_15648));
	notech_nor2 i_146051630(.A(n_346771358), .B(n_124126568), .Z(n_168473069
		));
	notech_ao3 i_146151629(.A(opc_10[20]), .B(n_63736), .C(n_337661004), .Z(n_169473079
		));
	notech_or4 i_2121523(.A(n_169473079), .B(n_204873416), .C(n_204373411), 
		.D(n_168473069), .Z(n_15642));
	notech_nor2 i_151151579(.A(n_363450925), .B(n_387664407), .Z(n_169573080
		));
	notech_ao3 i_151251578(.A(n_63776), .B(opc_10[23]), .C(n_387764408), .Z(n_170273087
		));
	notech_or4 i_2421622(.A(n_77826105), .B(n_205573423), .C(n_170273087), .D
		(n_169573080), .Z(n_13130));
	notech_nor2 i_154351547(.A(n_3466), .B(n_387664407), .Z(n_170373088));
	notech_ao3 i_154451546(.A(opc_10[21]), .B(n_63782), .C(n_387764408), .Z(n_171073095
		));
	notech_or4 i_2221620(.A(n_75626083), .B(n_206273430), .C(n_171073095), .D
		(n_170373088), .Z(n_13118));
	notech_or4 i_155951531(.A(n_57256), .B(n_346771358), .C(n_2829), .D(n_2845
		), .Z(n_171173096));
	notech_ao3 i_156051530(.A(opc_10[20]), .B(n_63756), .C(n_387764408), .Z(n_171873103
		));
	notech_nao3 i_2121619(.A(n_207073438), .B(n_171173096), .C(n_171873103),
		 .Z(n_13112));
	notech_or2 i_163051460(.A(n_363450925), .B(n_126226589), .Z(n_171973104)
		);
	notech_nand2 i_162951461(.A(sav_esp[23]), .B(n_61870), .Z(n_173073115)
		);
	notech_nao3 i_163151459(.A(n_63776), .B(opc_10[23]), .C(n_337961007), .Z
		(n_173173116));
	notech_nand3 i_2421782(.A(n_173173116), .B(n_208173449), .C(n_171973104)
		, .Z(n_15308));
	notech_or2 i_165551435(.A(n_126226589), .B(n_3464), .Z(n_173273117));
	notech_nand2 i_165451436(.A(sav_esp[22]), .B(n_61871), .Z(n_174373128)
		);
	notech_nao3 i_165651434(.A(opc_10[22]), .B(n_63764), .C(n_337961007), .Z
		(n_174473129));
	notech_nand3 i_2321781(.A(n_174473129), .B(n_209273460), .C(n_173273117)
		, .Z(n_15302));
	notech_or2 i_168051410(.A(n_3466), .B(n_126226589), .Z(n_174573130));
	notech_nand2 i_167951411(.A(sav_esp[21]), .B(n_61871), .Z(n_176273141)
		);
	notech_nao3 i_168151409(.A(opc_10[21]), .B(n_63764), .C(n_337961007), .Z
		(n_176373142));
	notech_nand3 i_2221780(.A(n_176373142), .B(n_210373471), .C(n_174573130)
		, .Z(n_15296));
	notech_or2 i_170551385(.A(n_346771358), .B(n_126226589), .Z(n_176473143)
		);
	notech_nand2 i_170451386(.A(sav_esp[20]), .B(n_61870), .Z(n_177573154)
		);
	notech_nao3 i_170651384(.A(opc_10[20]), .B(n_63764), .C(n_337961007), .Z
		(n_177673155));
	notech_nand3 i_2121779(.A(n_177673155), .B(n_211473482), .C(n_176473143)
		, .Z(n_15290));
	notech_nor2 i_175851332(.A(n_363450925), .B(n_301522040), .Z(n_177773156
		));
	notech_ao3 i_175951331(.A(n_63776), .B(opc_10[23]), .C(n_298922014), .Z(n_178473163
		));
	notech_or4 i_2421846(.A(n_77826105), .B(n_212073488), .C(n_178473163), .D
		(n_177773156), .Z(n_12782));
	notech_nor2 i_179251299(.A(n_3466), .B(n_301522040), .Z(n_178573164));
	notech_nand3 i_179151300(.A(n_57392), .B(n_32210), .C(opd[21]), .Z(n_179173170
		));
	notech_ao3 i_179351298(.A(opc_10[21]), .B(n_63782), .C(n_298922014), .Z(n_179273171
		));
	notech_or4 i_2221844(.A(n_75626083), .B(n_179273171), .C(n_178573164), .D
		(n_30285), .Z(n_12770));
	notech_or2 i_181051282(.A(n_346771358), .B(n_301522040), .Z(n_179373172)
		);
	notech_nao3 i_181151281(.A(opc_10[20]), .B(n_63782), .C(n_298922014), .Z
		(n_180073179));
	notech_nand3 i_2121843(.A(n_213673504), .B(n_180073179), .C(n_179373172)
		, .Z(n_12764));
	notech_or4 i_186651227(.A(n_340461032), .B(n_2830), .C(n_57256), .D(n_363450925
		), .Z(n_180173180));
	notech_nand2 i_3553039(.A(n_61625), .B(read_data[23]), .Z(n_180473183)
		);
	notech_or2 i_186551228(.A(n_25110), .B(nbus_11271[23]), .Z(n_180573184)
		);
	notech_or2 i_186051233(.A(n_365628696), .B(\nbus_11283[23] ), .Z(n_180673185
		));
	notech_or2 i_186351230(.A(n_365228692), .B(n_33170), .Z(n_180973188));
	notech_nao3 i_186451229(.A(n_63748), .B(opc_10[23]), .C(n_365428694), .Z
		(n_181073189));
	notech_nand3 i_2421910(.A(n_181073189), .B(n_214473512), .C(n_180173180)
		, .Z(n_12430));
	notech_or4 i_190351190(.A(n_340461032), .B(n_2830), .C(n_57256), .D(n_3466
		), .Z(n_181173190));
	notech_nand2 i_189551198(.A(tsc[53]), .B(n_30615), .Z(n_181273191));
	notech_nand2 i_3753037(.A(n_61625), .B(read_data[21]), .Z(n_181373192)
		);
	notech_or2 i_190251191(.A(n_25110), .B(nbus_11271[21]), .Z(n_181573194)
		);
	notech_or2 i_189751196(.A(n_365628696), .B(\nbus_11283[21] ), .Z(n_181673195
		));
	notech_or2 i_190051193(.A(n_365228692), .B(n_33288), .Z(n_181973198));
	notech_nao3 i_190151192(.A(opc_10[21]), .B(n_63764), .C(n_365428694), .Z
		(n_182173199));
	notech_nand3 i_2221908(.A(n_215373521), .B(n_182173199), .C(n_181173190)
		, .Z(n_12418));
	notech_nor2 i_208651008(.A(n_388064411), .B(n_363450925), .Z(n_182273200
		));
	notech_nao3 i_208551009(.A(n_57392), .B(opd[23]), .C(n_58701), .Z(n_183573207
		));
	notech_ao3 i_208751007(.A(n_63748), .B(opc_10[23]), .C(n_388164412), .Z(n_183673208
		));
	notech_or4 i_2417590(.A(n_77826105), .B(n_183673208), .C(n_182273200), .D
		(n_30284), .Z(n_11704));
	notech_or4 i_214050954(.A(n_444168025), .B(n_346771358), .C(n_340361031)
		, .D(n_2830), .Z(n_183773209));
	notech_nao3 i_213950955(.A(n_57392), .B(opd[20]), .C(n_58701), .Z(n_184573216
		));
	notech_nao3 i_214150953(.A(opc_10[20]), .B(n_63782), .C(n_388164412), .Z
		(n_184673217));
	notech_and4 i_2117587(.A(n_216873536), .B(n_183773209), .C(n_74526072), 
		.D(n_184673217), .Z(n_11686));
	notech_ao4 i_53452546(.A(n_30697), .B(n_33170), .C(n_30689), .D(n_109226419
		), .Z(n_184773218));
	notech_ao4 i_53352547(.A(n_30693), .B(\nbus_11290[23] ), .C(n_30695), .D
		(\nbus_11283[23] ), .Z(n_184873219));
	notech_nand3 i_51553072(.A(n_180473183), .B(n_184873219), .C(n_184773218
		), .Z(n_77826105));
	notech_ao4 i_54652534(.A(n_327960907), .B(n_31499), .C(n_117626503), .D(n_33170
		), .Z(n_185073221));
	notech_ao4 i_54452536(.A(n_442668010), .B(\nbus_11283[23] ), .C(n_442868012
		), .D(nbus_11271[23]), .Z(n_185173222));
	notech_ao4 i_54552535(.A(n_109226419), .B(n_117726504), .C(n_442568009),
		 .D(\nbus_11290[23] ), .Z(n_185273223));
	notech_nand3 i_54852532(.A(n_185273223), .B(n_185173222), .C(n_185073221
		), .Z(n_185473225));
	notech_ao4 i_58152500(.A(n_30697), .B(n_33288), .C(n_30689), .D(n_59465)
		, .Z(n_185773228));
	notech_ao4 i_57952501(.A(n_30693), .B(\nbus_11290[21] ), .C(n_30695), .D
		(\nbus_11283[21] ), .Z(n_185873229));
	notech_nand3 i_51353074(.A(n_181373192), .B(n_185873229), .C(n_185773228
		), .Z(n_75626083));
	notech_ao4 i_59352488(.A(n_327960907), .B(n_31494), .C(n_117626503), .D(n_33288
		), .Z(n_186373231));
	notech_ao4 i_59152490(.A(n_442668010), .B(\nbus_11283[21] ), .C(n_442868012
		), .D(nbus_11271[21]), .Z(n_186473232));
	notech_ao4 i_59252489(.A(n_59465), .B(n_117726504), .C(n_442568009), .D(\nbus_11290[21] 
		), .Z(n_186573233));
	notech_nand3 i_59552486(.A(n_186573233), .B(n_186473232), .C(n_186373231
		), .Z(n_186773235));
	notech_ao4 i_60452477(.A(n_33292), .B(n_30697), .C(n_59466), .D(n_30689)
		, .Z(n_187073238));
	notech_ao4 i_60352478(.A(n_30693), .B(\nbus_11290[20] ), .C(n_30695), .D
		(\nbus_11283[20] ), .Z(n_187173239));
	notech_and3 i_51253075(.A(n_375575066), .B(n_187173239), .C(n_187073238)
		, .Z(n_74526072));
	notech_ao4 i_61652465(.A(n_327960907), .B(n_31493), .C(n_117626503), .D(n_33292
		), .Z(n_187373241));
	notech_ao4 i_61452467(.A(n_442668010), .B(\nbus_11283[20] ), .C(n_442868012
		), .D(nbus_11271[20]), .Z(n_187473242));
	notech_ao4 i_61552466(.A(n_59466), .B(n_117726504), .C(n_442568009), .D(\nbus_11290[20] 
		), .Z(n_187573243));
	notech_and4 i_61952462(.A(n_187573243), .B(n_187473242), .C(n_187373241)
		, .D(n_74526072), .Z(n_187873246));
	notech_ao4 i_64852433(.A(n_305744491), .B(n_31499), .C(n_118426511), .D(n_33170
		), .Z(n_188073248));
	notech_ao4 i_64652435(.A(n_443268016), .B(\nbus_11283[23] ), .C(n_443168015
		), .D(nbus_11271[23]), .Z(n_188173249));
	notech_ao4 i_64752434(.A(n_109226419), .B(n_118526512), .C(n_443368017),
		 .D(\nbus_11290[23] ), .Z(n_188273250));
	notech_nand3 i_65052431(.A(n_188273250), .B(n_188173249), .C(n_188073248
		), .Z(n_188473252));
	notech_ao4 i_66452417(.A(n_305744491), .B(n_31496), .C(n_118426511), .D(n_33284
		), .Z(n_188773255));
	notech_ao4 i_66252419(.A(n_443268016), .B(\nbus_11283[22] ), .C(n_443168015
		), .D(nbus_11271[22]), .Z(n_188873256));
	notech_ao4 i_66352418(.A(n_59464), .B(n_118526512), .C(n_443368017), .D(\nbus_11290[22] 
		), .Z(n_188973257));
	notech_and4 i_66752414(.A(n_188973257), .B(n_188873256), .C(n_188773255)
		, .D(n_354467708), .Z(n_189273260));
	notech_ao4 i_68052401(.A(n_305744491), .B(n_31494), .C(n_118426511), .D(n_33288
		), .Z(n_189473262));
	notech_ao4 i_67852403(.A(n_443268016), .B(\nbus_11283[21] ), .C(n_443168015
		), .D(nbus_11271[21]), .Z(n_189573263));
	notech_ao4 i_67952402(.A(n_59465), .B(n_118526512), .C(n_443368017), .D(\nbus_11290[21] 
		), .Z(n_189673264));
	notech_nand3 i_68252399(.A(n_189673264), .B(n_189573263), .C(n_189473262
		), .Z(n_189873266));
	notech_ao4 i_69652385(.A(n_305744491), .B(n_31493), .C(n_118426511), .D(n_33292
		), .Z(n_190173269));
	notech_ao4 i_69452387(.A(n_443268016), .B(\nbus_11283[20] ), .C(n_443168015
		), .D(nbus_11271[20]), .Z(n_190273270));
	notech_ao4 i_69552386(.A(n_59466), .B(n_118526512), .C(n_443368017), .D(\nbus_11290[20] 
		), .Z(n_190373271));
	notech_and4 i_69952382(.A(n_190373271), .B(n_190273270), .C(n_190173269)
		, .D(n_74526072), .Z(n_190673274));
	notech_ao4 i_74452337(.A(n_379264323), .B(n_31499), .C(n_119226519), .D(n_33170
		), .Z(n_190873276));
	notech_ao4 i_74252339(.A(n_443768021), .B(\nbus_11283[23] ), .C(n_443668020
		), .D(nbus_11271[23]), .Z(n_190973277));
	notech_ao4 i_74352338(.A(n_109226419), .B(n_119326520), .C(n_443868022),
		 .D(\nbus_11290[23] ), .Z(n_191073278));
	notech_nand3 i_74652335(.A(n_191073278), .B(n_190973277), .C(n_190873276
		), .Z(n_191273280));
	notech_ao4 i_77652305(.A(n_379264323), .B(n_31494), .C(n_119226519), .D(n_33288
		), .Z(n_191573283));
	notech_ao4 i_77452307(.A(n_443768021), .B(\nbus_11283[21] ), .C(n_443668020
		), .D(nbus_11271[21]), .Z(n_191673284));
	notech_ao4 i_77552306(.A(n_59465), .B(n_119326520), .C(n_443868022), .D(\nbus_11290[21] 
		), .Z(n_191773285));
	notech_nand3 i_78052303(.A(n_191773285), .B(n_191673284), .C(n_191573283
		), .Z(n_191973287));
	notech_ao4 i_79452289(.A(n_379264323), .B(n_31493), .C(n_119226519), .D(n_33292
		), .Z(n_192273290));
	notech_ao4 i_79252291(.A(n_443768021), .B(\nbus_11283[20] ), .C(n_443668020
		), .D(nbus_11271[20]), .Z(n_192373291));
	notech_ao4 i_79352290(.A(n_59466), .B(n_119326520), .C(\nbus_11290[20] )
		, .D(n_443868022), .Z(n_192473292));
	notech_and4 i_79852286(.A(n_192473292), .B(n_192373291), .C(n_192273290)
		, .D(n_74526072), .Z(n_192773295));
	notech_ao4 i_84252243(.A(n_57363), .B(\nbus_11283[23] ), .C(n_303922064)
		, .D(nbus_11271[23]), .Z(n_192973297));
	notech_ao4 i_84352242(.A(n_57320), .B(n_109226419), .C(n_57362), .D(\nbus_11290[23] 
		), .Z(n_193173299));
	notech_ao4 i_84452241(.A(n_386864399), .B(n_31499), .C(n_57319), .D(n_33170
		), .Z(n_193273300));
	notech_and4 i_84752238(.A(n_193273300), .B(n_193173299), .C(n_192973297)
		, .D(n_180473183), .Z(n_193473302));
	notech_ao4 i_87452211(.A(n_57363), .B(\nbus_11283[21] ), .C(n_303922064)
		, .D(nbus_11271[21]), .Z(n_193673304));
	notech_ao4 i_87552210(.A(n_57320), .B(n_59465), .C(n_57362), .D(\nbus_11290[21] 
		), .Z(n_193873306));
	notech_ao4 i_87652209(.A(n_386864399), .B(n_31494), .C(n_57319), .D(n_33288
		), .Z(n_193973307));
	notech_and4 i_87952206(.A(n_193973307), .B(n_193873306), .C(n_193673304)
		, .D(n_181373192), .Z(n_194173309));
	notech_ao4 i_89052195(.A(n_57363), .B(\nbus_11283[20] ), .C(n_303922064)
		, .D(nbus_11271[20]), .Z(n_194373311));
	notech_ao4 i_89152194(.A(n_57320), .B(n_59466), .C(n_57362), .D(\nbus_11290[20] 
		), .Z(n_194573313));
	notech_ao4 i_89252193(.A(n_386864399), .B(n_31493), .C(n_57319), .D(n_33292
		), .Z(n_194673314));
	notech_and4 i_89552190(.A(n_194673314), .B(n_194573313), .C(n_194373311)
		, .D(n_375575066), .Z(n_194873316));
	notech_ao4 i_94052145(.A(n_58088), .B(n_31499), .C(n_324778256), .D(n_33170
		), .Z(n_195073318));
	notech_ao4 i_93852147(.A(n_57201), .B(\nbus_11283[23] ), .C(n_324978258)
		, .D(nbus_11271[23]), .Z(n_195173319));
	notech_ao4 i_93952146(.A(n_109226419), .B(n_324878257), .C(n_57200), .D(\nbus_11290[23] 
		), .Z(n_195273320));
	notech_nand3 i_94252143(.A(n_195273320), .B(n_195173319), .C(n_195073318
		), .Z(n_195473322));
	notech_ao4 i_97252113(.A(n_58088), .B(n_31494), .C(n_324778256), .D(n_33288
		), .Z(n_195773325));
	notech_ao4 i_97052115(.A(n_57201), .B(\nbus_11283[21] ), .C(n_324978258)
		, .D(nbus_11271[21]), .Z(n_195873326));
	notech_ao4 i_97152114(.A(n_59465), .B(n_324878257), .C(n_57200), .D(\nbus_11290[21] 
		), .Z(n_195973327));
	notech_nand3 i_97452111(.A(n_195973327), .B(n_195873326), .C(n_195773325
		), .Z(n_196173329));
	notech_ao4 i_98852097(.A(n_58088), .B(n_31493), .C(n_324778256), .D(n_33292
		), .Z(n_196473332));
	notech_ao4 i_98652099(.A(n_57201), .B(\nbus_11283[20] ), .C(n_324978258)
		, .D(nbus_11271[20]), .Z(n_196573333));
	notech_ao4 i_98752098(.A(n_59466), .B(n_324878257), .C(n_57200), .D(\nbus_11290[20] 
		), .Z(n_196673334));
	notech_and4 i_99152094(.A(n_196673334), .B(n_196573333), .C(n_196473332)
		, .D(n_74526072), .Z(n_196973337));
	notech_ao4 i_117851912(.A(n_59464), .B(n_122926556), .C(n_122626553), .D
		(\nbus_11290[22] ), .Z(n_197173339));
	notech_ao4 i_117951911(.A(n_331060938), .B(n_31496), .C(n_122826555), .D
		(n_33284), .Z(n_197273340));
	notech_nand2 i_118251908(.A(n_197273340), .B(n_197173339), .Z(n_197373341
		));
	notech_ao4 i_118051910(.A(n_61099), .B(n_30853), .C(n_57012), .D(n_31530
		), .Z(n_197473342));
	notech_ao4 i_117651914(.A(n_333360961), .B(n_33329), .C(n_333260960), .D
		(n_33328), .Z(n_197573343));
	notech_ao4 i_117751913(.A(n_122726554), .B(\nbus_11283[22] ), .C(nbus_11271
		[22]), .D(n_337361001), .Z(n_197673344));
	notech_nand3 i_118351907(.A(n_197673344), .B(n_197573343), .C(n_197473342
		), .Z(n_197873346));
	notech_ao4 i_120151889(.A(n_59465), .B(n_122926556), .C(n_122626553), .D
		(\nbus_11290[21] ), .Z(n_198173349));
	notech_ao4 i_120251888(.A(n_331060938), .B(n_31494), .C(n_122826555), .D
		(n_33288), .Z(n_198273350));
	notech_nand2 i_120551885(.A(n_198273350), .B(n_198173349), .Z(n_198373351
		));
	notech_ao4 i_120351887(.A(n_61099), .B(n_30852), .C(n_57006), .D(n_31529
		), .Z(n_198473352));
	notech_ao4 i_119951891(.A(n_333360961), .B(n_33331), .C(n_333260960), .D
		(n_33330), .Z(n_198573353));
	notech_ao4 i_120051890(.A(n_122726554), .B(\nbus_11283[21] ), .C(n_337361001
		), .D(nbus_11271[21]), .Z(n_198673354));
	notech_nand3 i_120651884(.A(n_198673354), .B(n_198573353), .C(n_198473352
		), .Z(n_198873356));
	notech_ao4 i_122451866(.A(n_59466), .B(n_122926556), .C(n_122626553), .D
		(\nbus_11290[20] ), .Z(n_199173359));
	notech_ao4 i_122551865(.A(n_331060938), .B(n_31493), .C(n_122826555), .D
		(n_33292), .Z(n_199273360));
	notech_nand2 i_122851862(.A(n_199273360), .B(n_199173359), .Z(n_199373361
		));
	notech_ao4 i_122651864(.A(n_61099), .B(n_30851), .C(n_57012), .D(n_31528
		), .Z(n_199473362));
	notech_ao4 i_122251868(.A(n_333360961), .B(n_33333), .C(n_333260960), .D
		(n_33332), .Z(n_199573363));
	notech_ao4 i_122351867(.A(n_122726554), .B(\nbus_11283[20] ), .C(n_337361001
		), .D(nbus_11271[20]), .Z(n_199673364));
	notech_nand3 i_122951861(.A(n_199673364), .B(n_199573363), .C(n_199473362
		), .Z(n_199873366));
	notech_ao4 i_134951741(.A(n_124826575), .B(n_101026337), .C(n_124526572)
		, .D(\nbus_11290[25] ), .Z(n_200173369));
	notech_ao4 i_135051740(.A(n_328660914), .B(n_31501), .C(n_124726574), .D
		(n_33172), .Z(n_200273370));
	notech_nand2 i_135351737(.A(n_200273370), .B(n_200173369), .Z(n_200373371
		));
	notech_ao4 i_135151739(.A(n_61103), .B(n_30831), .C(n_57012), .D(n_31533
		), .Z(n_200473372));
	notech_ao4 i_134751743(.A(n_330460932), .B(n_33335), .C(n_330560933), .D
		(n_33334), .Z(n_200573373));
	notech_ao4 i_134851742(.A(n_124626573), .B(\nbus_11283[25] ), .C(n_337561003
		), .D(nbus_11271[25]), .Z(n_200673374));
	notech_nand3 i_135451736(.A(n_200673374), .B(n_200573373), .C(n_200473372
		), .Z(n_200873376));
	notech_ao4 i_139551695(.A(n_109226419), .B(n_124826575), .C(n_124526572)
		, .D(\nbus_11290[23] ), .Z(n_201173379));
	notech_ao4 i_139651694(.A(n_328660914), .B(n_31499), .C(n_124726574), .D
		(n_33170), .Z(n_201273380));
	notech_nand2 i_139951691(.A(n_201273380), .B(n_201173379), .Z(n_201373381
		));
	notech_ao4 i_139751693(.A(n_61103), .B(n_30827), .C(n_57012), .D(n_31531
		), .Z(n_201473382));
	notech_ao4 i_139351697(.A(n_330460932), .B(n_33337), .C(n_330560933), .D
		(n_33336), .Z(n_201573383));
	notech_ao4 i_139451696(.A(n_124626573), .B(\nbus_11283[23] ), .C(n_337561003
		), .D(nbus_11271[23]), .Z(n_201673384));
	notech_nand3 i_140051690(.A(n_201673384), .B(n_201573383), .C(n_201473382
		), .Z(n_201873386));
	notech_ao4 i_141851672(.A(n_59464), .B(n_124826575), .C(n_124526572), .D
		(\nbus_11290[22] ), .Z(n_202173389));
	notech_ao4 i_141951671(.A(n_328660914), .B(n_31496), .C(n_124726574), .D
		(n_33284), .Z(n_202273390));
	notech_nand2 i_142251668(.A(n_202273390), .B(n_202173389), .Z(n_202373391
		));
	notech_ao4 i_142051670(.A(n_61103), .B(n_30826), .C(n_57012), .D(n_31530
		), .Z(n_202473392));
	notech_ao4 i_141651674(.A(n_330460932), .B(n_33339), .C(n_330560933), .D
		(n_33338), .Z(n_202573393));
	notech_ao4 i_141751673(.A(n_124626573), .B(\nbus_11283[22] ), .C(nbus_11271
		[22]), .D(n_337561003), .Z(n_202673394));
	notech_nand3 i_142351667(.A(n_202673394), .B(n_202573393), .C(n_202473392
		), .Z(n_202873396));
	notech_ao4 i_144151649(.A(n_59465), .B(n_124826575), .C(n_124526572), .D
		(\nbus_11290[21] ), .Z(n_203173399));
	notech_ao4 i_144251648(.A(n_328660914), .B(n_31494), .C(n_124726574), .D
		(n_33288), .Z(n_203273400));
	notech_nand2 i_144551645(.A(n_203273400), .B(n_203173399), .Z(n_203373401
		));
	notech_ao4 i_144351647(.A(n_61103), .B(n_30825), .C(n_57006), .D(n_31529
		), .Z(n_203473402));
	notech_ao4 i_143951651(.A(n_330460932), .B(n_33341), .C(n_330560933), .D
		(n_33340), .Z(n_203573403));
	notech_ao4 i_144051650(.A(n_124626573), .B(\nbus_11283[21] ), .C(n_337561003
		), .D(nbus_11271[21]), .Z(n_203673404));
	notech_nand3 i_144651644(.A(n_203673404), .B(n_203573403), .C(n_203473402
		), .Z(n_203873406));
	notech_ao4 i_146451626(.A(n_59466), .B(n_124826575), .C(n_124526572), .D
		(\nbus_11290[20] ), .Z(n_204173409));
	notech_ao4 i_146551625(.A(n_328660914), .B(n_31493), .C(n_124726574), .D
		(n_33292), .Z(n_204273410));
	notech_nand2 i_146851622(.A(n_204273410), .B(n_204173409), .Z(n_204373411
		));
	notech_ao4 i_146651624(.A(n_61103), .B(n_30824), .C(n_57006), .D(n_31528
		), .Z(n_204473412));
	notech_ao4 i_146251628(.A(n_330460932), .B(n_33343), .C(n_330560933), .D
		(n_33342), .Z(n_204573413));
	notech_ao4 i_146351627(.A(n_124626573), .B(\nbus_11283[20] ), .C(n_337561003
		), .D(nbus_11271[20]), .Z(n_204673414));
	notech_nand3 i_146951621(.A(n_204673414), .B(n_204573413), .C(n_204473412
		), .Z(n_204873416));
	notech_ao4 i_151551575(.A(n_305644490), .B(n_31499), .C(n_125326580), .D
		(n_33170), .Z(n_205173419));
	notech_ao4 i_151351577(.A(n_302744461), .B(\nbus_11283[23] ), .C(n_387564406
		), .D(nbus_11271[23]), .Z(n_205273420));
	notech_ao4 i_151451576(.A(n_109226419), .B(n_125426581), .C(n_302844462)
		, .D(\nbus_11290[23] ), .Z(n_205373421));
	notech_nand3 i_151751573(.A(n_205373421), .B(n_205273420), .C(n_205173419
		), .Z(n_205573423));
	notech_ao4 i_154751543(.A(n_305644490), .B(n_31494), .C(n_125326580), .D
		(n_33288), .Z(n_205873426));
	notech_ao4 i_154551545(.A(n_302744461), .B(\nbus_11283[21] ), .C(n_387564406
		), .D(nbus_11271[21]), .Z(n_205973427));
	notech_ao4 i_154651544(.A(n_59465), .B(n_125426581), .C(n_302844462), .D
		(\nbus_11290[21] ), .Z(n_206073428));
	notech_nand3 i_154951541(.A(n_206073428), .B(n_205973427), .C(n_205873426
		), .Z(n_206273430));
	notech_ao4 i_156351527(.A(n_305644490), .B(n_31493), .C(n_125326580), .D
		(n_33292), .Z(n_206573433));
	notech_ao4 i_156151529(.A(n_302744461), .B(\nbus_11283[20] ), .C(n_387564406
		), .D(nbus_11271[20]), .Z(n_206673434));
	notech_ao4 i_156251528(.A(n_59466), .B(n_125426581), .C(n_302844462), .D
		(\nbus_11290[20] ), .Z(n_206773435));
	notech_and4 i_156651524(.A(n_206773435), .B(n_206673434), .C(n_206573433
		), .D(n_74526072), .Z(n_207073438));
	notech_ao4 i_163551455(.A(n_126926596), .B(n_33170), .C(n_109226419), .D
		(n_127026597), .Z(n_207273440));
	notech_ao4 i_163651454(.A(n_337861006), .B(n_31499), .C(n_26600), .D(n_31531
		), .Z(n_207373441));
	notech_ao4 i_163251458(.A(n_126126588), .B(n_32082), .C(n_26585), .D(n_31014
		), .Z(n_207573443));
	notech_ao4 i_163351457(.A(n_337761005), .B(nbus_11271[23]), .C(n_125926586
		), .D(n_33344), .Z(n_207773445));
	notech_ao4 i_163451456(.A(n_126826595), .B(\nbus_11290[23] ), .C(n_126726594
		), .D(\nbus_11283[23] ), .Z(n_207873446));
	notech_and4 i_164051450(.A(n_207873446), .B(n_207773445), .C(n_207573443
		), .D(n_173073115), .Z(n_208073448));
	notech_and3 i_164151449(.A(n_207373441), .B(n_207273440), .C(n_208073448
		), .Z(n_208173449));
	notech_ao4 i_166051430(.A(n_126926596), .B(n_33284), .C(n_127026597), .D
		(n_59464), .Z(n_208373451));
	notech_ao4 i_166151429(.A(n_337861006), .B(n_31496), .C(n_26600), .D(n_31530
		), .Z(n_208473452));
	notech_ao4 i_165751433(.A(n_126126588), .B(n_32081), .C(n_26585), .D(n_31012
		), .Z(n_208673454));
	notech_ao4 i_165851432(.A(n_337761005), .B(nbus_11271[22]), .C(n_125926586
		), .D(n_33345), .Z(n_208873456));
	notech_ao4 i_165951431(.A(n_126826595), .B(\nbus_11290[22] ), .C(n_126726594
		), .D(\nbus_11283[22] ), .Z(n_208973457));
	notech_and4 i_166551425(.A(n_208973457), .B(n_208873456), .C(n_208673454
		), .D(n_174373128), .Z(n_209173459));
	notech_and3 i_166651424(.A(n_208473452), .B(n_208373451), .C(n_209173459
		), .Z(n_209273460));
	notech_ao4 i_168551405(.A(n_126926596), .B(n_33288), .C(n_59465), .D(n_127026597
		), .Z(n_209473462));
	notech_ao4 i_168651404(.A(n_337861006), .B(n_31494), .C(n_26600), .D(n_31529
		), .Z(n_209573463));
	notech_ao4 i_168251408(.A(n_126126588), .B(n_32080), .C(n_26585), .D(n_31010
		), .Z(n_209773465));
	notech_ao4 i_168351407(.A(n_337761005), .B(nbus_11271[21]), .C(n_125926586
		), .D(n_33346), .Z(n_209973467));
	notech_ao4 i_168451406(.A(n_126826595), .B(\nbus_11290[21] ), .C(n_126726594
		), .D(\nbus_11283[21] ), .Z(n_210073468));
	notech_and4 i_169051400(.A(n_210073468), .B(n_209973467), .C(n_209773465
		), .D(n_176273141), .Z(n_210273470));
	notech_and3 i_169151399(.A(n_209573463), .B(n_209473462), .C(n_210273470
		), .Z(n_210373471));
	notech_ao4 i_171051380(.A(n_33292), .B(n_126926596), .C(n_59466), .D(n_127026597
		), .Z(n_210573473));
	notech_ao4 i_171151379(.A(n_337861006), .B(n_31493), .C(n_26600), .D(n_31528
		), .Z(n_210673474));
	notech_ao4 i_170751383(.A(n_126126588), .B(n_32079), .C(n_26585), .D(n_31008
		), .Z(n_210873476));
	notech_ao4 i_170851382(.A(n_337761005), .B(nbus_11271[20]), .C(n_125926586
		), .D(n_33347), .Z(n_211073478));
	notech_ao4 i_170951381(.A(n_126826595), .B(\nbus_11290[20] ), .C(n_126726594
		), .D(\nbus_11283[20] ), .Z(n_211173479));
	notech_and4 i_171551375(.A(n_211173479), .B(n_211073478), .C(n_210873476
		), .D(n_177573154), .Z(n_211373481));
	notech_and3 i_171651374(.A(n_210673474), .B(n_210573473), .C(n_211373481
		), .Z(n_211473482));
	notech_ao4 i_176251328(.A(n_58083), .B(n_31499), .C(n_324178250), .D(n_33170
		), .Z(n_211673484));
	notech_ao4 i_176051330(.A(n_57213), .B(\nbus_11283[23] ), .C(n_301822043
		), .D(nbus_11271[23]), .Z(n_211773485));
	notech_ao4 i_176151329(.A(n_109226419), .B(n_324278251), .C(n_57217), .D
		(\nbus_11290[23] ), .Z(n_211873486));
	notech_nand3 i_176451326(.A(n_211873486), .B(n_211773485), .C(n_211673484
		), .Z(n_212073488));
	notech_ao4 i_179451297(.A(n_301822043), .B(nbus_11271[21]), .C(n_383264363
		), .D(n_61625), .Z(n_212373491));
	notech_ao4 i_179551296(.A(n_57217), .B(\nbus_11290[21] ), .C(n_57213), .D
		(\nbus_11283[21] ), .Z(n_212573493));
	notech_ao4 i_179651295(.A(n_324178250), .B(n_33288), .C(n_59465), .D(n_324278251
		), .Z(n_212673494));
	notech_and4 i_179951292(.A(n_212673494), .B(n_212573493), .C(n_212373491
		), .D(n_179173170), .Z(n_212873496));
	notech_ao4 i_181451278(.A(n_58083), .B(n_31493), .C(n_324178250), .D(n_33292
		), .Z(n_213173499));
	notech_ao4 i_181251280(.A(n_57213), .B(\nbus_11283[20] ), .C(n_301822043
		), .D(nbus_11271[20]), .Z(n_213273500));
	notech_ao4 i_181351279(.A(n_59466), .B(n_324278251), .C(\nbus_11290[20] 
		), .D(n_57217), .Z(n_213373501));
	notech_and4 i_181751275(.A(n_213373501), .B(n_213273500), .C(n_213173499
		), .D(n_74526072), .Z(n_213673504));
	notech_ao4 i_187151222(.A(n_109226419), .B(n_365328693), .C(n_365528695)
		, .D(\nbus_11290[23] ), .Z(n_213873506));
	notech_ao4 i_186751226(.A(n_382264353), .B(n_31499), .C(n_56036), .D(n_32571
		), .Z(n_213973507));
	notech_and3 i_186951224(.A(n_180473183), .B(n_213973507), .C(n_180573184
		), .Z(n_214173509));
	notech_and4 i_187351220(.A(n_213873506), .B(n_180673185), .C(n_214173509
		), .D(n_180973188), .Z(n_214473512));
	notech_ao4 i_190951184(.A(n_59465), .B(n_365328693), .C(n_365528695), .D
		(\nbus_11290[21] ), .Z(n_214673514));
	notech_ao4 i_190551188(.A(n_382264353), .B(n_31494), .C(n_61688), .D(n_31529
		), .Z(n_214873516));
	notech_and4 i_190751186(.A(n_5774), .B(n_214873516), .C(n_181273191), .D
		(n_181573194), .Z(n_215073518));
	notech_and4 i_191151182(.A(n_215073518), .B(n_214673514), .C(n_181673195
		), .D(n_181973198), .Z(n_215373521));
	notech_ao4 i_208851006(.A(n_131426641), .B(nbus_11271[23]), .C(n_56036),
		 .D(n_32551), .Z(n_215573523));
	notech_ao4 i_208951005(.A(n_387964410), .B(\nbus_11290[23] ), .C(n_387864409
		), .D(\nbus_11283[23] ), .Z(n_215773525));
	notech_ao4 i_209051004(.A(n_131526642), .B(n_33170), .C(n_109226419), .D
		(n_131626643), .Z(n_215873526));
	notech_and4 i_209351001(.A(n_215873526), .B(n_215773525), .C(n_215573523
		), .D(n_183573207), .Z(n_216073528));
	notech_ao4 i_214250952(.A(n_131426641), .B(nbus_11271[20]), .C(n_56036),
		 .D(n_32546), .Z(n_216373531));
	notech_ao4 i_214350951(.A(n_387964410), .B(\nbus_11290[20] ), .C(n_387864409
		), .D(\nbus_11283[20] ), .Z(n_216573533));
	notech_ao4 i_214450950(.A(n_33292), .B(n_131526642), .C(n_59466), .D(n_131626643
		), .Z(n_216673534));
	notech_and4 i_214750947(.A(n_216673534), .B(n_216573533), .C(n_216373531
		), .D(n_184573216), .Z(n_216873536));
	notech_and4 i_89045564(.A(n_286763769), .B(n_116742608), .C(n_29560), .D
		(n_386764398), .Z(n_217173539));
	notech_nand3 i_29852(.A(n_290663806), .B(instrc[117]), .C(n_63782), .Z(n_217373541
		));
	notech_or4 i_103445422(.A(n_318060808), .B(n_2577), .C(n_286263764), .D(n_386664397
		), .Z(n_217473542));
	notech_or4 i_103545421(.A(n_318060808), .B(n_2577), .C(n_286263764), .D(n_29553
		), .Z(n_217573543));
	notech_or2 i_103645420(.A(n_386964400), .B(n_29553), .Z(n_217673544));
	notech_or4 i_60440090(.A(n_61917), .B(n_61901), .C(n_61889), .D(n_1861),
		 .Z(n_218373551));
	notech_and3 i_8339993(.A(n_22752), .B(n_1832), .C(n_227173639), .Z(n_218573553
		));
	notech_ao4 i_8239994(.A(n_61625), .B(n_2974), .C(n_23367), .D(nbus_11291
		[1]), .Z(n_218673554));
	notech_and2 i_8039996(.A(n_1832), .B(n_367275008), .Z(n_218873556));
	notech_and2 i_7939997(.A(n_1832), .B(n_364274979), .Z(n_218973557));
	notech_and2 i_7839998(.A(n_361374951), .B(n_1832), .Z(n_219073558));
	notech_and4 i_8539991(.A(n_301274364), .B(n_242373791), .C(n_360074938),
		 .D(n_301474366), .Z(n_219173559));
	notech_and2 i_8639990(.A(n_25467), .B(n_1824), .Z(n_219273560));
	notech_ao4 i_7739999(.A(n_23367), .B(nbus_11291[8]), .C(n_220973577), .D
		(n_61623), .Z(n_219373561));
	notech_ao4 i_7640000(.A(n_23367), .B(nbus_11291[9]), .C(n_220973577), .D
		(n_61623), .Z(n_219573563));
	notech_ao4 i_7540001(.A(n_23367), .B(nbus_11291[10]), .C(n_220973577), .D
		(n_61623), .Z(n_219773565));
	notech_ao4 i_7440002(.A(n_23367), .B(nbus_11291[11]), .C(n_220973577), .D
		(n_61623), .Z(n_219973567));
	notech_ao4 i_7340003(.A(n_23367), .B(nbus_11291[12]), .C(n_220973577), .D
		(n_61623), .Z(n_220173569));
	notech_ao4 i_7240004(.A(n_23367), .B(nbus_11291[13]), .C(n_220973577), .D
		(n_61623), .Z(n_220373571));
	notech_ao4 i_7140005(.A(n_23367), .B(nbus_11291[14]), .C(n_220973577), .D
		(n_61625), .Z(n_220573573));
	notech_ao4 i_7040006(.A(n_23367), .B(nbus_11291[15]), .C(n_61625), .D(n_220973577
		), .Z(n_220773575));
	notech_and3 i_55639528(.A(n_25467), .B(n_2973), .C(n_1808), .Z(n_220973577
		));
	notech_and4 i_6940007(.A(n_23373), .B(n_23371), .C(n_301574367), .D(n_221173579
		), .Z(n_221073578));
	notech_or2 i_57839506(.A(n_23367), .B(nbus_11291[16]), .Z(n_221173579)
		);
	notech_and4 i_6840008(.A(n_23373), .B(n_23371), .C(n_301574367), .D(n_221373581
		), .Z(n_221273580));
	notech_or2 i_60239484(.A(n_23367), .B(nbus_11291[17]), .Z(n_221373581)
		);
	notech_and4 i_6740009(.A(n_23373), .B(n_23371), .C(n_301574367), .D(n_221573583
		), .Z(n_221473582));
	notech_or2 i_62639462(.A(n_23367), .B(nbus_11291[18]), .Z(n_221573583)
		);
	notech_and4 i_6640010(.A(n_23373), .B(n_23371), .C(n_301574367), .D(n_221773585
		), .Z(n_221673584));
	notech_or2 i_65439440(.A(n_23367), .B(nbus_11291[19]), .Z(n_221773585)
		);
	notech_and4 i_6540011(.A(n_23373), .B(n_23371), .C(n_301574367), .D(n_221973587
		), .Z(n_221873586));
	notech_or2 i_67639418(.A(n_23367), .B(nbus_11291[20]), .Z(n_221973587)
		);
	notech_and4 i_6440012(.A(n_23373), .B(n_23371), .C(n_301574367), .D(n_222173589
		), .Z(n_222073588));
	notech_or2 i_70039396(.A(n_23367), .B(nbus_11291[21]), .Z(n_222173589)
		);
	notech_and4 i_6340013(.A(n_23373), .B(n_23371), .C(n_301574367), .D(n_222373591
		), .Z(n_222273590));
	notech_or2 i_72639374(.A(n_23367), .B(nbus_11291[22]), .Z(n_222373591)
		);
	notech_and4 i_6240014(.A(n_23373), .B(n_23371), .C(n_301574367), .D(n_222573593
		), .Z(n_222473592));
	notech_or2 i_75039352(.A(n_57896), .B(nbus_11291[23]), .Z(n_222573593)
		);
	notech_and4 i_6140015(.A(n_23373), .B(n_23371), .C(n_301574367), .D(n_222773595
		), .Z(n_222673594));
	notech_or2 i_77339330(.A(n_57896), .B(nbus_11291[24]), .Z(n_222773595)
		);
	notech_and4 i_6040016(.A(n_23373), .B(n_23371), .C(n_301574367), .D(n_222973597
		), .Z(n_222873596));
	notech_or2 i_79639308(.A(n_57896), .B(nbus_11291[25]), .Z(n_222973597)
		);
	notech_and4 i_5940017(.A(n_23373), .B(n_23371), .C(n_301574367), .D(n_223173599
		), .Z(n_223073598));
	notech_or2 i_81939286(.A(n_57896), .B(nbus_11291[26]), .Z(n_223173599)
		);
	notech_and4 i_5840018(.A(n_23373), .B(n_23371), .C(n_301574367), .D(n_223373601
		), .Z(n_223273600));
	notech_or2 i_84139264(.A(n_57896), .B(nbus_11291[27]), .Z(n_223373601)
		);
	notech_and4 i_5740019(.A(n_23373), .B(n_57907), .C(n_301574367), .D(n_223573603
		), .Z(n_223473602));
	notech_or2 i_86339242(.A(n_57896), .B(nbus_11291[28]), .Z(n_223573603)
		);
	notech_and4 i_5640020(.A(n_23373), .B(n_57907), .C(n_301574367), .D(n_223773605
		), .Z(n_223673604));
	notech_or2 i_88639220(.A(n_57896), .B(nbus_11291[29]), .Z(n_223773605)
		);
	notech_and4 i_5540021(.A(n_23373), .B(n_57907), .C(n_301574367), .D(n_223973607
		), .Z(n_223873606));
	notech_or2 i_90839198(.A(n_57896), .B(nbus_11291[30]), .Z(n_223973607)
		);
	notech_and4 i_5440022(.A(n_23373), .B(n_57907), .C(n_301574367), .D(n_224173609
		), .Z(n_224073608));
	notech_or2 i_93039176(.A(n_57896), .B(nbus_11291[31]), .Z(n_224173609)
		);
	notech_nand2 i_12039956(.A(nbus_135[0]), .B(n_22746), .Z(n_224573613));
	notech_nao3 i_11339963(.A(opa_0[0]), .B(n_61688), .C(n_1803), .Z(n_225273620
		));
	notech_or2 i_10639970(.A(n_1828), .B(n_33169), .Z(n_225973627));
	notech_nand2 i_9939977(.A(n_6259), .B(n_23330), .Z(n_226673634));
	notech_or2 i_12139955(.A(n_57896), .B(nbus_11291[0]), .Z(n_227173639));
	notech_nand2 i_15139926(.A(nbus_135[1]), .B(n_22746), .Z(n_227473642));
	notech_nao3 i_14439933(.A(opa_0[1]), .B(n_61688), .C(n_1803), .Z(n_228173649
		));
	notech_or2 i_13739940(.A(n_1828), .B(n_33103), .Z(n_228873656));
	notech_nand2 i_21439865(.A(nbus_135[3]), .B(n_22746), .Z(n_230373671));
	notech_nao3 i_20739872(.A(opa_0[3]), .B(n_61688), .C(n_1803), .Z(n_231073678
		));
	notech_or2 i_20039879(.A(n_1828), .B(n_33118), .Z(n_231773685));
	notech_nand2 i_24639834(.A(nbus_135[4]), .B(n_22746), .Z(n_233473702));
	notech_nao3 i_23939841(.A(opa_0[4]), .B(n_61688), .C(n_1803), .Z(n_234173709
		));
	notech_or2 i_23239848(.A(n_1828), .B(n_33104), .Z(n_234873716));
	notech_nand2 i_27739803(.A(nbus_135[6]), .B(n_22746), .Z(n_236573733));
	notech_nao3 i_27039810(.A(opa_0[6]), .B(n_61684), .C(n_1803), .Z(n_237273740
		));
	notech_or2 i_26339817(.A(n_1828), .B(n_33166), .Z(n_237973747));
	notech_nao3 i_30039780(.A(nbus_138[7]), .B(n_61684), .C(n_1802), .Z(n_239673764
		));
	notech_nand3 i_29739783(.A(mul64[7]), .B(n_30648), .C(n_61684), .Z(n_239973767
		));
	notech_or2 i_29439786(.A(n_22979), .B(n_58902), .Z(n_240273770));
	notech_or2 i_29139789(.A(n_1828), .B(n_33165), .Z(n_240573773));
	notech_nao3 i_28839792(.A(nbus_14541[7]), .B(n_32241), .C(n_58506), .Z(n_240873776
		));
	notech_or4 i_28539795(.A(n_30926), .B(n_30691), .C(n_19548), .D(n_32458)
		, .Z(n_241173779));
	notech_or2 i_28239798(.A(n_23345), .B(\nbus_11290[7] ), .Z(n_241473782)
		);
	notech_or2 i_31139769(.A(n_57896), .B(nbus_11291[7]), .Z(n_242373791));
	notech_or2 i_32639754(.A(n_23345), .B(\nbus_11290[8] ), .Z(n_244273810)
		);
	notech_or2 i_35639724(.A(n_23345), .B(\nbus_11290[9] ), .Z(n_247173839)
		);
	notech_or2 i_38739694(.A(n_23345), .B(\nbus_11290[10] ), .Z(n_250073868)
		);
	notech_nao3 i_41739664(.A(resa_arithbox[11]), .B(n_61684), .C(n_27914), 
		.Z(n_252973897));
	notech_nao3 i_44739634(.A(resa_arithbox[12]), .B(n_61684), .C(n_27914), 
		.Z(n_255873926));
	notech_nao3 i_47739604(.A(nbus_14541[13]), .B(n_32241), .C(n_58506), .Z(n_258773955
		));
	notech_nao3 i_50739574(.A(nbus_14541[14]), .B(n_32241), .C(n_58506), .Z(n_261673984
		));
	notech_nao3 i_53739544(.A(nbus_14541[15]), .B(n_32241), .C(n_58506), .Z(n_264574013
		));
	notech_nao3 i_57639508(.A(n_318760815), .B(cr3[16]), .C(n_58506), .Z(n_266174029
		));
	notech_nand2 i_57339511(.A(cr0[16]), .B(n_23351), .Z(n_266474032));
	notech_nao3 i_57039514(.A(nbus_140[16]), .B(n_61684), .C(n_27920), .Z(n_266774035
		));
	notech_or4 i_56539519(.A(n_30926), .B(n_30691), .C(n_19548), .D(n_32467)
		, .Z(n_267274040));
	notech_or4 i_56239522(.A(n_61723), .B(n_61890), .C(n_25467), .D(nbus_11271
		[0]), .Z(n_267574043));
	notech_nao3 i_55939525(.A(nbus_138[16]), .B(n_61684), .C(n_27919), .Z(n_267874046
		));
	notech_nao3 i_60139485(.A(cr2_reg[17]), .B(n_32268), .C(n_58506), .Z(n_268774047
		));
	notech_nao3 i_59939486(.A(n_318760815), .B(cr3[17]), .C(n_58506), .Z(n_269274050
		));
	notech_nand2 i_59639489(.A(\nbus_14542[17] ), .B(n_23351), .Z(n_269574053
		));
	notech_nao3 i_59339492(.A(nbus_140[17]), .B(n_61684), .C(n_27920), .Z(n_269874056
		));
	notech_or4 i_58839497(.A(n_30926), .B(n_30691), .C(n_19548), .D(n_32468)
		, .Z(n_270374061));
	notech_or4 i_58539500(.A(n_61889), .B(n_25467), .C(n_61723), .D(nbus_11271
		[1]), .Z(n_270674064));
	notech_nao3 i_58239503(.A(nbus_138[17]), .B(n_61684), .C(n_27919), .Z(n_270974067
		));
	notech_nao3 i_62539463(.A(cr2_reg[18]), .B(n_32268), .C(n_58506), .Z(n_271074068
		));
	notech_nao3 i_62439464(.A(n_318760815), .B(cr3[18]), .C(n_58506), .Z(n_271574071
		));
	notech_nand2 i_62139467(.A(\nbus_14542[18] ), .B(n_23351), .Z(n_271874074
		));
	notech_nao3 i_61739470(.A(nbus_140[18]), .B(n_61684), .C(n_27920), .Z(n_272174077
		));
	notech_or4 i_61239475(.A(n_30926), .B(n_30691), .C(n_19548), .D(n_32469)
		, .Z(n_272674082));
	notech_or4 i_60939478(.A(n_61890), .B(n_25467), .C(n_61723), .D(nbus_11271
		[2]), .Z(n_273374085));
	notech_nao3 i_60639481(.A(nbus_138[18]), .B(n_61688), .C(n_27919), .Z(n_273674088
		));
	notech_nao3 i_65339441(.A(cr2_reg[19]), .B(n_32268), .C(n_58506), .Z(n_273774089
		));
	notech_nao3 i_65239442(.A(n_318760815), .B(cr3[19]), .C(n_58506), .Z(n_274074092
		));
	notech_nand2 i_64739445(.A(\nbus_14542[19] ), .B(n_23351), .Z(n_274374095
		));
	notech_nao3 i_64339448(.A(nbus_140[19]), .B(n_61689), .C(n_27920), .Z(n_274674098
		));
	notech_or4 i_63739453(.A(n_30926), .B(n_30691), .C(n_19548), .D(n_32470)
		, .Z(n_275174103));
	notech_or4 i_63239456(.A(n_61890), .B(n_25467), .C(n_61723), .D(nbus_11271
		[3]), .Z(n_275474106));
	notech_nao3 i_62939459(.A(nbus_138[19]), .B(n_61689), .C(n_27919), .Z(n_275774109
		));
	notech_nao3 i_67539419(.A(cr2_reg[20]), .B(n_32268), .C(n_58506), .Z(n_275874110
		));
	notech_nao3 i_67439420(.A(n_318760815), .B(cr3[20]), .C(n_58506), .Z(n_276174113
		));
	notech_nand2 i_67139423(.A(\nbus_14542[20] ), .B(n_23351), .Z(n_276474116
		));
	notech_nao3 i_66839426(.A(nbus_140[20]), .B(n_61689), .C(n_27920), .Z(n_276774119
		));
	notech_or4 i_66339431(.A(n_30926), .B(n_30691), .C(n_19548), .D(n_32471)
		, .Z(n_277274124));
	notech_or4 i_66039434(.A(n_61889), .B(n_25467), .C(n_61723), .D(nbus_11271
		[4]), .Z(n_277574127));
	notech_nao3 i_65739437(.A(nbus_138[20]), .B(n_61689), .C(n_27919), .Z(n_277874130
		));
	notech_nao3 i_69839398(.A(n_318760815), .B(cr3[21]), .C(n_58506), .Z(n_278274134
		));
	notech_nand2 i_69439401(.A(\nbus_14542[21] ), .B(n_23351), .Z(n_278574137
		));
	notech_nao3 i_69139404(.A(nbus_140[21]), .B(n_61689), .C(n_27920), .Z(n_278874140
		));
	notech_or4 i_68539409(.A(n_30926), .B(n_30691), .C(n_19548), .D(n_32472)
		, .Z(n_279374145));
	notech_or4 i_68239412(.A(n_61718), .B(n_61889), .C(n_25467), .D(nbus_11271
		[5]), .Z(n_279674148));
	notech_nao3 i_67939415(.A(nbus_138[21]), .B(n_61689), .C(n_27919), .Z(n_279974151
		));
	notech_nao3 i_72539375(.A(cr2_reg[22]), .B(n_32268), .C(n_58506), .Z(n_280074152
		));
	notech_nao3 i_72439376(.A(cr3[22]), .B(n_318760815), .C(n_58506), .Z(n_280374155
		));
	notech_nand2 i_72139379(.A(\nbus_14542[22] ), .B(n_23351), .Z(n_280674158
		));
	notech_nao3 i_71839382(.A(nbus_140[22]), .B(n_61693), .C(n_27920), .Z(n_280974161
		));
	notech_or4 i_71339387(.A(n_30926), .B(n_30691), .C(n_19548), .D(n_32473)
		, .Z(n_281474166));
	notech_or4 i_70939390(.A(n_61718), .B(n_61889), .C(n_25467), .D(nbus_11271
		[6]), .Z(n_281774169));
	notech_nao3 i_70339393(.A(nbus_138[22]), .B(n_61689), .C(n_27919), .Z(n_282074172
		));
	notech_nao3 i_74939353(.A(cr2_reg[23]), .B(n_32268), .C(n_58506), .Z(n_282174173
		));
	notech_nao3 i_74839354(.A(n_318760815), .B(cr3[23]), .C(n_58506), .Z(n_282474176
		));
	notech_nand2 i_74539357(.A(\nbus_14542[23] ), .B(n_23351), .Z(n_282774179
		));
	notech_nao3 i_74239360(.A(nbus_140[23]), .B(n_61689), .C(n_27920), .Z(n_283074182
		));
	notech_nand2 i_73539365(.A(readio_data[23]), .B(n_30272), .Z(n_283574187
		));
	notech_or4 i_73239368(.A(n_61889), .B(n_25467), .C(n_61718), .D(nbus_11271
		[7]), .Z(n_283874190));
	notech_nao3 i_72939371(.A(nbus_138[23]), .B(n_61689), .C(n_27919), .Z(n_284174193
		));
	notech_nao3 i_77239331(.A(cr2_reg[24]), .B(n_32268), .C(n_58506), .Z(n_284274194
		));
	notech_nao3 i_77139332(.A(n_318760815), .B(cr3[24]), .C(n_58506), .Z(n_284574197
		));
	notech_nand2 i_76839335(.A(\nbus_14542[24] ), .B(n_23351), .Z(n_284874200
		));
	notech_nao3 i_76539338(.A(nbus_140[24]), .B(n_61688), .C(n_27920), .Z(n_285174203
		));
	notech_or4 i_76039343(.A(n_30926), .B(n_30691), .C(n_19548), .D(n_32475)
		, .Z(n_285674208));
	notech_or4 i_75739346(.A(n_61718), .B(n_61889), .C(n_25467), .D(nbus_11271
		[8]), .Z(n_285974211));
	notech_nao3 i_75439349(.A(nbus_138[24]), .B(n_61688), .C(n_27919), .Z(n_286274214
		));
	notech_nao3 i_79539309(.A(cr2_reg[25]), .B(n_32268), .C(n_58501), .Z(n_286374215
		));
	notech_nao3 i_79439310(.A(n_318760815), .B(cr3[25]), .C(n_58501), .Z(n_286674218
		));
	notech_nao3 i_79139313(.A(\nbus_14542[25] ), .B(n_32249), .C(n_58501), .Z
		(n_286974221));
	notech_nao3 i_78839316(.A(nbus_140[25]), .B(n_61688), .C(n_27920), .Z(n_287274224
		));
	notech_or4 i_78339321(.A(n_30926), .B(n_30691), .C(n_19548), .D(n_32476)
		, .Z(n_287774229));
	notech_or4 i_77939324(.A(n_61718), .B(n_61885), .C(n_58541), .D(nbus_11271
		[9]), .Z(n_288074232));
	notech_nao3 i_77639327(.A(nbus_138[25]), .B(n_61688), .C(n_27919), .Z(n_288374235
		));
	notech_nao3 i_81839287(.A(cr2_reg[26]), .B(n_32268), .C(n_58501), .Z(n_288474236
		));
	notech_nao3 i_81739288(.A(n_318760815), .B(cr3[26]), .C(n_58501), .Z(n_288774239
		));
	notech_nand2 i_81439291(.A(\nbus_14542[26] ), .B(n_23351), .Z(n_289074242
		));
	notech_nao3 i_81139294(.A(nbus_140[26]), .B(n_61688), .C(n_27920), .Z(n_289374245
		));
	notech_or4 i_80639299(.A(n_30926), .B(n_30691), .C(n_19548), .D(n_32478)
		, .Z(n_289874250));
	notech_or4 i_80239302(.A(n_61723), .B(n_61885), .C(n_58541), .D(nbus_11271
		[10]), .Z(n_290174253));
	notech_nao3 i_79939305(.A(nbus_138[26]), .B(n_61689), .C(n_27919), .Z(n_290474256
		));
	notech_nao3 i_84039265(.A(cr2_reg[27]), .B(n_32268), .C(n_58501), .Z(n_290574257
		));
	notech_nao3 i_83939266(.A(n_318760815), .B(cr3[27]), .C(n_58501), .Z(n_290874260
		));
	notech_nand2 i_83639269(.A(\nbus_14542[27] ), .B(n_23351), .Z(n_291174263
		));
	notech_nao3 i_83339272(.A(nbus_140[27]), .B(n_61689), .C(n_27920), .Z(n_291474266
		));
	notech_or4 i_82839277(.A(n_30926), .B(n_30691), .C(n_19548), .D(n_32480)
		, .Z(n_291974271));
	notech_or4 i_82539280(.A(n_61723), .B(n_61885), .C(n_58541), .D(nbus_11271
		[11]), .Z(n_292274274));
	notech_nao3 i_82239283(.A(nbus_138[27]), .B(n_61689), .C(n_58523), .Z(n_292574277
		));
	notech_nao3 i_86239243(.A(cr2_reg[28]), .B(n_32268), .C(n_58501), .Z(n_292674278
		));
	notech_nao3 i_86139244(.A(n_318760815), .B(cr3[28]), .C(n_58501), .Z(n_292974281
		));
	notech_nand2 i_85839247(.A(\nbus_14542[28] ), .B(n_23351), .Z(n_293274284
		));
	notech_nao3 i_85539250(.A(opa_0[28]), .B(n_61689), .C(n_27922), .Z(n_293574287
		));
	notech_or2 i_85039255(.A(n_23345), .B(\nbus_11290[28] ), .Z(n_294074292)
		);
	notech_or4 i_84739258(.A(n_61723), .B(n_61885), .C(n_58541), .D(nbus_11271
		[12]), .Z(n_294374295));
	notech_nao3 i_84439261(.A(nbus_138[28]), .B(n_61689), .C(n_58523), .Z(n_294674298
		));
	notech_nao3 i_88539221(.A(cr2_reg[29]), .B(n_32268), .C(n_58501), .Z(n_294774299
		));
	notech_nao3 i_88439222(.A(n_318760815), .B(cr3[29]), .C(n_58501), .Z(n_295074302
		));
	notech_nand2 i_88139225(.A(\nbus_14542[29] ), .B(n_23351), .Z(n_295374305
		));
	notech_nao3 i_87839228(.A(nbus_140[29]), .B(n_61684), .C(n_27920), .Z(n_295674308
		));
	notech_nand2 i_87339233(.A(readio_data[29]), .B(n_30272), .Z(n_296174313
		));
	notech_or4 i_87039236(.A(n_61718), .B(n_61885), .C(n_58541), .D(nbus_11271
		[13]), .Z(n_296474316));
	notech_nao3 i_86639239(.A(nbus_138[29]), .B(n_61679), .C(n_58523), .Z(n_296774319
		));
	notech_nao3 i_90739199(.A(cr2_reg[30]), .B(n_58601), .C(n_58501), .Z(n_296874320
		));
	notech_nao3 i_90639200(.A(n_318760815), .B(cr3[30]), .C(n_58501), .Z(n_297174323
		));
	notech_nand2 i_90339203(.A(\nbus_14542[30] ), .B(n_23351), .Z(n_297474326
		));
	notech_nao3 i_90039206(.A(nbus_140[30]), .B(n_61679), .C(n_27920), .Z(n_297774329
		));
	notech_nand2 i_89539211(.A(readio_data[30]), .B(n_30272), .Z(n_298274334
		));
	notech_or4 i_89239214(.A(n_61718), .B(n_61885), .C(n_58541), .D(nbus_11271
		[14]), .Z(n_298574337));
	notech_nao3 i_88939217(.A(nbus_138[30]), .B(n_61679), .C(n_58523), .Z(n_298874340
		));
	notech_nao3 i_92939177(.A(cr2_reg[31]), .B(n_58601), .C(n_58501), .Z(n_298974341
		));
	notech_nao3 i_92839178(.A(n_318760815), .B(cr3[31]), .C(n_58501), .Z(n_299274344
		));
	notech_nand2 i_92539181(.A(\nbus_14542[31] ), .B(n_23351), .Z(n_299574347
		));
	notech_nao3 i_92239184(.A(nbus_140[31]), .B(n_61675), .C(n_27920), .Z(n_299874350
		));
	notech_nand2 i_91739189(.A(readio_data[31]), .B(n_30272), .Z(n_300374355
		));
	notech_or4 i_91439192(.A(n_61885), .B(n_58541), .C(n_61723), .D(nbus_11271
		[15]), .Z(n_300674358));
	notech_nao3 i_91139195(.A(nbus_138[31]), .B(n_61675), .C(n_58523), .Z(n_300974361
		));
	notech_or4 i_211438034(.A(n_61917), .B(n_61901), .C(n_61885), .D(nbus_11273
		[7]), .Z(n_301074362));
	notech_or4 i_145740077(.A(n_25680), .B(n_63764), .C(n_61958), .D(n_61625
		), .Z(n_301274364));
	notech_or4 i_145640078(.A(n_25680), .B(\opcode[1] ), .C(n_61935), .D(n_61628
		), .Z(n_301374365));
	notech_and2 i_188938251(.A(n_23379), .B(n_301374365), .Z(n_301474366));
	notech_and3 i_194540063(.A(n_23379), .B(n_301374365), .C(n_301274364), .Z
		(n_301574367));
	notech_or4 i_151240074(.A(n_25680), .B(\opcode[1] ), .C(n_63764), .D(n_61628
		), .Z(n_301874370));
	notech_ao4 i_188438256(.A(n_301874370), .B(n_31507), .C(n_224073608), .D
		(\nbus_11283[31] ), .Z(n_301974371));
	notech_or4 i_69740084(.A(n_32396), .B(n_28008), .C(n_60157), .D(n_61625)
		, .Z(n_302174373));
	notech_ao4 i_188238258(.A(n_218373551), .B(n_33414), .C(n_302174373), .D
		(n_32803), .Z(n_302274374));
	notech_and4 i_188638254(.A(n_302274374), .B(n_301974371), .C(n_300674358
		), .D(n_300974361), .Z(n_302474376));
	notech_ao4 i_187938261(.A(n_23334), .B(nbus_11271[31]), .C(n_23379), .D(n_32059
		), .Z(n_302574377));
	notech_ao4 i_187838262(.A(n_30612), .B(n_33413), .C(n_23329), .D(n_32489
		), .Z(n_302774379));
	notech_and4 i_188738253(.A(n_302574377), .B(n_302774379), .C(n_302474376
		), .D(n_300374355), .Z(n_302974381));
	notech_ao4 i_187338266(.A(n_32374), .B(n_30688), .C(n_27814), .D(n_32450
		), .Z(n_303074382));
	notech_ao4 i_187038268(.A(n_23345), .B(\nbus_11290[31] ), .C(n_23353), .D
		(n_31199), .Z(n_303274384));
	notech_and4 i_187538264(.A(n_303274384), .B(n_303074382), .C(n_299574347
		), .D(n_299874350), .Z(n_303474386));
	notech_ao4 i_186738271(.A(n_1828), .B(n_33206), .C(n_1827), .D(n_32421),
		 .Z(n_303574387));
	notech_and4 i_186938269(.A(n_317751253), .B(n_303574387), .C(n_298974341
		), .D(n_299274344), .Z(n_303874390));
	notech_ao4 i_186238276(.A(n_301874370), .B(n_31506), .C(\nbus_11283[30] 
		), .D(n_223873606), .Z(n_304074392));
	notech_ao4 i_186038278(.A(n_57978), .B(n_33412), .C(n_302174373), .D(n_32802
		), .Z(n_304274394));
	notech_and4 i_186438274(.A(n_304274394), .B(n_304074392), .C(n_298574337
		), .D(n_298874340), .Z(n_304474396));
	notech_ao4 i_185738281(.A(n_23334), .B(nbus_11271[30]), .C(n_23379), .D(n_32058
		), .Z(n_304574397));
	notech_ao4 i_185638282(.A(n_30612), .B(n_33411), .C(n_23329), .D(n_32488
		), .Z(n_304774399));
	notech_and4 i_186538273(.A(n_304574397), .B(n_304774399), .C(n_304474396
		), .D(n_298274334), .Z(n_304974401));
	notech_ao4 i_185238286(.A(n_30688), .B(n_32373), .C(n_27814), .D(n_32449
		), .Z(n_305074402));
	notech_ao4 i_185038288(.A(n_23345), .B(\nbus_11290[30] ), .C(n_23353), .D
		(n_31198), .Z(n_305274404));
	notech_and4 i_185438284(.A(n_305274404), .B(n_305074402), .C(n_297474326
		), .D(n_297774329), .Z(n_305474406));
	notech_ao4 i_184738291(.A(n_1828), .B(n_33194), .C(n_1827), .D(n_32420),
		 .Z(n_305574407));
	notech_and4 i_184938289(.A(n_317751253), .B(n_305574407), .C(n_296874320
		), .D(n_297174323), .Z(n_305874410));
	notech_ao4 i_184238296(.A(n_301874370), .B(n_31505), .C(n_223673604), .D
		(\nbus_11283[29] ), .Z(n_306074412));
	notech_ao4 i_184038298(.A(n_218373551), .B(n_33410), .C(n_302174373), .D
		(n_32801), .Z(n_306274414));
	notech_and4 i_184438294(.A(n_306274414), .B(n_306074412), .C(n_296474316
		), .D(n_296774319), .Z(n_306474416));
	notech_ao4 i_183738301(.A(n_23334), .B(nbus_11271[29]), .C(n_23379), .D(n_32057
		), .Z(n_306574417));
	notech_ao4 i_183638302(.A(n_30612), .B(n_33409), .C(n_23329), .D(n_32483
		), .Z(n_306774419));
	notech_and4 i_184538293(.A(n_306574417), .B(n_306774419), .C(n_306474416
		), .D(n_296174313), .Z(n_306974421));
	notech_ao4 i_183238306(.A(n_30688), .B(n_32371), .C(n_27814), .D(n_32448
		), .Z(n_307074422));
	notech_ao4 i_183038308(.A(n_23345), .B(\nbus_11290[29] ), .C(n_23353), .D
		(n_31197), .Z(n_307274424));
	notech_and4 i_183438304(.A(n_307274424), .B(n_307074422), .C(n_295374305
		), .D(n_295674308), .Z(n_307474426));
	notech_ao4 i_182638311(.A(n_1828), .B(n_33197), .C(n_1827), .D(n_32419),
		 .Z(n_307574427));
	notech_and4 i_182938309(.A(n_317751253), .B(n_307574427), .C(n_294774299
		), .D(n_295074302), .Z(n_307874430));
	notech_ao4 i_182038316(.A(n_301874370), .B(n_31504), .C(n_223473602), .D
		(\nbus_11283[28] ), .Z(n_308074432));
	notech_ao4 i_181838318(.A(n_218373551), .B(n_33408), .C(n_302174373), .D
		(n_32800), .Z(n_308274434));
	notech_and4 i_182338314(.A(n_308274434), .B(n_308074432), .C(n_294374295
		), .D(n_294674298), .Z(n_308474436));
	notech_ao4 i_181538321(.A(n_23334), .B(nbus_11271[28]), .C(n_23379), .D(n_32056
		), .Z(n_308574437));
	notech_ao4 i_181438322(.A(n_23329), .B(n_32482), .C(n_1826), .D(n_32528)
		, .Z(n_308774439));
	notech_and4 i_182438313(.A(n_308574437), .B(n_308774439), .C(n_308474436
		), .D(n_294074292), .Z(n_308974441));
	notech_ao4 i_181038326(.A(n_27814), .B(n_32447), .C(n_30612), .D(n_33407
		), .Z(n_309074442));
	notech_ao4 i_180838328(.A(n_23353), .B(n_31196), .C(n_23341), .D(n_32751
		), .Z(n_309274444));
	notech_and4 i_181238324(.A(n_309274444), .B(n_309074442), .C(n_293274284
		), .D(n_293574287), .Z(n_309474446));
	notech_ao4 i_180538331(.A(n_1828), .B(n_33196), .C(n_1827), .D(n_32418),
		 .Z(n_309574447));
	notech_and4 i_180738329(.A(n_317751253), .B(n_309574447), .C(n_292674278
		), .D(n_292974281), .Z(n_309874450));
	notech_ao4 i_179938336(.A(n_301874370), .B(n_31503), .C(\nbus_11283[27] 
		), .D(n_223273600), .Z(n_310074452));
	notech_ao4 i_179738338(.A(n_218373551), .B(n_33406), .C(n_302174373), .D
		(n_32799), .Z(n_310274454));
	notech_and4 i_180138334(.A(n_310274454), .B(n_310074452), .C(n_292274274
		), .D(n_292574277), .Z(n_310474456));
	notech_ao4 i_179438341(.A(n_1826), .B(n_32527), .C(n_23379), .D(n_32055)
		, .Z(n_310574457));
	notech_ao4 i_179338342(.A(n_23334), .B(nbus_11271[27]), .C(n_30612), .D(n_33405
		), .Z(n_310774459));
	notech_and4 i_180238333(.A(n_310574457), .B(n_310774459), .C(n_310474456
		), .D(n_291974271), .Z(n_310974461));
	notech_ao4 i_178938346(.A(n_30688), .B(n_32370), .C(n_27814), .D(n_32446
		), .Z(n_311074462));
	notech_ao4 i_178738348(.A(n_23345), .B(\nbus_11290[27] ), .C(n_23353), .D
		(n_31195), .Z(n_311274464));
	notech_and4 i_179138344(.A(n_311274464), .B(n_311074462), .C(n_291174263
		), .D(n_291474266), .Z(n_311474466));
	notech_ao4 i_178438351(.A(n_1828), .B(n_33195), .C(n_1827), .D(n_32417),
		 .Z(n_311574467));
	notech_and4 i_178638349(.A(n_317751253), .B(n_311574467), .C(n_290574257
		), .D(n_290874260), .Z(n_311874470));
	notech_ao4 i_177838356(.A(n_301874370), .B(n_31502), .C(\nbus_11283[26] 
		), .D(n_223073598), .Z(n_312074472));
	notech_ao4 i_177638358(.A(n_57978), .B(n_33404), .C(n_302174373), .D(n_32798
		), .Z(n_312274474));
	notech_and4 i_178038354(.A(n_312274474), .B(n_312074472), .C(n_290174253
		), .D(n_290474256), .Z(n_312474476));
	notech_ao4 i_177338361(.A(n_1826), .B(n_32526), .C(n_23379), .D(n_32054)
		, .Z(n_312574477));
	notech_ao4 i_177238362(.A(n_23334), .B(nbus_11271[26]), .C(n_30612), .D(n_33403
		), .Z(n_312774479));
	notech_and4 i_178138353(.A(n_312574477), .B(n_312774479), .C(n_312474476
		), .D(n_289874250), .Z(n_312974481));
	notech_ao4 i_176638366(.A(n_30688), .B(n_32369), .C(n_27814), .D(n_32445
		), .Z(n_313074482));
	notech_ao4 i_176438368(.A(n_23345), .B(\nbus_11290[26] ), .C(n_23353), .D
		(n_31194), .Z(n_313274484));
	notech_and4 i_176938364(.A(n_313274484), .B(n_313074482), .C(n_289074242
		), .D(n_289374245), .Z(n_313474486));
	notech_ao4 i_176138371(.A(n_1828), .B(n_33198), .C(n_1827), .D(n_32416),
		 .Z(n_313574487));
	notech_and4 i_176338369(.A(n_317751253), .B(n_313574487), .C(n_288474236
		), .D(n_288774239), .Z(n_313874490));
	notech_ao4 i_175638376(.A(n_301874370), .B(n_31501), .C(\nbus_11283[25] 
		), .D(n_222873596), .Z(n_314074492));
	notech_ao4 i_175438378(.A(n_57978), .B(n_33402), .C(n_302174373), .D(n_32797
		), .Z(n_314274494));
	notech_and4 i_175838374(.A(n_314274494), .B(n_314074492), .C(n_288074232
		), .D(n_288374235), .Z(n_314474496));
	notech_ao4 i_175138381(.A(n_1826), .B(n_32525), .C(n_23379), .D(n_32053)
		, .Z(n_314574497));
	notech_ao4 i_175038382(.A(n_23334), .B(nbus_11271[25]), .C(n_30612), .D(n_33401
		), .Z(n_314774499));
	notech_and4 i_175938373(.A(n_314574497), .B(n_314774499), .C(n_314474496
		), .D(n_287774229), .Z(n_314974501));
	notech_ao4 i_174638386(.A(n_30688), .B(n_32367), .C(n_27814), .D(n_32444
		), .Z(n_315074502));
	notech_ao4 i_174438388(.A(n_23345), .B(\nbus_11290[25] ), .C(n_23353), .D
		(n_31193), .Z(n_315374504));
	notech_and4 i_174838384(.A(n_315374504), .B(n_315074502), .C(n_286974221
		), .D(n_287274224), .Z(n_315574506));
	notech_ao4 i_174138391(.A(n_1828), .B(n_33172), .C(n_1827), .D(n_32415),
		 .Z(n_315674507));
	notech_and4 i_174338389(.A(n_317751253), .B(n_315674507), .C(n_286374215
		), .D(n_286674218), .Z(n_316074510));
	notech_ao4 i_173638396(.A(n_301874370), .B(n_31500), .C(\nbus_11283[24] 
		), .D(n_222673594), .Z(n_316274512));
	notech_ao4 i_173438398(.A(n_57978), .B(n_33400), .C(n_302174373), .D(n_32796
		), .Z(n_316474514));
	notech_and4 i_173838394(.A(n_316474514), .B(n_316274512), .C(n_285974211
		), .D(n_286274214), .Z(n_316674516));
	notech_ao4 i_173138401(.A(n_1826), .B(n_32524), .C(n_23379), .D(n_32052)
		, .Z(n_316774517));
	notech_ao4 i_173038402(.A(n_23334), .B(nbus_11271[24]), .C(n_30612), .D(n_33399
		), .Z(n_316974519));
	notech_and4 i_173938393(.A(n_316774517), .B(n_316974519), .C(n_316674516
		), .D(n_285674208), .Z(n_317174521));
	notech_ao4 i_172638406(.A(n_30688), .B(n_32366), .C(n_27814), .D(n_32443
		), .Z(n_317274522));
	notech_ao4 i_172438408(.A(n_23345), .B(\nbus_11290[24] ), .C(n_23353), .D
		(n_31192), .Z(n_317474524));
	notech_and4 i_172838404(.A(n_317474524), .B(n_317274522), .C(n_284874200
		), .D(n_285174203), .Z(n_317674526));
	notech_ao4 i_172138411(.A(n_1828), .B(n_33171), .C(n_1827), .D(n_32414),
		 .Z(n_317774527));
	notech_and4 i_172338409(.A(n_317751253), .B(n_317774527), .C(n_284274194
		), .D(n_284574197), .Z(n_318074530));
	notech_ao4 i_171638416(.A(n_301874370), .B(n_31499), .C(n_222473592), .D
		(n_58420), .Z(n_318274532));
	notech_ao4 i_171438418(.A(n_57978), .B(n_33398), .C(n_302174373), .D(n_32795
		), .Z(n_318474534));
	notech_and4 i_171838414(.A(n_318474534), .B(n_318274532), .C(n_283874190
		), .D(n_284174193), .Z(n_318674536));
	notech_ao4 i_171138421(.A(n_23334), .B(nbus_11271[23]), .C(n_32051), .D(n_23379
		), .Z(n_318774537));
	notech_ao4 i_171038422(.A(n_30612), .B(n_33397), .C(n_23329), .D(n_32474
		), .Z(n_318974539));
	notech_and4 i_171938413(.A(n_318774537), .B(n_318974539), .C(n_318674536
		), .D(n_283574187), .Z(n_319174541));
	notech_ao4 i_170638426(.A(n_30688), .B(n_32365), .C(n_27814), .D(n_32442
		), .Z(n_319274542));
	notech_ao4 i_170438428(.A(n_23345), .B(n_58902), .C(n_23353), .D(n_31191
		), .Z(n_319474544));
	notech_and4 i_170838424(.A(n_319474544), .B(n_319274542), .C(n_282774179
		), .D(n_283074182), .Z(n_319774546));
	notech_ao4 i_170138431(.A(n_1828), .B(n_33170), .C(n_1827), .D(n_32413),
		 .Z(n_319874547));
	notech_and4 i_170338429(.A(n_317751253), .B(n_319874547), .C(n_282174173
		), .D(n_282474176), .Z(n_320274550));
	notech_ao4 i_169638436(.A(n_301874370), .B(n_31496), .C(n_222273590), .D
		(\nbus_11283[22] ), .Z(n_320474552));
	notech_ao4 i_169438438(.A(n_57978), .B(n_33396), .C(n_302174373), .D(n_32794
		), .Z(n_320674554));
	notech_and4 i_169838434(.A(n_320674554), .B(n_320474552), .C(n_281774169
		), .D(n_282074172), .Z(n_320874556));
	notech_ao4 i_169138441(.A(n_1826), .B(n_32523), .C(n_23379), .D(n_32050)
		, .Z(n_320974557));
	notech_ao4 i_169038442(.A(n_23334), .B(nbus_11271[22]), .C(n_30612), .D(n_33395
		), .Z(n_321174559));
	notech_and4 i_169938433(.A(n_320974557), .B(n_321174559), .C(n_320874556
		), .D(n_281474166), .Z(n_321374561));
	notech_ao4 i_168638446(.A(n_30688), .B(n_32364), .C(n_27814), .D(n_32441
		), .Z(n_321474562));
	notech_ao4 i_168438448(.A(n_23345), .B(\nbus_11290[22] ), .C(n_23353), .D
		(n_31190), .Z(n_321674564));
	notech_and4 i_168838444(.A(n_321674564), .B(n_321474562), .C(n_280674158
		), .D(n_280974161), .Z(n_321874566));
	notech_ao4 i_168138451(.A(n_1828), .B(n_33284), .C(n_1827), .D(n_32412),
		 .Z(n_321974567));
	notech_and4 i_168338449(.A(n_321974567), .B(n_280074152), .C(n_280374155
		), .D(n_317751253), .Z(n_322274570));
	notech_ao4 i_167638456(.A(n_301874370), .B(n_31494), .C(n_222073588), .D
		(n_58402), .Z(n_322474572));
	notech_ao4 i_167438458(.A(n_57978), .B(n_33394), .C(n_302174373), .D(n_32793
		), .Z(n_322774574));
	notech_and4 i_167838454(.A(n_322774574), .B(n_322474572), .C(n_279674148
		), .D(n_279974151), .Z(n_322974576));
	notech_ao4 i_167138461(.A(n_1826), .B(n_32519), .C(n_23379), .D(n_32049)
		, .Z(n_323074577));
	notech_ao4 i_167038462(.A(n_23334), .B(nbus_11271[21]), .C(n_30612), .D(n_33393
		), .Z(n_323374579));
	notech_and3 i_167338459(.A(n_323074577), .B(n_323374579), .C(n_279374145
		), .Z(n_323474580));
	notech_ao4 i_166538466(.A(n_30688), .B(n_32363), .C(n_27814), .D(n_32440
		), .Z(n_323674582));
	notech_ao4 i_166238468(.A(n_23345), .B(n_58884), .C(n_23353), .D(n_31189
		), .Z(n_323874584));
	notech_and4 i_166738464(.A(n_323874584), .B(n_323674582), .C(n_278574137
		), .D(n_278874140), .Z(n_324074586));
	notech_ao4 i_165938471(.A(n_57867), .B(n_33288), .C(n_1827), .D(n_32411)
		, .Z(n_324174587));
	notech_ao4 i_165838472(.A(n_1834), .B(n_301074362), .C(n_23383), .D(n_31216
		), .Z(n_324374589));
	notech_and4 i_166838463(.A(n_324174587), .B(n_324374589), .C(n_324074586
		), .D(n_278274134), .Z(n_324574591));
	notech_ao4 i_165138476(.A(n_301874370), .B(n_31493), .C(n_221873586), .D
		(n_58393), .Z(n_324674592));
	notech_ao4 i_164938478(.A(n_218373551), .B(n_33392), .C(n_302174373), .D
		(n_32792), .Z(n_324874594));
	notech_and4 i_165338474(.A(n_324874594), .B(n_324674592), .C(n_277574127
		), .D(n_277874130), .Z(n_325074596));
	notech_ao4 i_164638481(.A(n_1826), .B(n_32518), .C(n_23379), .D(n_32048)
		, .Z(n_325174597));
	notech_ao4 i_164538482(.A(n_23334), .B(nbus_11271[20]), .C(n_30612), .D(n_33391
		), .Z(n_325374599));
	notech_and4 i_165538473(.A(n_325174597), .B(n_325374599), .C(n_325074596
		), .D(n_277274124), .Z(n_325574601));
	notech_ao4 i_164138486(.A(n_30688), .B(n_32362), .C(n_27814), .D(n_32439
		), .Z(n_325674602));
	notech_ao4 i_163938488(.A(n_23345), .B(n_58857), .C(n_23353), .D(n_31188
		), .Z(n_325874604));
	notech_and4 i_164338484(.A(n_325874604), .B(n_325674602), .C(n_276474116
		), .D(n_276774119), .Z(n_326074606));
	notech_ao4 i_163638491(.A(n_57867), .B(n_33292), .C(n_1827), .D(n_32410)
		, .Z(n_326174607));
	notech_and4 i_163838489(.A(n_317751253), .B(n_326174607), .C(n_275874110
		), .D(n_276174113), .Z(n_326474610));
	notech_ao4 i_163138496(.A(n_57928), .B(n_31492), .C(n_221673584), .D(\nbus_11283[19] 
		), .Z(n_326674612));
	notech_ao4 i_162938498(.A(n_218373551), .B(n_33390), .C(n_302174373), .D
		(n_32791), .Z(n_326974614));
	notech_and4 i_163338494(.A(n_326974614), .B(n_326674612), .C(n_275474106
		), .D(n_275774109), .Z(n_327274616));
	notech_ao4 i_162538501(.A(n_1826), .B(n_32517), .C(n_23379), .D(n_32047)
		, .Z(n_327374617));
	notech_ao4 i_162438502(.A(n_23334), .B(nbus_11271[19]), .C(n_30612), .D(n_33389
		), .Z(n_327574619));
	notech_and4 i_163438493(.A(n_327374617), .B(n_327574619), .C(n_327274616
		), .D(n_275174103), .Z(n_327774621));
	notech_ao4 i_162038506(.A(n_30688), .B(n_32360), .C(n_27814), .D(n_32438
		), .Z(n_327874622));
	notech_ao4 i_161738508(.A(n_58512), .B(\nbus_11290[19] ), .C(n_23353), .D
		(n_31187), .Z(n_328074624));
	notech_and4 i_162238504(.A(n_328074624), .B(n_327874622), .C(n_274374095
		), .D(n_274674098), .Z(n_328274626));
	notech_ao4 i_161438511(.A(n_57867), .B(n_33202), .C(n_1827), .D(n_32409)
		, .Z(n_328374627));
	notech_and4 i_161638509(.A(n_317751253), .B(n_328374627), .C(n_273774089
		), .D(n_274074092), .Z(n_328674630));
	notech_ao4 i_160938516(.A(n_57928), .B(n_31491), .C(n_221473582), .D(\nbus_11283[18] 
		), .Z(n_328874632));
	notech_ao4 i_160738518(.A(n_218373551), .B(n_33388), .C(n_302174373), .D
		(n_32790), .Z(n_329074634));
	notech_and4 i_161138514(.A(n_329074634), .B(n_328874632), .C(n_273374085
		), .D(n_273674088), .Z(n_329274636));
	notech_ao4 i_160438521(.A(n_1826), .B(n_32516), .C(n_23379), .D(n_32046)
		, .Z(n_329374637));
	notech_ao4 i_160338522(.A(n_23334), .B(nbus_11271[18]), .C(n_30612), .D(n_33387
		), .Z(n_329574639));
	notech_and4 i_161238513(.A(n_329374637), .B(n_329574639), .C(n_329274636
		), .D(n_272674082), .Z(n_329774641));
	notech_ao4 i_159938526(.A(n_30688), .B(n_32359), .C(n_27814), .D(n_32437
		), .Z(n_329874642));
	notech_ao4 i_159738528(.A(n_58512), .B(\nbus_11290[18] ), .C(n_23353), .D
		(n_31186), .Z(n_330074644));
	notech_and4 i_160138524(.A(n_330074644), .B(n_329874642), .C(n_271874074
		), .D(n_272174077), .Z(n_330274646));
	notech_ao4 i_159438531(.A(n_57867), .B(n_33201), .C(n_1827), .D(n_32408)
		, .Z(n_330374647));
	notech_and4 i_159638529(.A(n_57878), .B(n_330374647), .C(n_271074068), .D
		(n_271574071), .Z(n_330674650));
	notech_ao4 i_158938536(.A(n_57928), .B(n_31490), .C(n_221273580), .D(\nbus_11283[17] 
		), .Z(n_330874652));
	notech_ao4 i_158738538(.A(n_218373551), .B(n_33386), .C(n_302174373), .D
		(n_32788), .Z(n_331074654));
	notech_and4 i_159138534(.A(n_331074654), .B(n_330874652), .C(n_270674064
		), .D(n_270974067), .Z(n_331274656));
	notech_ao4 i_158438541(.A(n_1826), .B(n_32515), .C(n_23379), .D(n_32045)
		, .Z(n_331374657));
	notech_ao4 i_158338542(.A(n_23334), .B(nbus_11271[17]), .C(n_30612), .D(n_33385
		), .Z(n_331574659));
	notech_and4 i_159238533(.A(n_331374657), .B(n_331574659), .C(n_331274656
		), .D(n_270374061), .Z(n_331774661));
	notech_ao4 i_157938546(.A(n_30688), .B(n_32358), .C(n_27814), .D(n_32436
		), .Z(n_331874662));
	notech_ao4 i_157738548(.A(n_58512), .B(\nbus_11290[17] ), .C(n_58492), .D
		(n_31185), .Z(n_332074664));
	notech_and4 i_158138544(.A(n_332074664), .B(n_331874662), .C(n_269574053
		), .D(n_269874056), .Z(n_332474666));
	notech_ao4 i_157438551(.A(n_57867), .B(n_33200), .C(n_1827), .D(n_32406)
		, .Z(n_332574667));
	notech_and4 i_157638549(.A(n_57878), .B(n_332574667), .C(n_268774047), .D
		(n_269274050), .Z(n_332874670));
	notech_ao4 i_156938556(.A(n_57928), .B(n_31489), .C(n_221073578), .D(\nbus_11283[16] 
		), .Z(n_333074672));
	notech_ao4 i_156738558(.A(n_218373551), .B(n_33384), .C(n_302174373), .D
		(n_32787), .Z(n_333274674));
	notech_and4 i_157138554(.A(n_333274674), .B(n_333074672), .C(n_267574043
		), .D(n_267874046), .Z(n_333474676));
	notech_ao4 i_156438561(.A(n_1826), .B(n_32513), .C(n_57998), .D(n_32044)
		, .Z(n_333574677));
	notech_ao4 i_156338562(.A(n_23334), .B(nbus_11271[16]), .C(n_30612), .D(n_33383
		), .Z(n_333774679));
	notech_and3 i_156638559(.A(n_333574677), .B(n_333774679), .C(n_267274040
		), .Z(n_333874680));
	notech_ao4 i_155938566(.A(n_30688), .B(n_32357), .C(n_58215), .D(n_32435
		), .Z(n_334074682));
	notech_ao4 i_155638568(.A(n_58512), .B(\nbus_11290[16] ), .C(n_58492), .D
		(n_31184), .Z(n_334274684));
	notech_and4 i_156138564(.A(n_334274684), .B(n_334074682), .C(n_266474032
		), .D(n_266774035), .Z(n_334474686));
	notech_ao4 i_155238571(.A(n_57867), .B(n_33199), .C(n_1827), .D(n_32405)
		, .Z(n_334574687));
	notech_ao4 i_155138572(.A(n_1834), .B(n_301074362), .C(n_23383), .D(n_31215
		), .Z(n_334774689));
	notech_and4 i_156238563(.A(n_334574687), .B(n_334774689), .C(n_334474686
		), .D(n_266174029), .Z(n_334974691));
	notech_or4 i_155440072(.A(n_25485), .B(\opcode[1] ), .C(n_63764), .D(n_61625
		), .Z(n_335174693));
	notech_ao4 i_154638577(.A(n_335174693), .B(\nbus_11283[31] ), .C(n_220773575
		), .D(nbus_11273[15]), .Z(n_335274694));
	notech_nao3 i_154440073(.A(n_27843), .B(n_61679), .C(n_30696), .Z(n_335374695
		));
	notech_ao4 i_154538578(.A(n_57928), .B(n_31488), .C(n_335374695), .D(n_32852
		), .Z(n_335474696));
	notech_ao4 i_154238580(.A(n_301374365), .B(\nbus_11290[7] ), .C(n_301274364
		), .D(n_31480), .Z(n_335674698));
	notech_ao4 i_154138581(.A(n_58007), .B(nbus_11271[15]), .C(n_57998), .D(n_32043
		), .Z(n_335774699));
	notech_and4 i_154838575(.A(n_335774699), .B(n_335674698), .C(n_335474696
		), .D(n_335274694), .Z(n_335974701));
	notech_ao4 i_153838584(.A(n_58512), .B(\nbus_11290[15] ), .C(n_57917), .D
		(nbus_11273[7]), .Z(n_336074702));
	notech_ao4 i_153738585(.A(n_23329), .B(n_32466), .C(n_1826), .D(n_32512)
		, .Z(n_336174703));
	notech_ao4 i_153538587(.A(n_58215), .B(n_32434), .C(n_57987), .D(n_33382
		), .Z(n_336374705));
	notech_and4 i_154038582(.A(n_336374705), .B(n_336174703), .C(n_336074702
		), .D(n_264574013), .Z(n_336574707));
	notech_ao4 i_153038591(.A(n_30611), .B(n_31063), .C(n_22979), .D(\nbus_11290[31] 
		), .Z(n_336774709));
	notech_ao4 i_152938592(.A(n_57867), .B(n_33248), .C(n_57745), .D(n_32403
		), .Z(n_336874710));
	notech_ao4 i_152738594(.A(n_23383), .B(n_31214), .C(n_23359), .D(n_31610
		), .Z(n_337074712));
	notech_ao4 i_152638595(.A(n_22968), .B(n_32836), .C(n_22967), .D(n_32819
		), .Z(n_337174713));
	notech_and4 i_153338589(.A(n_337174713), .B(n_337074712), .C(n_336874710
		), .D(n_336774709), .Z(n_337374715));
	notech_ao4 i_152338598(.A(n_22976), .B(n_32356), .C(n_28089), .D(n_33381
		), .Z(n_337474716));
	notech_ao4 i_152238599(.A(n_22980), .B(n_32767), .C(n_22977), .D(n_32786
		), .Z(n_337574717));
	notech_ao4 i_152038601(.A(n_22985), .B(n_33380), .C(n_22984), .D(n_32750
		), .Z(n_337774719));
	notech_and4 i_152538596(.A(n_57878), .B(n_337774719), .C(n_337574717), .D
		(n_337474716), .Z(n_337974721));
	notech_ao4 i_151638605(.A(n_335174693), .B(\nbus_11283[30] ), .C(n_220573573
		), .D(nbus_11273[14]), .Z(n_338174723));
	notech_ao4 i_151538606(.A(n_57928), .B(n_31487), .C(n_335374695), .D(n_32851
		), .Z(n_338274724));
	notech_ao4 i_151338608(.A(n_301374365), .B(\nbus_11290[6] ), .C(n_301274364
		), .D(n_31479), .Z(n_338474726));
	notech_ao4 i_151138609(.A(n_57917), .B(nbus_11273[6]), .C(n_57998), .D(n_32042
		), .Z(n_338574727));
	notech_and4 i_151838603(.A(n_338574727), .B(n_338474726), .C(n_338274724
		), .D(n_338174723), .Z(n_338774729));
	notech_ao4 i_150838612(.A(n_1826), .B(n_32511), .C(n_58512), .D(\nbus_11290[14] 
		), .Z(n_338874730));
	notech_ao4 i_150738613(.A(n_57987), .B(n_33379), .C(n_23329), .D(n_32465
		), .Z(n_338974731));
	notech_ao4 i_150538615(.A(n_58215), .B(n_32433), .C(n_58007), .D(nbus_11271
		[14]), .Z(n_339174733));
	notech_and4 i_151038610(.A(n_339174733), .B(n_338974731), .C(n_338874730
		), .D(n_261673984), .Z(n_339374735));
	notech_ao4 i_150138619(.A(n_57745), .B(n_32399), .C(n_30611), .D(n_31062
		), .Z(n_339574737));
	notech_ao4 i_150038620(.A(n_23359), .B(n_31609), .C(n_57867), .D(n_33215
		), .Z(n_339674738));
	notech_ao4 i_149838622(.A(n_22979), .B(\nbus_11290[30] ), .C(n_23383), .D
		(n_31213), .Z(n_339874740));
	notech_ao4 i_149738623(.A(n_22968), .B(n_32835), .C(n_22967), .D(n_32818
		), .Z(n_339974741));
	notech_and4 i_150338617(.A(n_339974741), .B(n_339874740), .C(n_339674738
		), .D(n_339574737), .Z(n_340174743));
	notech_ao4 i_149438626(.A(n_22976), .B(n_32355), .C(n_28089), .D(n_33378
		), .Z(n_340274744));
	notech_ao4 i_149338627(.A(n_22980), .B(n_32766), .C(n_22977), .D(n_32784
		), .Z(n_340374745));
	notech_ao4 i_149138629(.A(n_22985), .B(n_33377), .C(n_22984), .D(n_32749
		), .Z(n_340574747));
	notech_and4 i_149638624(.A(n_57878), .B(n_340574747), .C(n_340374745), .D
		(n_340274744), .Z(n_340774749));
	notech_ao4 i_148538633(.A(n_335174693), .B(\nbus_11283[29] ), .C(n_220373571
		), .D(nbus_11273[13]), .Z(n_340974751));
	notech_ao4 i_148438634(.A(n_57928), .B(n_31486), .C(n_335374695), .D(n_32850
		), .Z(n_341074752));
	notech_ao4 i_148138636(.A(n_301374365), .B(\nbus_11290[5] ), .C(n_301274364
		), .D(n_31478), .Z(n_341274754));
	notech_ao4 i_148038637(.A(n_57917), .B(nbus_11273[5]), .C(n_57998), .D(n_32041
		), .Z(n_341374755));
	notech_and4 i_148838631(.A(n_341374755), .B(n_341274754), .C(n_341074752
		), .D(n_340974751), .Z(n_341574757));
	notech_ao4 i_147738640(.A(n_1826), .B(n_32510), .C(n_58512), .D(\nbus_11290[13] 
		), .Z(n_341674758));
	notech_ao4 i_147638641(.A(n_57987), .B(n_33376), .C(n_23329), .D(n_32464
		), .Z(n_341774759));
	notech_ao4 i_147438643(.A(n_58215), .B(n_32432), .C(nbus_11271[13]), .D(n_58007
		), .Z(n_341974761));
	notech_and4 i_147938638(.A(n_341974761), .B(n_341774759), .C(n_341674758
		), .D(n_258773955), .Z(n_342174763));
	notech_ao4 i_147038647(.A(n_57745), .B(n_32398), .C(n_30611), .D(n_31061
		), .Z(n_342374765));
	notech_ao4 i_146938648(.A(n_23359), .B(n_31608), .C(n_57867), .D(n_33213
		), .Z(n_342474766));
	notech_ao4 i_146738650(.A(n_22979), .B(\nbus_11290[29] ), .C(n_23383), .D
		(n_31212), .Z(n_342674768));
	notech_ao4 i_146638651(.A(n_22968), .B(n_32834), .C(n_22967), .D(n_32817
		), .Z(n_342774769));
	notech_and4 i_147238645(.A(n_342774769), .B(n_342674768), .C(n_342474766
		), .D(n_342374765), .Z(n_342974771));
	notech_ao4 i_146238654(.A(n_22976), .B(n_32354), .C(n_28089), .D(n_33375
		), .Z(n_343074772));
	notech_ao4 i_146138655(.A(n_22980), .B(n_32765), .C(n_22977), .D(n_32783
		), .Z(n_343174773));
	notech_ao4 i_145938657(.A(n_22985), .B(n_33374), .C(n_22984), .D(n_32748
		), .Z(n_343374775));
	notech_and4 i_146538652(.A(n_57878), .B(n_343374775), .C(n_343174773), .D
		(n_343074772), .Z(n_343574777));
	notech_ao4 i_145238661(.A(n_335174693), .B(\nbus_11283[28] ), .C(n_220173569
		), .D(nbus_11273[12]), .Z(n_343774779));
	notech_ao4 i_145138662(.A(n_57928), .B(n_31485), .C(n_335374695), .D(n_32849
		), .Z(n_343874780));
	notech_ao4 i_144938664(.A(n_301374365), .B(\nbus_11290[4] ), .C(n_301274364
		), .D(n_31477), .Z(n_344074782));
	notech_ao4 i_144838665(.A(n_57917), .B(nbus_11273[4]), .C(n_57998), .D(n_32040
		), .Z(n_344174783));
	notech_and4 i_145538659(.A(n_344174783), .B(n_344074782), .C(n_343874780
		), .D(n_343774779), .Z(n_344374785));
	notech_ao4 i_144538668(.A(n_58512), .B(\nbus_11290[12] ), .C(n_22979), .D
		(\nbus_11290[28] ), .Z(n_344474786));
	notech_ao4 i_144438669(.A(n_23329), .B(n_32463), .C(n_57887), .D(n_32509
		), .Z(n_344574787));
	notech_ao4 i_144238671(.A(n_58007), .B(nbus_11271[12]), .C(n_57987), .D(n_33373
		), .Z(n_344774789));
	notech_and4 i_144738666(.A(n_344774789), .B(n_344574787), .C(n_344474786
		), .D(n_255873926), .Z(n_344974791));
	notech_ao4 i_143838675(.A(n_30611), .B(n_31060), .C(n_58492), .D(n_31183
		), .Z(n_345174793));
	notech_ao4 i_143738676(.A(n_57867), .B(n_33250), .C(n_57745), .D(n_32395
		), .Z(n_345274794));
	notech_ao4 i_143538678(.A(n_23383), .B(n_31211), .C(n_23359), .D(n_31607
		), .Z(n_345474796));
	notech_ao4 i_143438679(.A(n_22968), .B(n_32833), .C(n_22967), .D(n_32816
		), .Z(n_345574797));
	notech_and4 i_144038673(.A(n_345574797), .B(n_345474796), .C(n_345274794
		), .D(n_345174793), .Z(n_345774799));
	notech_ao4 i_143138682(.A(n_22976), .B(n_32352), .C(n_28089), .D(n_33372
		), .Z(n_345874800));
	notech_ao4 i_143038683(.A(n_22980), .B(n_32764), .C(n_22977), .D(n_32782
		), .Z(n_345974801));
	notech_ao4 i_142838685(.A(n_22985), .B(n_33371), .C(n_22984), .D(n_32747
		), .Z(n_346174803));
	notech_and4 i_143338680(.A(n_57878), .B(n_346174803), .C(n_345974801), .D
		(n_345874800), .Z(n_346374805));
	notech_ao4 i_142438689(.A(n_335174693), .B(\nbus_11283[27] ), .C(n_219973567
		), .D(nbus_11273[11]), .Z(n_346574807));
	notech_ao4 i_142338690(.A(n_57928), .B(n_31484), .C(n_335374695), .D(n_32848
		), .Z(n_346674808));
	notech_ao4 i_142138692(.A(n_301374365), .B(\nbus_11290[3] ), .C(n_301274364
		), .D(n_31476), .Z(n_346874810));
	notech_ao4 i_142038693(.A(n_57917), .B(nbus_11273[3]), .C(n_57998), .D(n_32039
		), .Z(n_346974811));
	notech_and4 i_142638687(.A(n_346974811), .B(n_346874810), .C(n_346674808
		), .D(n_346574807), .Z(n_347174813));
	notech_ao4 i_141738696(.A(n_57867), .B(n_33258), .C(n_58512), .D(\nbus_11290[11] 
		), .Z(n_347274814));
	notech_ao4 i_141638697(.A(n_23329), .B(n_32462), .C(n_57887), .D(n_32507
		), .Z(n_347374815));
	notech_ao4 i_141438699(.A(n_58007), .B(nbus_11271[11]), .C(n_57987), .D(n_33370
		), .Z(n_347574817));
	notech_and4 i_141938694(.A(n_347574817), .B(n_347374815), .C(n_347274814
		), .D(n_252973897), .Z(n_347774819));
	notech_ao4 i_141038703(.A(n_30611), .B(n_31059), .C(n_58492), .D(n_31182
		), .Z(n_347974821));
	notech_ao4 i_140938704(.A(n_23359), .B(n_31230), .C(n_57745), .D(n_32392
		), .Z(n_348074822));
	notech_ao4 i_140738706(.A(n_22979), .B(\nbus_11290[27] ), .C(n_23383), .D
		(n_31210), .Z(n_348274824));
	notech_ao4 i_140638707(.A(n_22968), .B(n_32832), .C(n_22967), .D(n_32815
		), .Z(n_348374825));
	notech_and4 i_141238701(.A(n_348374825), .B(n_348274824), .C(n_348074822
		), .D(n_347974821), .Z(n_348574827));
	notech_ao4 i_140338710(.A(n_22976), .B(n_32351), .C(n_28089), .D(n_33369
		), .Z(n_348674828));
	notech_ao4 i_140238711(.A(n_22980), .B(n_32763), .C(n_22977), .D(n_32781
		), .Z(n_348774829));
	notech_ao4 i_140038713(.A(n_22985), .B(n_33368), .C(n_22984), .D(n_32746
		), .Z(n_348974831));
	notech_and4 i_140538708(.A(n_57878), .B(n_348974831), .C(n_348774829), .D
		(n_348674828), .Z(n_349174833));
	notech_ao4 i_139638717(.A(n_335174693), .B(\nbus_11283[26] ), .C(n_219773565
		), .D(nbus_11273[10]), .Z(n_349374835));
	notech_ao4 i_139538718(.A(n_57928), .B(n_31483), .C(n_335374695), .D(n_32847
		), .Z(n_349474836));
	notech_ao4 i_139238720(.A(n_301374365), .B(\nbus_11290[2] ), .C(n_301274364
		), .D(n_31474), .Z(n_349674838));
	notech_ao4 i_139138721(.A(n_57917), .B(nbus_11273[2]), .C(n_57998), .D(n_32038
		), .Z(n_349774839));
	notech_and4 i_139838715(.A(n_349774839), .B(n_349674838), .C(n_349474836
		), .D(n_349374835), .Z(n_349974841));
	notech_ao4 i_138738724(.A(n_23329), .B(n_32461), .C(n_57887), .D(n_32504
		), .Z(n_350074842));
	notech_ao4 i_138638725(.A(n_58007), .B(nbus_11271[10]), .C(n_57987), .D(n_33367
		), .Z(n_350174843));
	notech_ao4 i_138438727(.A(n_58492), .B(n_31181), .C(n_58215), .D(n_32431
		), .Z(n_350474845));
	notech_and4 i_138938722(.A(n_350474845), .B(n_350174843), .C(n_350074842
		), .D(n_250073868), .Z(n_350974847));
	notech_ao4 i_138038731(.A(n_57745), .B(n_32389), .C(n_30611), .D(n_31058
		), .Z(n_351174849));
	notech_ao4 i_137938732(.A(n_23359), .B(n_31229), .C(n_57867), .D(n_33204
		), .Z(n_351274850));
	notech_ao4 i_137738734(.A(n_22979), .B(\nbus_11290[26] ), .C(n_23383), .D
		(n_31209), .Z(n_351474852));
	notech_ao4 i_137638735(.A(n_22968), .B(n_32831), .C(n_22967), .D(n_32814
		), .Z(n_351574853));
	notech_and4 i_138238729(.A(n_351574853), .B(n_351474852), .C(n_351274850
		), .D(n_351174849), .Z(n_351774855));
	notech_ao4 i_137338738(.A(n_22976), .B(n_32350), .C(n_28089), .D(n_33366
		), .Z(n_351874856));
	notech_ao4 i_137238739(.A(n_22980), .B(n_32762), .C(n_22977), .D(n_32780
		), .Z(n_351974857));
	notech_ao4 i_137038741(.A(n_22985), .B(n_33365), .C(n_22984), .D(n_32745
		), .Z(n_352174859));
	notech_and4 i_137538736(.A(n_57878), .B(n_352174859), .C(n_351974857), .D
		(n_351874856), .Z(n_352374861));
	notech_ao4 i_136638745(.A(n_335174693), .B(\nbus_11283[25] ), .C(n_219573563
		), .D(nbus_11273[9]), .Z(n_352574863));
	notech_ao4 i_136538746(.A(n_57928), .B(n_31482), .C(n_335374695), .D(n_32846
		), .Z(n_352674864));
	notech_ao4 i_136338748(.A(n_301374365), .B(n_59005), .C(n_301274364), .D
		(n_31473), .Z(n_352874866));
	notech_ao4 i_136238749(.A(n_57917), .B(nbus_11273[1]), .C(n_57998), .D(n_32037
		), .Z(n_352974867));
	notech_and4 i_136838743(.A(n_352974867), .B(n_352874866), .C(n_352674864
		), .D(n_352574863), .Z(n_353174869));
	notech_ao4 i_135938752(.A(n_23329), .B(n_32460), .C(n_57887), .D(n_32503
		), .Z(n_353274870));
	notech_ao4 i_135838753(.A(n_58007), .B(nbus_11271[9]), .C(n_57987), .D(n_33364
		), .Z(n_353374871));
	notech_ao4 i_135638755(.A(n_58492), .B(n_31180), .C(n_58215), .D(n_32430
		), .Z(n_353574873));
	notech_and4 i_136138750(.A(n_353574873), .B(n_353374871), .C(n_353274870
		), .D(n_247173839), .Z(n_353774875));
	notech_ao4 i_135238759(.A(n_57745), .B(n_32387), .C(n_30611), .D(n_31057
		), .Z(n_353974877));
	notech_ao4 i_135138760(.A(n_23359), .B(n_31228), .C(n_57867), .D(n_33168
		), .Z(n_354074878));
	notech_ao4 i_134938762(.A(n_22979), .B(\nbus_11290[25] ), .C(n_23383), .D
		(n_31208), .Z(n_354274880));
	notech_ao4 i_134838763(.A(n_22968), .B(n_32830), .C(n_22967), .D(n_32813
		), .Z(n_354374881));
	notech_and4 i_135438757(.A(n_354374881), .B(n_354274880), .C(n_354074878
		), .D(n_353974877), .Z(n_354574883));
	notech_ao4 i_134538766(.A(n_22976), .B(n_32349), .C(n_28089), .D(n_33363
		), .Z(n_354674884));
	notech_ao4 i_134438767(.A(n_22980), .B(n_32761), .C(n_22977), .D(n_32778
		), .Z(n_354774885));
	notech_ao4 i_134238769(.A(n_22985), .B(n_33362), .C(n_22984), .D(n_32744
		), .Z(n_354974887));
	notech_and4 i_134738764(.A(n_57878), .B(n_354974887), .C(n_354774885), .D
		(n_354674884), .Z(n_355174889));
	notech_ao4 i_133838773(.A(n_335174693), .B(\nbus_11283[24] ), .C(n_219373561
		), .D(nbus_11273[8]), .Z(n_355374891));
	notech_ao4 i_133738774(.A(n_57928), .B(n_31481), .C(n_335374695), .D(n_32845
		), .Z(n_355474892));
	notech_ao4 i_133538776(.A(n_301374365), .B(\nbus_11290[0] ), .C(n_301274364
		), .D(n_31472), .Z(n_355674894));
	notech_ao4 i_133438777(.A(n_57917), .B(nbus_11273[0]), .C(n_57998), .D(n_32036
		), .Z(n_355774895));
	notech_and4 i_134038771(.A(n_355774895), .B(n_355674894), .C(n_355474892
		), .D(n_355374891), .Z(n_355974897));
	notech_ao4 i_133138780(.A(n_23329), .B(n_32459), .C(n_57887), .D(n_32502
		), .Z(n_356074898));
	notech_ao4 i_133038781(.A(n_58007), .B(nbus_11271[8]), .C(n_57987), .D(n_33361
		), .Z(n_356174899));
	notech_ao4 i_132838783(.A(n_58492), .B(n_31179), .C(n_58215), .D(n_32429
		), .Z(n_356374901));
	notech_and4 i_133338778(.A(n_356374901), .B(n_356174899), .C(n_356074898
		), .D(n_244273810), .Z(n_356574903));
	notech_ao4 i_132438787(.A(n_57745), .B(n_32385), .C(n_30611), .D(n_31056
		), .Z(n_356774905));
	notech_ao4 i_132338788(.A(n_23359), .B(n_31227), .C(n_57867), .D(n_33253
		), .Z(n_356874906));
	notech_ao4 i_132138790(.A(n_22979), .B(\nbus_11290[24] ), .C(n_23383), .D
		(n_31207), .Z(n_357074908));
	notech_ao4 i_132038791(.A(n_22968), .B(n_32829), .C(n_22967), .D(n_32812
		), .Z(n_357174909));
	notech_and4 i_132638785(.A(n_357174909), .B(n_357074908), .C(n_356874906
		), .D(n_356774905), .Z(n_357374911));
	notech_ao4 i_131738794(.A(n_22976), .B(n_32348), .C(n_28089), .D(n_33360
		), .Z(n_357474912));
	notech_ao4 i_131638795(.A(n_22980), .B(n_32760), .C(n_22977), .D(n_32777
		), .Z(n_357574913));
	notech_ao4 i_131438797(.A(n_22985), .B(n_33359), .C(n_22984), .D(n_32743
		), .Z(n_357774915));
	notech_and4 i_131938792(.A(n_57878), .B(n_357774915), .C(n_357574913), .D
		(n_357474912), .Z(n_357974917));
	notech_ao4 i_130038810(.A(n_57917), .B(nbus_11273[15]), .C(n_57998), .D(n_32035
		), .Z(n_358174919));
	notech_ao4 i_129838812(.A(n_57887), .B(n_32501), .C(n_58007), .D(nbus_11271
		[7]), .Z(n_358374921));
	notech_and4 i_130238808(.A(n_358374921), .B(n_358174919), .C(n_241173779
		), .D(n_241473782), .Z(n_358574923));
	notech_ao4 i_129538815(.A(n_58215), .B(n_32428), .C(n_57987), .D(n_33357
		), .Z(n_358674924));
	notech_ao4 i_129338817(.A(n_57745), .B(n_32384), .C(n_31055), .D(n_30611
		), .Z(n_358874926));
	notech_and4 i_129738813(.A(n_358874926), .B(n_358674924), .C(n_240573773
		), .D(n_240873776), .Z(n_359074928));
	notech_ao4 i_128738821(.A(n_23383), .B(n_31206), .C(n_23359), .D(n_31226
		), .Z(n_359274930));
	notech_ao4 i_128538823(.A(n_22968), .B(n_32828), .C(n_22967), .D(n_32811
		), .Z(n_359474932));
	notech_and4 i_128938819(.A(n_359474932), .B(n_240273770), .C(n_359274930
		), .D(n_239973767), .Z(n_359674934));
	notech_ao4 i_128238826(.A(n_22977), .B(n_32776), .C(n_22976), .D(n_32347
		), .Z(n_359774935));
	notech_or4 i_131338798(.A(n_27922), .B(n_30687), .C(n_61625), .D(opa[7])
		, .Z(n_359974937));
	notech_ao4 i_131238799(.A(n_22752), .B(n_30270), .C(n_61625), .D(n_219273560
		), .Z(n_360074938));
	notech_ao4 i_130938802(.A(n_219173559), .B(nbus_11273[7]), .C(n_359974937
		), .D(n_27829), .Z(n_360274940));
	notech_ao4 i_130838803(.A(n_22984), .B(n_32742), .C(n_57907), .D(\nbus_11290[15] 
		), .Z(n_360374941));
	notech_ao4 i_130538805(.A(n_22742), .B(n_31480), .C(n_22985), .D(n_33358
		), .Z(n_360574943));
	notech_ao4 i_130438806(.A(n_30610), .B(n_32701), .C(n_22745), .D(n_32844
		), .Z(n_360674944));
	notech_and4 i_18160(.A(n_360674944), .B(n_360574943), .C(n_360374941), .D
		(n_360274940), .Z(n_360874946));
	notech_and4 i_128438824(.A(n_57878), .B(n_360874946), .C(n_359774935), .D
		(n_239673764), .Z(n_361074948));
	notech_or4 i_128038828(.A(n_27922), .B(n_30687), .C(n_61625), .D(opa[6])
		, .Z(n_361274950));
	notech_ao4 i_127938829(.A(nbus_11291[6]), .B(n_57896), .C(n_22752), .D(n_30271
		), .Z(n_361374951));
	notech_ao4 i_127538833(.A(nbus_11273[6]), .B(n_219073558), .C(n_105014667
		), .D(n_361274950), .Z(n_361474952));
	notech_ao4 i_127438834(.A(n_57917), .B(nbus_11273[14]), .C(n_57998), .D(n_32034
		), .Z(n_361574953));
	notech_ao4 i_127238836(.A(n_58007), .B(nbus_11271[6]), .C(n_57907), .D(\nbus_11290[14] 
		), .Z(n_361774955));
	notech_ao4 i_127138837(.A(n_57887), .B(n_32500), .C(n_58512), .D(\nbus_11290[6] 
		), .Z(n_361874956));
	notech_and4 i_127738831(.A(n_361874956), .B(n_361774955), .C(n_361574953
		), .D(n_361474952), .Z(n_362074958));
	notech_ao4 i_126838840(.A(n_57987), .B(n_33356), .C(n_23329), .D(n_32457
		), .Z(n_362174959));
	notech_ao4 i_126738841(.A(n_58492), .B(n_31178), .C(n_58215), .D(n_32427
		), .Z(n_362274960));
	notech_ao4 i_126538843(.A(n_57745), .B(n_32382), .C(n_30611), .D(n_31054
		), .Z(n_362474962));
	notech_and4 i_127038838(.A(n_362474962), .B(n_362274960), .C(n_362174959
		), .D(n_237973747), .Z(n_362674964));
	notech_ao4 i_126138847(.A(n_23383), .B(n_31205), .C(n_23359), .D(n_31225
		), .Z(n_362874966));
	notech_ao4 i_126038848(.A(n_22967), .B(n_32810), .C(n_22979), .D(\nbus_11290[22] 
		), .Z(n_362974967));
	notech_ao4 i_125838850(.A(n_28089), .B(n_32591), .C(n_22968), .D(n_32827
		), .Z(n_363174969));
	notech_and4 i_126338845(.A(n_363174969), .B(n_362974967), .C(n_362874966
		), .D(n_237273740), .Z(n_363374971));
	notech_ao4 i_125538853(.A(n_22980), .B(n_32759), .C(n_22977), .D(n_32775
		), .Z(n_363474972));
	notech_ao4 i_125438854(.A(n_22985), .B(n_33355), .C(n_22984), .D(n_32741
		), .Z(n_363574973));
	notech_ao4 i_125238856(.A(n_22745), .B(n_32843), .C(n_22742), .D(n_31479
		), .Z(n_363774975));
	notech_and4 i_125738851(.A(n_363774975), .B(n_363574973), .C(n_363474972
		), .D(n_236573733), .Z(n_363974976));
	notech_nao3 i_125138857(.A(n_27826), .B(n_27832), .C(n_30687), .Z(n_364174978
		));
	notech_ao4 i_125038858(.A(n_22752), .B(n_27832), .C(n_57896), .D(nbus_11291
		[4]), .Z(n_364274979));
	notech_mux2 i_124638862(.S(opa[4]), .A(n_364174978), .B(n_218973557), .Z
		(n_364374980));
	notech_ao4 i_124538863(.A(n_23379), .B(n_32032), .C(n_58007), .D(nbus_11271
		[4]), .Z(n_364474981));
	notech_ao4 i_124338865(.A(n_57907), .B(\nbus_11290[12] ), .C(n_57917), .D
		(nbus_11273[12]), .Z(n_364674983));
	notech_ao4 i_124238866(.A(n_57887), .B(n_32494), .C(n_58512), .D(\nbus_11290[4] 
		), .Z(n_364774984));
	notech_and4 i_124838860(.A(n_364774984), .B(n_364674983), .C(n_364474981
		), .D(n_364374980), .Z(n_365074986));
	notech_ao4 i_123938869(.A(n_57987), .B(n_33354), .C(n_23329), .D(n_32456
		), .Z(n_365174987));
	notech_ao4 i_123838870(.A(n_58492), .B(n_31176), .C(n_58215), .D(n_32426
		), .Z(n_365274988));
	notech_ao4 i_123638872(.A(n_57745), .B(n_32381), .C(n_30611), .D(n_31053
		), .Z(n_365474990));
	notech_and4 i_124138867(.A(n_365474990), .B(n_365274988), .C(n_365174987
		), .D(n_234873716), .Z(n_365674992));
	notech_ao4 i_123238876(.A(n_23383), .B(n_31204), .C(n_23359), .D(n_31223
		), .Z(n_365874994));
	notech_ao4 i_123138877(.A(n_22967), .B(n_32808), .C(n_22979), .D(n_58857
		), .Z(n_365974995));
	notech_ao4 i_122938879(.A(n_28089), .B(n_32588), .C(n_22968), .D(n_32825
		), .Z(n_366174997));
	notech_and4 i_123438874(.A(n_366174997), .B(n_365974995), .C(n_365874994
		), .D(n_234173709), .Z(n_366374999));
	notech_ao4 i_122638882(.A(n_22980), .B(n_32758), .C(n_22977), .D(n_32773
		), .Z(n_366475000));
	notech_ao4 i_122538883(.A(n_22985), .B(n_33353), .C(n_22984), .D(n_32740
		), .Z(n_366575001));
	notech_ao4 i_122338885(.A(n_22745), .B(n_32842), .C(n_22742), .D(n_31477
		), .Z(n_366775003));
	notech_and4 i_122838880(.A(n_366775003), .B(n_366575001), .C(n_366475000
		), .D(n_233473702), .Z(n_366975005));
	notech_nand2 i_122238886(.A(n_27833), .B(nbus_11273[3]), .Z(n_367175007)
		);
	notech_ao4 i_122138887(.A(n_22752), .B(n_27833), .C(n_57896), .D(nbus_11291
		[3]), .Z(n_367275008));
	notech_ao4 i_121738891(.A(nbus_11273[3]), .B(n_218873556), .C(n_22752), 
		.D(n_367175007), .Z(n_367375009));
	notech_ao4 i_121638892(.A(n_57998), .B(n_32031), .C(n_58007), .D(nbus_11271
		[3]), .Z(n_367475010));
	notech_ao4 i_121438894(.A(n_57907), .B(\nbus_11290[11] ), .C(n_57917), .D
		(nbus_11273[11]), .Z(n_367675012));
	notech_ao4 i_121338895(.A(n_23329), .B(n_32455), .C(n_57887), .D(n_32493
		), .Z(n_367775013));
	notech_and4 i_121938889(.A(n_367775013), .B(n_367675012), .C(n_367475010
		), .D(n_367375009), .Z(n_367975015));
	notech_ao4 i_121038898(.A(n_58215), .B(n_32425), .C(n_57987), .D(n_33352
		), .Z(n_368075016));
	notech_ao4 i_120938899(.A(n_58512), .B(\nbus_11290[3] ), .C(n_23353), .D
		(n_31175), .Z(n_368175017));
	notech_ao4 i_120738901(.A(n_57745), .B(n_32380), .C(n_30611), .D(n_31052
		), .Z(n_368375019));
	notech_and4 i_121238896(.A(n_368375019), .B(n_368175017), .C(n_368075016
		), .D(n_231773685), .Z(n_368575021));
	notech_ao4 i_120338905(.A(n_23383), .B(n_31203), .C(n_23359), .D(n_31222
		), .Z(n_368875023));
	notech_ao4 i_120238906(.A(n_22967), .B(n_32807), .C(n_22979), .D(\nbus_11290[19] 
		), .Z(n_368975024));
	notech_ao4 i_120038908(.A(n_28089), .B(n_32587), .C(n_22968), .D(n_32824
		), .Z(n_369175026));
	notech_and4 i_120538903(.A(n_369175026), .B(n_368975024), .C(n_368875023
		), .D(n_231073678), .Z(n_369375028));
	notech_ao4 i_119738911(.A(n_22980), .B(n_32757), .C(n_22977), .D(n_32772
		), .Z(n_369475029));
	notech_ao4 i_119638912(.A(n_22985), .B(n_33351), .C(n_22984), .D(n_32739
		), .Z(n_369575030));
	notech_ao4 i_119438914(.A(n_22745), .B(n_32841), .C(n_22742), .D(n_31476
		), .Z(n_369775032));
	notech_and4 i_119938909(.A(n_369775032), .B(n_369575030), .C(n_369475029
		), .D(n_230373671), .Z(n_369975034));
	notech_ao4 i_116038947(.A(n_22752), .B(n_316151269), .C(n_218673554), .D
		(nbus_11273[1]), .Z(n_370175036));
	notech_ao4 i_115938948(.A(n_57917), .B(nbus_11273[9]), .C(n_57998), .D(n_32029
		), .Z(n_370275037));
	notech_ao4 i_115738950(.A(n_57887), .B(n_32491), .C(n_57907), .D(\nbus_11290[9] 
		), .Z(n_370475039));
	notech_ao4 i_115638951(.A(n_57987), .B(n_33350), .C(n_23329), .D(n_32453
		), .Z(n_370575040));
	notech_and4 i_116238945(.A(n_370575040), .B(n_370475039), .C(n_370275037
		), .D(n_370175036), .Z(n_3707));
	notech_ao4 i_115338954(.A(n_58215), .B(n_32423), .C(n_58007), .D(nbus_11271
		[1]), .Z(n_3708));
	notech_ao4 i_115238955(.A(n_58512), .B(\nbus_11290[1] ), .C(n_58492), .D
		(n_31173), .Z(n_3709));
	notech_ao4 i_115038957(.A(n_57745), .B(n_32377), .C(n_30611), .D(n_31051
		), .Z(n_3711));
	notech_and4 i_115538952(.A(n_3711), .B(n_3709), .C(n_3708), .D(n_228873656
		), .Z(n_3713));
	notech_ao4 i_114638961(.A(n_23383), .B(n_31201), .C(n_23359), .D(n_31219
		), .Z(n_371575042));
	notech_ao4 i_114538962(.A(n_22967), .B(n_32805), .C(n_22979), .D(\nbus_11290[17] 
		), .Z(n_371675043));
	notech_ao4 i_114338964(.A(n_28089), .B(n_32585), .C(n_22968), .D(n_32822
		), .Z(n_371875045));
	notech_and4 i_114838959(.A(n_371875045), .B(n_371675043), .C(n_371575042
		), .D(n_228173649), .Z(n_372075047));
	notech_ao4 i_114038967(.A(n_22980), .B(n_32754), .C(n_22977), .D(n_32770
		), .Z(n_372175048));
	notech_ao4 i_113938968(.A(n_22985), .B(n_33349), .C(n_22984), .D(n_32737
		), .Z(n_372275049));
	notech_ao4 i_113738970(.A(n_22745), .B(n_32839), .C(n_22742), .D(n_31473
		), .Z(n_372475051));
	notech_and4 i_114238965(.A(n_372475051), .B(n_372275049), .C(n_372175048
		), .D(n_227473642), .Z(n_3726));
	notech_ao4 i_113238975(.A(n_57998), .B(n_32028), .C(nbus_11273[0]), .D(n_218573553
		), .Z(n_3729));
	notech_ao4 i_113138976(.A(n_57907), .B(\nbus_11290[8] ), .C(n_57917), .D
		(nbus_11273[8]), .Z(n_3730));
	notech_ao4 i_112938978(.A(n_23329), .B(n_32452), .C(n_57887), .D(n_32490
		), .Z(n_3732));
	notech_and4 i_113438973(.A(n_3732), .B(n_3730), .C(n_3729), .D(n_226673634
		), .Z(n_3734));
	notech_ao4 i_112638981(.A(n_58215), .B(n_32422), .C(n_58007), .D(nbus_11271
		[0]), .Z(n_3735));
	notech_ao4 i_112538982(.A(n_58512), .B(\nbus_11290[0] ), .C(n_58492), .D
		(n_31172), .Z(n_3736));
	notech_ao4 i_112338984(.A(n_57745), .B(n_32376), .C(n_30611), .D(n_32451
		), .Z(n_3738));
	notech_and4 i_112838979(.A(n_3738), .B(n_3736), .C(n_3735), .D(n_225973627
		), .Z(n_3740));
	notech_ao4 i_111938988(.A(n_23383), .B(n_31200), .C(n_23359), .D(n_31217
		), .Z(n_374275054));
	notech_ao4 i_111838989(.A(n_22967), .B(n_32804), .C(n_22979), .D(\nbus_11290[16] 
		), .Z(n_374375055));
	notech_ao4 i_111638991(.A(n_28089), .B(n_32584), .C(n_22968), .D(n_32821
		), .Z(n_374575057));
	notech_and4 i_112138986(.A(n_374575057), .B(n_374375055), .C(n_374275054
		), .D(n_225273620), .Z(n_3747));
	notech_ao4 i_111338994(.A(n_22980), .B(n_32753), .C(n_22977), .D(n_32769
		), .Z(n_374875059));
	notech_ao4 i_111238995(.A(n_22985), .B(n_33348), .C(n_22984), .D(n_32736
		), .Z(n_374975060));
	notech_ao4 i_111038997(.A(n_22745), .B(n_32838), .C(n_22742), .D(n_31472
		), .Z(n_375175062));
	notech_and4 i_111538992(.A(n_375175062), .B(n_374975060), .C(n_374875059
		), .D(n_224573613), .Z(n_375375064));
	notech_and4 i_621764(.A(n_144272827), .B(n_144172826), .C(n_143672821), 
		.D(n_144072825), .Z(n_15200));
	notech_and4 i_521763(.A(n_145972844), .B(n_145872843), .C(n_145372838), 
		.D(n_145772842), .Z(n_15194));
	notech_nand2 i_3353041(.A(n_61625), .B(read_data[20]), .Z(n_375575066)
		);
	notech_nao3 i_29854(.A(n_29557), .B(n_63764), .C(n_386664397), .Z(n_303922064
		));
	notech_or2 i_29871(.A(n_444168025), .B(n_57062), .Z(n_303822063));
	notech_nao3 i_136146413(.A(n_290663806), .B(instrc[117]), .C(n_217173539
		), .Z(n_299122016));
	notech_and4 i_118746467(.A(n_29550), .B(n_30697), .C(n_57612), .D(n_217673544
		), .Z(n_57319));
	notech_and4 i_118646466(.A(n_29540), .B(n_30689), .C(n_57611), .D(n_217573543
		), .Z(n_57320));
	notech_and3 i_114346465(.A(n_29533), .B(n_217473542), .C(n_30693), .Z(n_57362
		));
	notech_ao4 i_114246464(.A(n_335360981), .B(n_61625), .C(n_386664397), .D
		(n_386964400), .Z(n_57363));
	notech_ao4 i_175244761(.A(n_30860), .B(n_61103), .C(n_321271180), .D(n_336760995
		), .Z(n_271670708));
	notech_or4 i_87555981(.A(n_318060808), .B(n_2577), .C(n_286263764), .D(n_29560
		), .Z(n_57611));
	notech_or2 i_87455982(.A(n_386964400), .B(n_29560), .Z(n_57612));
	notech_and4 i_175944754(.A(n_271270705), .B(n_271070703), .C(n_253370528
		), .D(n_253670531), .Z(n_271570707));
	notech_nand3 i_3217758(.A(n_303474386), .B(n_302974381), .C(n_303874390)
		, .Z(n_17234));
	notech_nand3 i_3117757(.A(n_305474406), .B(n_304974401), .C(n_305874410)
		, .Z(n_17228));
	notech_nand3 i_3017756(.A(n_307474426), .B(n_306974421), .C(n_307874430)
		, .Z(n_17222));
	notech_nand3 i_2917755(.A(n_309874450), .B(n_309474446), .C(n_308974441)
		, .Z(n_17216));
	notech_nand3 i_2817754(.A(n_311474466), .B(n_310974461), .C(n_311874470)
		, .Z(n_17210));
	notech_nand3 i_2717753(.A(n_313474486), .B(n_312974481), .C(n_313874490)
		, .Z(n_17204));
	notech_nand3 i_2617752(.A(n_315574506), .B(n_314974501), .C(n_316074510)
		, .Z(n_17198));
	notech_nand3 i_2517751(.A(n_317674526), .B(n_317174521), .C(n_318074530)
		, .Z(n_17192));
	notech_nand3 i_2417750(.A(n_319774546), .B(n_319174541), .C(n_320274550)
		, .Z(n_17186));
	notech_nand3 i_2317749(.A(n_321874566), .B(n_321374561), .C(n_322274570)
		, .Z(n_17180));
	notech_nand3 i_2217748(.A(n_322974576), .B(n_324574591), .C(n_323474580)
		, .Z(n_17174));
	notech_nand3 i_2117747(.A(n_326474610), .B(n_326074606), .C(n_325574601)
		, .Z(n_17168));
	notech_nand3 i_2017746(.A(n_328674630), .B(n_328274626), .C(n_327774621)
		, .Z(n_17162));
	notech_nand3 i_1917745(.A(n_330674650), .B(n_330274646), .C(n_329774641)
		, .Z(n_17156));
	notech_nand3 i_1817744(.A(n_332874670), .B(n_332474666), .C(n_331774661)
		, .Z(n_17150));
	notech_nand3 i_1717743(.A(n_333474676), .B(n_334974691), .C(n_333874680)
		, .Z(n_17144));
	notech_and4 i_1617742(.A(n_337974721), .B(n_337374715), .C(n_336574707),
		 .D(n_335974701), .Z(n_17138));
	notech_and4 i_1517741(.A(n_340774749), .B(n_340174743), .C(n_339374735),
		 .D(n_338774729), .Z(n_17132));
	notech_and4 i_1417740(.A(n_343574777), .B(n_342974771), .C(n_342174763),
		 .D(n_341574757), .Z(n_17126));
	notech_and4 i_1317739(.A(n_346374805), .B(n_345774799), .C(n_344974791),
		 .D(n_344374785), .Z(n_17120));
	notech_and4 i_1217738(.A(n_349174833), .B(n_348574827), .C(n_347774819),
		 .D(n_347174813), .Z(n_17114));
	notech_and4 i_1117737(.A(n_352374861), .B(n_351774855), .C(n_350974847),
		 .D(n_349974841), .Z(n_17108));
	notech_and4 i_1017736(.A(n_355174889), .B(n_354574883), .C(n_353774875),
		 .D(n_353174869), .Z(n_17102));
	notech_and4 i_917735(.A(n_357974917), .B(n_357374911), .C(n_356574903), 
		.D(n_355974897), .Z(n_17096));
	notech_and4 i_817734(.A(n_361074948), .B(n_359674934), .C(n_359074928), 
		.D(n_358574923), .Z(n_17090));
	notech_and4 i_717733(.A(n_363974976), .B(n_363374971), .C(n_362674964), 
		.D(n_362074958), .Z(n_17084));
	notech_and4 i_517731(.A(n_366975005), .B(n_366374999), .C(n_365674992), 
		.D(n_365074986), .Z(n_17072));
	notech_and4 i_417730(.A(n_369975034), .B(n_369375028), .C(n_368575021), 
		.D(n_367975015), .Z(n_17066));
	notech_and4 i_217728(.A(n_3726), .B(n_372075047), .C(n_3713), .D(n_3707)
		, .Z(n_17054));
	notech_and4 i_117727(.A(n_375375064), .B(n_3747), .C(n_3740), .D(n_3734)
		, .Z(n_17048));
	notech_or4 i_71240086(.A(n_61889), .B(n_1834), .C(n_61725), .D(nbus_11273
		[7]), .Z(n_317751253));
	notech_xor2 i_165440070(.A(nbus_11273[1]), .B(opa[0]), .Z(n_316151269)
		);
	notech_ao4 i_175544758(.A(n_58042), .B(n_31472), .C(n_327660904), .D(n_249870493
		), .Z(n_271270705));
	notech_ao4 i_175744756(.A(\nbus_11290[0] ), .B(n_250170496), .C(nbus_11273
		[0]), .D(n_250070495), .Z(n_271070703));
	notech_and4 i_176544748(.A(n_270770700), .B(n_270570698), .C(n_270470697
		), .D(n_253970534), .Z(n_270970702));
	notech_ao4 i_176044753(.A(n_318871159), .B(n_33311), .C(n_309771080), .D
		(n_33103), .Z(n_270770700));
	notech_ao4 i_176244751(.A(n_334360971), .B(n_309671079), .C(n_61099), .D
		(n_30861), .Z(n_270570698));
	notech_ao4 i_176344750(.A(n_334060968), .B(n_321271180), .C(n_31473), .D
		(n_58042), .Z(n_270470697));
	notech_and4 i_177144742(.A(n_270170694), .B(n_269970692), .C(n_269870691
		), .D(n_254670541), .Z(n_270370696));
	notech_ao4 i_176644747(.A(n_30896), .B(n_262170616), .C(n_30891), .D(n_57441
		), .Z(n_270170694));
	notech_ao4 i_176844745(.A(n_30914), .B(n_249870493), .C(n_30916), .D(n_249970494
		), .Z(n_269970692));
	notech_ao4 i_176944744(.A(n_250370498), .B(n_262270617), .C(n_310271084)
		, .D(n_250270497), .Z(n_269870691));
	notech_and4 i_177744736(.A(n_269570688), .B(n_269370686), .C(n_269270685
		), .D(n_255370548), .Z(n_269770690));
	notech_ao4 i_177244741(.A(n_318871159), .B(n_33312), .C(n_310371085), .D
		(n_33253), .Z(n_269570688));
	notech_ao4 i_177444739(.A(n_5269), .B(n_310771089), .C(n_61099), .D(n_30873
		), .Z(n_269370686));
	notech_ao4 i_177544738(.A(n_30326), .B(n_33313), .C(n_309871081), .D(n_300722032
		), .Z(n_269270685));
	notech_ao4 i_178444729(.A(n_57117), .B(n_31779), .C(n_57616), .D(n_33314
		), .Z(n_268970682));
	notech_ao4 i_178544728(.A(n_57141), .B(n_31747), .C(n_57157), .D(n_33315
		), .Z(n_268870681));
	notech_and2 i_178944724(.A(n_268670679), .B(n_268570678), .Z(n_268770680
		));
	notech_ao4 i_178744726(.A(n_57168), .B(n_31843), .C(n_30590), .D(n_32004
		), .Z(n_268670679));
	notech_ao4 i_178844725(.A(n_57192), .B(n_31715), .C(n_30679), .D(n_31939
		), .Z(n_268570678));
	notech_and4 i_179744716(.A(n_268270675), .B(n_268170674), .C(n_267970672
		), .D(n_267870671), .Z(n_268470677));
	notech_ao4 i_179144722(.A(n_57062), .B(n_31683), .C(n_57072), .D(n_31811
		), .Z(n_268270675));
	notech_ao4 i_179244721(.A(n_57086), .B(n_31875), .C(n_57103), .D(n_31580
		), .Z(n_268170674));
	notech_ao4 i_179444719(.A(n_58701), .B(n_31972), .C(n_59100), .D(n_31907
		), .Z(n_267970672));
	notech_ao4 i_179544718(.A(n_57218), .B(n_31416), .C(n_57230), .D(n_31651
		), .Z(n_267870671));
	notech_and4 i_178344730(.A(n_267570668), .B(n_267270665), .C(n_267070663
		), .D(n_256070555), .Z(n_267770670));
	notech_ao4 i_177844735(.A(n_267470667), .B(n_299422019), .C(n_265570648)
		, .D(nbus_11273[8]), .Z(n_267570668));
	notech_nao3 i_59146421(.A(n_61935), .B(opa[8]), .C(\opcode[1] ), .Z(n_267470667
		));
	notech_ao4 i_178044733(.A(n_299222017), .B(\nbus_11290[8] ), .C(n_267170664
		), .D(n_265370646), .Z(n_267270665));
	notech_nand2 i_10546427(.A(opc_10[8]), .B(n_63764), .Z(n_267170664));
	notech_ao4 i_178144732(.A(n_266970662), .B(n_265070645), .C(n_266870661)
		, .D(n_264970644), .Z(n_267070663));
	notech_nand2 i_60646419(.A(opc[8]), .B(n_63764), .Z(n_266970662));
	notech_nao3 i_60246420(.A(n_63792), .B(opa[8]), .C(\opcode[1] ), .Z(n_266870661
		));
	notech_and4 i_186244651(.A(n_266570658), .B(n_266370656), .C(n_258670581
		), .D(n_258370578), .Z(n_266770660));
	notech_ao4 i_185844655(.A(n_318871159), .B(n_33316), .C(n_310371085), .D
		(n_33215), .Z(n_266570658));
	notech_ao4 i_186044653(.A(n_61103), .B(n_30879), .C(n_309871081), .D(n_385364384
		), .Z(n_266370656));
	notech_and4 i_186744646(.A(n_266070653), .B(n_265870651), .C(n_258970584
		), .D(n_259270587), .Z(n_266270655));
	notech_ao4 i_186344650(.A(n_31487), .B(n_30325), .C(n_377264303), .D(n_265370646
		), .Z(n_266070653));
	notech_ao4 i_186544648(.A(\nbus_11290[14] ), .B(n_251370508), .C(nbus_11273
		[14]), .D(n_251270507), .Z(n_265870651));
	notech_or2 i_126546415(.A(n_299422019), .B(n_321871184), .Z(n_265570648)
		);
	notech_nao3 i_156146410(.A(n_56820), .B(n_3382), .C(n_310271084), .Z(n_265370646
		));
	notech_nao3 i_157846409(.A(n_56820), .B(n_3382), .C(n_299422019), .Z(n_265070645
		));
	notech_or2 i_164046406(.A(n_58274), .B(n_299422019), .Z(n_264970644));
	notech_and4 i_188744626(.A(n_264670641), .B(n_264470639), .C(n_259570590
		), .D(n_259870593), .Z(n_264870643));
	notech_ao4 i_188344630(.A(n_309971082), .B(\nbus_11283[31] ), .C(n_310671088
		), .D(\nbus_11290[31] ), .Z(n_264670641));
	notech_ao4 i_188544628(.A(n_311771098), .B(n_33206), .C(n_318971160), .D
		(n_31539), .Z(n_264470639));
	notech_and4 i_189244621(.A(n_264170636), .B(n_263970634), .C(n_260170596
		), .D(n_260470599), .Z(n_264370638));
	notech_ao4 i_188844625(.A(n_311471096), .B(n_31507), .C(n_61103), .D(n_30893
		), .Z(n_264170636));
	notech_ao4 i_189044623(.A(n_300822033), .B(n_311571097), .C(n_262470619)
		, .D(n_311271094), .Z(n_263970634));
	notech_ao4 i_189344620(.A(n_57117), .B(n_31802), .C(n_57609), .D(n_33317
		), .Z(n_263670631));
	notech_ao4 i_189444619(.A(n_57141), .B(n_31770), .C(n_57157), .D(n_33318
		), .Z(n_263570630));
	notech_and2 i_189844615(.A(n_263370628), .B(n_263270627), .Z(n_263470629
		));
	notech_ao4 i_189644617(.A(n_57168), .B(n_31866), .C(n_30590), .D(n_32027
		), .Z(n_263370628));
	notech_ao4 i_189744616(.A(n_57192), .B(n_31738), .C(n_30679), .D(n_31963
		), .Z(n_263270627));
	notech_and4 i_190644607(.A(n_262970624), .B(n_262870623), .C(n_262670621
		), .D(n_262570620), .Z(n_263170626));
	notech_ao4 i_190044613(.A(n_57062), .B(n_31706), .C(n_57072), .D(n_31834
		), .Z(n_262970624));
	notech_ao4 i_190144612(.A(n_57086), .B(n_31898), .C(n_58701), .D(n_31995
		), .Z(n_262870623));
	notech_ao4 i_190344610(.A(n_59100), .B(n_31930), .C(n_57218), .D(n_31439
		), .Z(n_262670621));
	notech_ao4 i_190444609(.A(n_57230), .B(n_31674), .C(n_57103), .D(n_31603
		), .Z(n_262570620));
	notech_nand2 i_2246428(.A(opc_10[31]), .B(n_63782), .Z(n_262470619));
	notech_and2 i_105046417(.A(n_310971091), .B(n_310571087), .Z(n_262270617
		));
	notech_or2 i_28166(.A(n_58274), .B(n_57441), .Z(n_262170616));
	notech_nand2 i_86045592(.A(\add_len_pc[31] ), .B(n_5680), .Z(n_260470599
		));
	notech_nand3 i_86345589(.A(n_2026), .B(n_6792), .C(n_32388), .Z(n_260170596
		));
	notech_or2 i_86645586(.A(n_5243), .B(n_311871099), .Z(n_259870593));
	notech_or2 i_87045583(.A(n_319071161), .B(nbus_11271[31]), .Z(n_259570590
		));
	notech_nao3 i_82045619(.A(n_63792), .B(opc[14]), .C(n_265070645), .Z(n_259270587
		));
	notech_nand2 i_82745616(.A(\add_len_pc[14] ), .B(n_5680), .Z(n_258970584
		));
	notech_or2 i_83045613(.A(n_97342414), .B(n_310771089), .Z(n_258670581)
		);
	notech_nao3 i_83345610(.A(n_19655), .B(read_data[14]), .C(n_60454), .Z(n_258370578
		));
	notech_nand2 i_72445715(.A(opd[8]), .B(n_300322028), .Z(n_256070555));
	notech_nao3 i_73145708(.A(n_19655), .B(read_data[8]), .C(n_60454), .Z(n_255370548
		));
	notech_nand2 i_70345735(.A(\add_len_pc[1] ), .B(n_5680), .Z(n_254670541)
		);
	notech_nao3 i_71045728(.A(n_19655), .B(read_data[1]), .C(n_60454), .Z(n_253970534
		));
	notech_nao3 i_68645751(.A(n_63792), .B(opc_10[0]), .C(n_249970494), .Z(n_253670531
		));
	notech_nand2 i_68945748(.A(\add_len_pc[0] ), .B(n_5680), .Z(n_253370528)
		);
	notech_or2 i_69245745(.A(n_101142452), .B(n_309671079), .Z(n_253070525)
		);
	notech_nao3 i_69545742(.A(n_19655), .B(read_data[0]), .C(n_60453), .Z(n_252770522
		));
	notech_or2 i_85645595(.A(n_262270617), .B(n_57501), .Z(n_251470509));
	notech_and3 i_1046397(.A(n_310671088), .B(n_309671079), .C(n_310871090),
		 .Z(n_251370508));
	notech_and3 i_946398(.A(n_309971082), .B(n_309771080), .C(n_310471086), 
		.Z(n_251270507));
	notech_ao4 i_1846393(.A(n_60175), .B(nbus_11273[1]), .C(n_30919), .D(n_58274
		), .Z(n_250770502));
	notech_ao4 i_1746394(.A(n_60175), .B(\nbus_11290[1] ), .C(n_30920), .D(n_58274
		), .Z(n_250570500));
	notech_ao4 i_1646395(.A(\nbus_11290[1] ), .B(n_57501), .C(nbus_11273[1])
		, .D(n_321871184), .Z(n_250370498));
	notech_mux2 i_1446396(.S(n_32304), .A(n_250770502), .B(n_250570500), .Z(n_250270497
		));
	notech_and3 i_2046391(.A(n_310871090), .B(n_310771089), .C(n_310671088),
		 .Z(n_250170496));
	notech_and3 i_1946392(.A(n_310471086), .B(n_309971082), .C(n_310371085),
		 .Z(n_250070495));
	notech_nao3 i_159346407(.A(n_56820), .B(n_3382), .C(n_310171083), .Z(n_249970494
		));
	notech_nao3 i_158346408(.A(n_56820), .B(n_3382), .C(n_57441), .Z(n_249870493
		));
	notech_and4 i_126548516(.A(n_246070456), .B(n_58055), .C(n_249470489), .D
		(n_249370488), .Z(n_249770492));
	notech_ao4 i_125948522(.A(n_24528), .B(n_33295), .C(n_24527), .D(n_33294
		), .Z(n_249470489));
	notech_and3 i_126448517(.A(n_249070485), .B(n_249270487), .C(n_214770148
		), .Z(n_249370488));
	notech_ao4 i_126148520(.A(n_381064341), .B(n_33118), .C(n_338361011), .D
		(n_380964340), .Z(n_249270487));
	notech_ao4 i_126248519(.A(n_31511), .B(n_60453), .C(n_61103), .D(n_30762
		), .Z(n_249070485));
	notech_ao4 i_126648515(.A(n_338161009), .B(n_24717), .C(n_74522848), .D(n_24421
		), .Z(n_248770482));
	notech_ao4 i_126748514(.A(n_74622849), .B(n_380764338), .C(n_74822851), 
		.D(n_24430), .Z(n_248670481));
	notech_and3 i_127248509(.A(n_215770157), .B(n_248270477), .C(n_248470479
		), .Z(n_248570480));
	notech_ao4 i_126948512(.A(n_75522858), .B(n_24428), .C(n_75622859), .D(n_24425
		), .Z(n_248470479));
	notech_ao4 i_127048511(.A(n_75222855), .B(n_24429), .C(n_74922852), .D(n_24424
		), .Z(n_248270477));
	notech_and4 i_127848503(.A(n_58055), .B(n_247970474), .C(n_247770472), .D
		(n_216270162), .Z(n_248170476));
	notech_ao4 i_127448507(.A(n_32186), .B(n_33296), .C(n_248736166), .D(nbus_11271
		[16]), .Z(n_247970474));
	notech_ao4 i_127648505(.A(n_57370), .B(\nbus_11290[16] ), .C(n_57325), .D
		(n_5444), .Z(n_247770472));
	notech_and4 i_128348498(.A(n_247470469), .B(n_247270467), .C(n_216570165
		), .D(n_216870168), .Z(n_247670471));
	notech_ao4 i_127948502(.A(n_60453), .B(n_31524), .C(n_385264383), .D(n_31489
		), .Z(n_247470469));
	notech_ao4 i_128148500(.A(n_58100), .B(n_320051171), .C(n_240370399), .D
		(n_242836107), .Z(n_247270467));
	notech_and4 i_129748484(.A(n_58055), .B(n_246970464), .C(n_246770462), .D
		(n_217370173), .Z(n_247170466));
	notech_ao4 i_129348488(.A(n_32186), .B(n_33297), .C(n_248736166), .D(nbus_11271
		[18]), .Z(n_246970464));
	notech_ao4 i_129548486(.A(n_57370), .B(\nbus_11290[18] ), .C(n_57325), .D
		(n_5436), .Z(n_246770462));
	notech_and4 i_130248479(.A(n_246470459), .B(n_246170457), .C(n_217770176
		), .D(n_218170179), .Z(n_246670461));
	notech_ao4 i_129848483(.A(n_60453), .B(n_31526), .C(n_385264383), .D(n_31491
		), .Z(n_246470459));
	notech_ao4 i_130048481(.A(n_58100), .B(n_319825274), .C(n_235370349), .D
		(n_242836107), .Z(n_246170457));
	notech_ao4 i_449721(.A(n_28240), .B(nbus_11273[3]), .C(n_331360941), .D(\nbus_11290[3] 
		), .Z(n_246070456));
	notech_and4 i_199047803(.A(n_245770453), .B(n_245670452), .C(n_245470450
		), .D(n_245370449), .Z(n_245970455));
	notech_ao4 i_198447809(.A(n_309771080), .B(n_33166), .C(n_100542446), .D
		(n_309671079), .Z(n_245770453));
	notech_ao4 i_198547808(.A(n_58042), .B(n_31479), .C(n_31514), .D(n_318971160
		), .Z(n_245670452));
	notech_ao4 i_198747806(.A(n_318871159), .B(n_33298), .C(n_61099), .D(n_30871
		), .Z(n_245470450));
	notech_ao4 i_198847805(.A(n_321271180), .B(n_337261000), .C(n_30326), .D
		(n_33299), .Z(n_245370449));
	notech_and4 i_199747796(.A(n_245070446), .B(n_244970445), .C(n_244770443
		), .D(n_244670442), .Z(n_245270448));
	notech_ao4 i_199147802(.A(n_249970494), .B(n_325260880), .C(n_249870493)
		, .D(n_325360881), .Z(n_245070446));
	notech_ao4 i_199247801(.A(n_262170616), .B(n_324960877), .C(n_57441), .D
		(n_325160879), .Z(n_244970445));
	notech_ao4 i_199447799(.A(n_243270428), .B(n_325460882), .C(n_243170427)
		, .D(n_325660884), .Z(n_244770443));
	notech_ao4 i_199547798(.A(n_242970425), .B(n_325560883), .C(n_242870424)
		, .D(n_325760885), .Z(n_244670442));
	notech_and4 i_200447789(.A(n_244370439), .B(n_244270438), .C(n_244070436
		), .D(n_243970435), .Z(n_244570441));
	notech_ao4 i_199847795(.A(n_309771080), .B(n_33165), .C(n_100242443), .D
		(n_309671079), .Z(n_244370439));
	notech_ao4 i_199947794(.A(n_58042), .B(n_31480), .C(n_318971160), .D(n_31515
		), .Z(n_244270438));
	notech_ao4 i_200147792(.A(n_318871159), .B(n_33300), .C(n_61097), .D(n_30872
		), .Z(n_244070436));
	notech_ao4 i_200247791(.A(n_336060988), .B(n_321271180), .C(n_30326), .D
		(n_33301), .Z(n_243970435));
	notech_and4 i_201147782(.A(n_243670432), .B(n_243570431), .C(n_243370429
		), .D(n_243070426), .Z(n_243870434));
	notech_ao4 i_200547788(.A(n_324660874), .B(n_249970494), .C(n_324560873)
		, .D(n_249870493), .Z(n_243670432));
	notech_ao4 i_200647787(.A(n_324160869), .B(n_262170616), .C(n_324060868)
		, .D(n_57441), .Z(n_243570431));
	notech_ao4 i_200847785(.A(n_324760875), .B(n_243270428), .C(n_324260870)
		, .D(n_243170427), .Z(n_243370429));
	notech_or2 i_849717(.A(n_262170616), .B(n_32304), .Z(n_243270428));
	notech_or2 i_949716(.A(n_57441), .B(n_32304), .Z(n_243170427));
	notech_ao4 i_200947784(.A(n_324360871), .B(n_242970425), .C(n_324460872)
		, .D(n_242870424), .Z(n_243070426));
	notech_or2 i_1049715(.A(n_262170616), .B(n_57449), .Z(n_242970425));
	notech_or2 i_1149714(.A(n_57441), .B(n_57449), .Z(n_242870424));
	notech_and4 i_201647777(.A(n_242570421), .B(n_242370419), .C(n_221770214
		), .D(n_222070217), .Z(n_242770423));
	notech_ao4 i_201247781(.A(n_309971082), .B(\nbus_11283[16] ), .C(n_310671088
		), .D(\nbus_11290[16] ), .Z(n_242570421));
	notech_ao4 i_201447779(.A(n_311771098), .B(n_33199), .C(n_318971160), .D
		(n_31524), .Z(n_242370419));
	notech_and4 i_202147772(.A(n_242070416), .B(n_241870414), .C(n_222370220
		), .D(n_222670223), .Z(n_242270418));
	notech_ao4 i_201747776(.A(n_311471096), .B(n_31489), .C(n_61097), .D(n_30882
		), .Z(n_242070416));
	notech_ao4 i_201947774(.A(n_320051171), .B(n_311571097), .C(n_240370399)
		, .D(n_311271094), .Z(n_241870414));
	notech_ao4 i_202247771(.A(n_57122), .B(n_31787), .C(n_33302), .D(n_57616
		), .Z(n_241570411));
	notech_ao4 i_202347770(.A(n_31755), .B(n_57141), .C(n_57157), .D(n_33303
		), .Z(n_241470410));
	notech_and2 i_202747766(.A(n_241270408), .B(n_241170407), .Z(n_241370409
		));
	notech_ao4 i_202547768(.A(n_31851), .B(n_57168), .C(n_32012), .D(n_30590
		), .Z(n_241270408));
	notech_ao4 i_202647767(.A(n_57192), .B(n_31723), .C(n_30679), .D(n_31948
		), .Z(n_241170407));
	notech_and4 i_203547758(.A(n_240870404), .B(n_240770403), .C(n_240570401
		), .D(n_240470400), .Z(n_241070406));
	notech_ao4 i_202947764(.A(n_31691), .B(n_57062), .C(n_30473), .D(n_31819
		), .Z(n_240870404));
	notech_ao4 i_203047763(.A(n_31883), .B(n_57091), .C(n_57103), .D(n_31588
		), .Z(n_240770403));
	notech_ao4 i_203247761(.A(n_58702), .B(n_31980), .C(n_31915), .D(n_59100
		), .Z(n_240570401));
	notech_ao4 i_203347760(.A(n_57218), .B(n_31424), .C(n_31659), .D(n_57230
		), .Z(n_240470400));
	notech_nand2 i_2549748(.A(opc_10[16]), .B(n_63782), .Z(n_240370399));
	notech_and4 i_204047753(.A(n_240070396), .B(n_239870394), .C(n_224570242
		), .D(n_224870245), .Z(n_240270398));
	notech_ao4 i_203647757(.A(n_309971082), .B(\nbus_11283[17] ), .C(n_310671088
		), .D(\nbus_11290[17] ), .Z(n_240070396));
	notech_ao4 i_203847755(.A(n_311771098), .B(n_33200), .C(n_318971160), .D
		(n_31525), .Z(n_239870394));
	notech_and4 i_204547748(.A(n_239570391), .B(n_239370389), .C(n_225170248
		), .D(n_225470251), .Z(n_239770393));
	notech_ao4 i_204147752(.A(n_311471096), .B(n_31490), .C(n_61097), .D(n_30883
		), .Z(n_239570391));
	notech_ao4 i_204347750(.A(n_319951172), .B(n_311571097), .C(n_237870374)
		, .D(n_311271094), .Z(n_239370389));
	notech_ao4 i_204647747(.A(n_57122), .B(n_31788), .C(n_57616), .D(n_33304
		), .Z(n_239070386));
	notech_ao4 i_204747746(.A(n_57141), .B(n_31756), .C(n_57157), .D(n_33305
		), .Z(n_238970385));
	notech_and2 i_205147742(.A(n_238770383), .B(n_238670382), .Z(n_238870384
		));
	notech_ao4 i_204947744(.A(n_57168), .B(n_31852), .C(n_30590), .D(n_32013
		), .Z(n_238770383));
	notech_ao4 i_205047743(.A(n_57192), .B(n_31724), .C(n_30679), .D(n_31949
		), .Z(n_238670382));
	notech_and4 i_205947734(.A(n_238370379), .B(n_238270378), .C(n_238070376
		), .D(n_237970375), .Z(n_238570381));
	notech_ao4 i_205347740(.A(n_57062), .B(n_31692), .C(n_30473), .D(n_31820
		), .Z(n_238370379));
	notech_ao4 i_205447739(.A(n_57091), .B(n_31884), .C(n_57103), .D(n_31589
		), .Z(n_238270378));
	notech_ao4 i_205647737(.A(n_58701), .B(n_31981), .C(n_59099), .D(n_31916
		), .Z(n_238070376));
	notech_ao4 i_205747736(.A(n_57218), .B(n_31425), .C(n_57230), .D(n_31660
		), .Z(n_237970375));
	notech_nand2 i_2649747(.A(opc_10[17]), .B(n_63764), .Z(n_237870374));
	notech_and4 i_206447729(.A(n_237570371), .B(n_237370369), .C(n_227370270
		), .D(n_227670273), .Z(n_237770373));
	notech_ao4 i_206047733(.A(n_309971082), .B(\nbus_11283[18] ), .C(n_310671088
		), .D(\nbus_11290[18] ), .Z(n_237570371));
	notech_ao4 i_206247731(.A(n_311771098), .B(n_33201), .C(n_318971160), .D
		(n_31526), .Z(n_237370369));
	notech_and4 i_206947724(.A(n_237070366), .B(n_236870364), .C(n_227970276
		), .D(n_228270279), .Z(n_237270368));
	notech_ao4 i_206547728(.A(n_311471096), .B(n_31491), .C(n_61097), .D(n_30884
		), .Z(n_237070366));
	notech_ao4 i_206747726(.A(n_319825274), .B(n_311571097), .C(n_235370349)
		, .D(n_311271094), .Z(n_236870364));
	notech_ao4 i_207047723(.A(n_57122), .B(n_31789), .C(n_57616), .D(n_33306
		), .Z(n_236570361));
	notech_ao4 i_207147722(.A(n_57136), .B(n_31757), .C(n_57158), .D(n_33307
		), .Z(n_236470360));
	notech_and2 i_207547718(.A(n_236270358), .B(n_236170357), .Z(n_236370359
		));
	notech_ao4 i_207347720(.A(n_57168), .B(n_31853), .C(n_30590), .D(n_32014
		), .Z(n_236270358));
	notech_ao4 i_207447719(.A(n_57192), .B(n_31725), .C(n_30679), .D(n_31950
		), .Z(n_236170357));
	notech_and4 i_208347710(.A(n_235870354), .B(n_235770353), .C(n_235570351
		), .D(n_235470350), .Z(n_236070356));
	notech_ao4 i_207747716(.A(n_57062), .B(n_31693), .C(n_30473), .D(n_31821
		), .Z(n_235870354));
	notech_ao4 i_207847715(.A(n_57091), .B(n_31885), .C(n_57103), .D(n_31590
		), .Z(n_235770353));
	notech_ao4 i_208047713(.A(n_58701), .B(n_31982), .C(n_59099), .D(n_31917
		), .Z(n_235570351));
	notech_ao4 i_208147712(.A(n_57218), .B(n_31426), .C(n_57230), .D(n_31661
		), .Z(n_235470350));
	notech_nand2 i_2749746(.A(opc_10[18]), .B(n_63782), .Z(n_235370349));
	notech_and4 i_208847705(.A(n_235070346), .B(n_234870344), .C(n_230170298
		), .D(n_230470301), .Z(n_235270348));
	notech_ao4 i_208447709(.A(n_309971082), .B(\nbus_11283[19] ), .C(n_310671088
		), .D(\nbus_11290[19] ), .Z(n_235070346));
	notech_ao4 i_208647707(.A(n_311771098), .B(n_33202), .C(n_318971160), .D
		(n_31527), .Z(n_234870344));
	notech_and4 i_209347700(.A(n_234570341), .B(n_234370339), .C(n_230770304
		), .D(n_231070307), .Z(n_234770343));
	notech_ao4 i_208947704(.A(n_311471096), .B(n_31492), .C(n_61097), .D(n_30885
		), .Z(n_234570341));
	notech_ao4 i_209147702(.A(n_319725273), .B(n_311571097), .C(n_232870324)
		, .D(n_311271094), .Z(n_234370339));
	notech_ao4 i_209447699(.A(n_57122), .B(n_31790), .C(n_57616), .D(n_33308
		), .Z(n_234070336));
	notech_ao4 i_209547698(.A(n_57136), .B(n_31758), .C(n_57157), .D(n_33309
		), .Z(n_233970335));
	notech_and2 i_209947694(.A(n_233770333), .B(n_233670332), .Z(n_233870334
		));
	notech_ao4 i_209747696(.A(n_57168), .B(n_31854), .C(n_57178), .D(n_32015
		), .Z(n_233770333));
	notech_ao4 i_209847695(.A(n_57192), .B(n_31726), .C(n_30679), .D(n_31951
		), .Z(n_233670332));
	notech_and4 i_210747686(.A(n_233370329), .B(n_233270328), .C(n_233070326
		), .D(n_232970325), .Z(n_233570331));
	notech_ao4 i_210147692(.A(n_57062), .B(n_31694), .C(n_57072), .D(n_31822
		), .Z(n_233370329));
	notech_ao4 i_210247691(.A(n_57091), .B(n_31886), .C(n_58701), .D(n_31983
		), .Z(n_233270328));
	notech_ao4 i_210447689(.A(n_59099), .B(n_31918), .C(n_57218), .D(n_31427
		), .Z(n_233070326));
	notech_ao4 i_210547688(.A(n_57230), .B(n_31662), .C(n_57103), .D(n_31591
		), .Z(n_232970325));
	notech_nand2 i_2849745(.A(opc_10[19]), .B(n_63782), .Z(n_232870324));
	notech_nand2 i_104448709(.A(\add_len_pc[19] ), .B(n_5680), .Z(n_231070307
		));
	notech_nand3 i_104748706(.A(n_2026), .B(n_6780), .C(n_32388), .Z(n_230770304
		));
	notech_or2 i_105048703(.A(n_5356), .B(n_311871099), .Z(n_230470301));
	notech_or2 i_105348700(.A(n_319071161), .B(nbus_11271[19]), .Z(n_230170298
		));
	notech_nand2 i_101648737(.A(\add_len_pc[18] ), .B(n_5680), .Z(n_228270279
		));
	notech_nand3 i_101948734(.A(n_2026), .B(n_6779), .C(n_32388), .Z(n_227970276
		));
	notech_or2 i_102248731(.A(n_5436), .B(n_311871099), .Z(n_227670273));
	notech_or2 i_102548728(.A(n_319071161), .B(nbus_11271[18]), .Z(n_227370270
		));
	notech_nand2 i_98848765(.A(\add_len_pc[17] ), .B(n_5680), .Z(n_225470251
		));
	notech_nand3 i_99148762(.A(n_2026), .B(n_6778), .C(n_32388), .Z(n_225170248
		));
	notech_or2 i_99448759(.A(n_5397), .B(n_311871099), .Z(n_224870245));
	notech_or2 i_99748756(.A(n_319071161), .B(nbus_11271[17]), .Z(n_224570242
		));
	notech_nand2 i_96048793(.A(\add_len_pc[16] ), .B(n_5680), .Z(n_222670223
		));
	notech_nand3 i_96348790(.A(n_2026), .B(n_6777), .C(n_32388), .Z(n_222370220
		));
	notech_or2 i_96648787(.A(n_5444), .B(n_311871099), .Z(n_222070217));
	notech_or2 i_96948784(.A(n_319071161), .B(nbus_11271[16]), .Z(n_221770214
		));
	notech_nand2 i_12749603(.A(sav_ecx[18]), .B(n_61870), .Z(n_218170179));
	notech_or2 i_13049600(.A(n_57326), .B(n_33201), .Z(n_217770176));
	notech_or2 i_13349597(.A(n_57369), .B(\nbus_11283[18] ), .Z(n_217370173)
		);
	notech_nand2 i_10549625(.A(sav_ecx[16]), .B(n_61870), .Z(n_216870168));
	notech_or2 i_10849622(.A(n_57326), .B(n_33199), .Z(n_216570165));
	notech_or2 i_11149619(.A(n_57369), .B(\nbus_11283[16] ), .Z(n_216270162)
		);
	notech_or4 i_8849641(.A(n_60175), .B(n_380764338), .C(nbus_11273[3]), .D
		(n_32241), .Z(n_215770157));
	notech_or2 i_9749632(.A(n_381164342), .B(n_31476), .Z(n_214770148));
	notech_and4 i_201551079(.A(n_211970121), .B(n_211770119), .C(n_211670118
		), .D(n_212270124), .Z(n_212470126));
	notech_and3 i_201251082(.A(n_58055), .B(n_212170123), .C(n_197569998), .Z
		(n_212270124));
	notech_ao4 i_200851086(.A(n_57369), .B(\nbus_11283[22] ), .C(n_248736166
		), .D(nbus_11271[22]), .Z(n_212170123));
	notech_ao4 i_201151083(.A(n_61097), .B(n_30774), .C(n_385264383), .D(n_31496
		), .Z(n_211970121));
	notech_ao4 i_201051084(.A(n_60453), .B(n_31530), .C(n_57326), .D(n_33284
		), .Z(n_211770119));
	notech_ao4 i_200951085(.A(n_59464), .B(n_57325), .C(n_57370), .D(\nbus_11290[22] 
		), .Z(n_211670118));
	notech_and4 i_174951341(.A(n_210770114), .B(n_210670113), .C(n_210470111
		), .D(n_210370110), .Z(n_211470116));
	notech_ao4 i_174651344(.A(n_31500), .B(n_58083), .C(n_324178250), .D(n_33171
		), .Z(n_210770114));
	notech_ao4 i_174551345(.A(n_324278251), .B(n_106826395), .C(n_57217), .D
		(\nbus_11290[24] ), .Z(n_210670113));
	notech_ao4 i_174451346(.A(n_57213), .B(\nbus_11283[24] ), .C(n_301822043
		), .D(nbus_11271[24]), .Z(n_210470111));
	notech_and2 i_174351347(.A(n_5774), .B(n_443068014), .Z(n_210370110));
	notech_nand3 i_48152594(.A(n_208970101), .B(n_208870100), .C(n_209970106
		), .Z(n_210070107));
	notech_and3 i_48052595(.A(n_209770104), .B(n_209570103), .C(n_196369986)
		, .Z(n_209970106));
	notech_ao4 i_47452601(.A(n_309971082), .B(n_58393), .C(n_319071161), .D(nbus_11271
		[20]), .Z(n_209770104));
	notech_ao4 i_47752598(.A(n_311471096), .B(n_31493), .C(n_318871159), .D(n_33293
		), .Z(n_209570103));
	notech_ao4 i_47652599(.A(n_318971160), .B(n_31528), .C(n_311771098), .D(n_33292
		), .Z(n_208970101));
	notech_ao4 i_47552600(.A(n_59466), .B(n_311871099), .C(n_58857), .D(n_310671088
		), .Z(n_208870100));
	notech_ao4 i_45552620(.A(n_57230), .B(n_31663), .C(n_57218), .D(n_31428)
		, .Z(n_208570097));
	notech_ao4 i_45452621(.A(n_59099), .B(n_31919), .C(n_58701), .D(n_31984)
		, .Z(n_208470096));
	notech_and2 i_45852617(.A(n_208270094), .B(n_208070093), .Z(n_208370095)
		);
	notech_ao4 i_45352622(.A(n_57103), .B(n_31592), .C(n_57086), .D(n_31887)
		, .Z(n_208270094));
	notech_ao4 i_45252623(.A(n_57072), .B(n_31823), .C(n_57062), .D(n_31695)
		, .Z(n_208070093));
	notech_and4 i_46052615(.A(n_207770090), .B(n_207670089), .C(n_207470087)
		, .D(n_207370086), .Z(n_207970092));
	notech_ao4 i_45152624(.A(n_30679), .B(n_31952), .C(n_57192), .D(n_31727)
		, .Z(n_207770090));
	notech_ao4 i_45052625(.A(n_57178), .B(n_32016), .C(n_57168), .D(n_31855)
		, .Z(n_207670089));
	notech_ao4 i_44952626(.A(n_57157), .B(n_33291), .C(n_57136), .D(n_31759)
		, .Z(n_207470087));
	notech_ao4 i_44852627(.A(n_57609), .B(n_33290), .C(n_57117), .D(n_31791)
		, .Z(n_207370086));
	notech_nand3 i_42852647(.A(n_206470077), .B(n_206370076), .C(n_206970082
		), .Z(n_207070083));
	notech_and3 i_42752648(.A(n_206770080), .B(n_206670079), .C(n_193569958)
		, .Z(n_206970082));
	notech_ao4 i_42152654(.A(n_309971082), .B(n_58402), .C(n_319071161), .D(nbus_11271
		[21]), .Z(n_206770080));
	notech_ao4 i_42452651(.A(n_311471096), .B(n_31494), .C(n_318871159), .D(n_33289
		), .Z(n_206670079));
	notech_ao4 i_42352652(.A(n_318971160), .B(n_31529), .C(n_311771098), .D(n_33288
		), .Z(n_206470077));
	notech_ao4 i_42252653(.A(n_59465), .B(n_311871099), .C(n_310671088), .D(n_58884
		), .Z(n_206370076));
	notech_ao4 i_40252673(.A(n_31664), .B(n_57230), .C(n_31429), .D(n_57218)
		, .Z(n_206070073));
	notech_ao4 i_40152674(.A(n_31920), .B(n_59099), .C(n_58701), .D(n_31985)
		, .Z(n_205970072));
	notech_and2 i_40552670(.A(n_205770070), .B(n_205670069), .Z(n_205870071)
		);
	notech_ao4 i_40052675(.A(n_31593), .B(n_57103), .C(n_31888), .D(n_57086)
		, .Z(n_205770070));
	notech_ao4 i_39952676(.A(n_31824), .B(n_57072), .C(n_31696), .D(n_57062)
		, .Z(n_205670069));
	notech_and4 i_40752668(.A(n_205370066), .B(n_205270065), .C(n_204970063)
		, .D(n_204870062), .Z(n_205570068));
	notech_ao4 i_39852677(.A(n_30679), .B(n_31953), .C(n_57192), .D(n_31728)
		, .Z(n_205370066));
	notech_ao4 i_39752678(.A(n_57178), .B(n_32017), .C(n_31856), .D(n_57168)
		, .Z(n_205270065));
	notech_ao4 i_39652679(.A(n_57157), .B(n_33287), .C(n_31760), .D(n_57136)
		, .Z(n_204970063));
	notech_ao4 i_39552680(.A(n_57609), .B(n_33286), .C(n_31792), .D(n_57117)
		, .Z(n_204870062));
	notech_nand3 i_37552700(.A(n_203870053), .B(n_203770052), .C(n_204470058
		), .Z(n_204570059));
	notech_and3 i_37452701(.A(n_204270056), .B(n_204170055), .C(n_190769930)
		, .Z(n_204470058));
	notech_ao4 i_36852707(.A(\nbus_11283[22] ), .B(n_309971082), .C(nbus_11271
		[22]), .D(n_319071161), .Z(n_204270056));
	notech_ao4 i_37152704(.A(n_311471096), .B(n_31496), .C(n_318871159), .D(n_33285
		), .Z(n_204170055));
	notech_ao4 i_37052705(.A(n_318971160), .B(n_31530), .C(n_311771098), .D(n_33284
		), .Z(n_203870053));
	notech_ao4 i_36952706(.A(n_59464), .B(n_311871099), .C(n_310671088), .D(\nbus_11290[22] 
		), .Z(n_203770052));
	notech_ao4 i_34952726(.A(n_57230), .B(n_31665), .C(n_57218), .D(n_31430)
		, .Z(n_203170049));
	notech_ao4 i_34852727(.A(n_59100), .B(n_31921), .C(n_58701), .D(n_31986)
		, .Z(n_203070048));
	notech_and2 i_35252723(.A(n_202870046), .B(n_202770045), .Z(n_202970047)
		);
	notech_ao4 i_34752728(.A(n_57103), .B(n_31594), .C(n_57086), .D(n_31889)
		, .Z(n_202870046));
	notech_ao4 i_34652729(.A(n_57072), .B(n_31825), .C(n_57062), .D(n_31697)
		, .Z(n_202770045));
	notech_and4 i_35452721(.A(n_202270042), .B(n_202170041), .C(n_201770039)
		, .D(n_201670038), .Z(n_202470044));
	notech_ao4 i_34552730(.A(n_30679), .B(n_31954), .C(n_57192), .D(n_31729)
		, .Z(n_202270042));
	notech_ao4 i_34452731(.A(n_57178), .B(n_32018), .C(n_57168), .D(n_31857)
		, .Z(n_202170041));
	notech_ao4 i_34352732(.A(n_57157), .B(n_33283), .C(n_57136), .D(n_31761)
		, .Z(n_201770039));
	notech_ao4 i_34252733(.A(n_57609), .B(n_33282), .C(n_57117), .D(n_31793)
		, .Z(n_201670038));
	notech_nand3 i_32252753(.A(n_200770029), .B(n_200670028), .C(n_201270034
		), .Z(n_201370035));
	notech_and3 i_32152754(.A(n_201070032), .B(n_200970031), .C(n_187969902)
		, .Z(n_201270034));
	notech_ao4 i_31552760(.A(n_309971082), .B(n_58420), .C(n_319071161), .D(nbus_11271
		[23]), .Z(n_201070032));
	notech_ao4 i_31852757(.A(n_311471096), .B(n_31499), .C(n_318871159), .D(n_33281
		), .Z(n_200970031));
	notech_ao4 i_31752758(.A(n_318971160), .B(n_31531), .C(n_311771098), .D(n_33170
		), .Z(n_200770029));
	notech_ao4 i_31652759(.A(n_311871099), .B(n_109226419), .C(n_310671088),
		 .D(n_58902), .Z(n_200670028));
	notech_nand3 i_26952806(.A(n_199670019), .B(n_199570018), .C(n_200170024
		), .Z(n_200270025));
	notech_and3 i_26852807(.A(n_199970022), .B(n_199870021), .C(n_186769890)
		, .Z(n_200170024));
	notech_ao4 i_26252813(.A(n_309971082), .B(\nbus_11283[24] ), .C(n_319071161
		), .D(nbus_11271[24]), .Z(n_199970022));
	notech_ao4 i_26552810(.A(n_311471096), .B(n_31500), .C(n_318871159), .D(n_33280
		), .Z(n_199870021));
	notech_ao4 i_26452811(.A(n_56992), .B(n_31532), .C(n_311771098), .D(n_33171
		), .Z(n_199670019));
	notech_ao4 i_26352812(.A(n_311871099), .B(n_106826395), .C(n_310671088),
		 .D(\nbus_11290[24] ), .Z(n_199570018));
	notech_nand3 i_24652829(.A(n_198670009), .B(n_198570008), .C(n_199170014
		), .Z(n_199270015));
	notech_and3 i_24552830(.A(n_198970012), .B(n_198870011), .C(n_185469878)
		, .Z(n_199170014));
	notech_ao4 i_23952836(.A(n_309971082), .B(\nbus_11283[25] ), .C(n_319071161
		), .D(nbus_11271[25]), .Z(n_198970012));
	notech_ao4 i_24252833(.A(n_311471096), .B(n_31501), .C(n_57034), .D(n_33279
		), .Z(n_198870011));
	notech_ao4 i_24152834(.A(n_56992), .B(n_31533), .C(n_311771098), .D(n_33172
		), .Z(n_198670009));
	notech_ao4 i_24052835(.A(n_311871099), .B(n_101026337), .C(n_310671088),
		 .D(\nbus_11290[25] ), .Z(n_198570008));
	notech_nand3 i_2317013(.A(n_212470126), .B(n_198470007), .C(n_197469997)
		, .Z(n_12067));
	notech_nao3 i_200651088(.A(opc_10[22]), .B(n_63782), .C(n_242836107), .Z
		(n_198470007));
	notech_nao3 i_199651098(.A(\regs_1_0[22] ), .B(n_19680), .C(n_57006), .Z
		(n_197569998));
	notech_or2 i_200551089(.A(n_3464), .B(n_58100), .Z(n_197469997));
	notech_nand3 i_2521847(.A(n_211470116), .B(n_197369996), .C(n_196669989)
		, .Z(n_12788));
	notech_nao3 i_174251348(.A(n_63792), .B(opc_10[24]), .C(n_298922014), .Z
		(n_197369996));
	notech_or4 i_174151349(.A(n_340461032), .B(n_2845), .C(n_444168025), .D(n_364628688
		), .Z(n_196669989));
	notech_or4 i_2120691(.A(n_196569988), .B(n_196469987), .C(n_210070107), 
		.D(n_195469977), .Z(n_20014));
	notech_ao3 i_47352602(.A(opc_10[20]), .B(n_63734), .C(n_311271094), .Z(n_196569988
		));
	notech_and2 i_47152604(.A(n_3458), .B(n_5680), .Z(n_196469987));
	notech_nand2 i_47052605(.A(sav_epc[20]), .B(n_61870), .Z(n_196369986));
	notech_nor2 i_47252603(.A(n_346771358), .B(n_311571097), .Z(n_195469977)
		);
	notech_or4 i_2220692(.A(n_193769960), .B(n_193669959), .C(n_207070083), 
		.D(n_192669949), .Z(n_20020));
	notech_ao3 i_42052655(.A(opc_10[21]), .B(n_63782), .C(n_311271094), .Z(n_193769960
		));
	notech_and2 i_41852657(.A(n_3459), .B(n_5680), .Z(n_193669959));
	notech_nand2 i_41752658(.A(sav_epc[21]), .B(n_61866), .Z(n_193569958));
	notech_nor2 i_41952656(.A(n_3466), .B(n_311571097), .Z(n_192669949));
	notech_or4 i_2320693(.A(n_190969932), .B(n_190869931), .C(n_204570059), 
		.D(n_189869921), .Z(n_20026));
	notech_ao3 i_36752708(.A(opc_10[22]), .B(n_63764), .C(n_311271094), .Z(n_190969932
		));
	notech_and2 i_36552710(.A(n_3460), .B(n_5680), .Z(n_190869931));
	notech_nand2 i_36452711(.A(sav_epc[22]), .B(n_61866), .Z(n_190769930));
	notech_nor2 i_36652709(.A(n_3464), .B(n_311571097), .Z(n_189869921));
	notech_or4 i_2420694(.A(n_188169904), .B(n_188069903), .C(n_201370035), 
		.D(n_187069893), .Z(n_20032));
	notech_ao3 i_31452761(.A(n_63792), .B(opc_10[23]), .C(n_311271094), .Z(n_188169904
		));
	notech_and2 i_31252763(.A(n_3461), .B(n_5680), .Z(n_188069903));
	notech_nand2 i_31152764(.A(sav_epc[23]), .B(n_61866), .Z(n_187969902));
	notech_nor2 i_31352762(.A(n_311571097), .B(n_363450925), .Z(n_187069893)
		);
	notech_or4 i_2520695(.A(n_186969892), .B(n_186869891), .C(n_200270025), 
		.D(n_185869881), .Z(n_20038));
	notech_ao3 i_26152814(.A(n_63792), .B(opc_10[24]), .C(n_311271094), .Z(n_186969892
		));
	notech_and2 i_26052815(.A(n_3462), .B(n_5680), .Z(n_186869891));
	notech_nand2 i_25852817(.A(sav_epc[24]), .B(n_61866), .Z(n_186769890));
	notech_nor2 i_25952816(.A(n_311571097), .B(n_364628688), .Z(n_185869881)
		);
	notech_or4 i_2620696(.A(n_185769880), .B(n_185569879), .C(n_199270015), 
		.D(n_183669869), .Z(n_20044));
	notech_ao3 i_23852837(.A(n_63792), .B(opc_10[25]), .C(n_311271094), .Z(n_185769880
		));
	notech_and2 i_23652839(.A(n_3463), .B(n_5680), .Z(n_185569879));
	notech_nand2 i_23552840(.A(sav_epc[25]), .B(n_61866), .Z(n_185469878));
	notech_nor2 i_23752838(.A(n_311571097), .B(n_363350926), .Z(n_183669869)
		);
	notech_and4 i_106254926(.A(n_58055), .B(n_182069854), .C(n_181869852), .D
		(n_157869616), .Z(n_182269856));
	notech_ao4 i_105854930(.A(n_32186), .B(n_33272), .C(n_248736166), .D(nbus_11271
		[26]), .Z(n_182069854));
	notech_ao4 i_106054928(.A(n_57370), .B(\nbus_11290[26] ), .C(n_57325), .D
		(n_5720), .Z(n_181869852));
	notech_and4 i_106754921(.A(n_181469849), .B(n_181269847), .C(n_158169619
		), .D(n_158469622), .Z(n_181669851));
	notech_ao4 i_106354925(.A(n_60454), .B(n_31534), .C(n_385264383), .D(n_31502
		), .Z(n_181469849));
	notech_ao4 i_106554923(.A(n_58100), .B(n_284231523), .C(n_175169787), .D
		(n_242836107), .Z(n_181269847));
	notech_and4 i_107254916(.A(n_58055), .B(n_180969844), .C(n_180769842), .D
		(n_158969627), .Z(n_181169846));
	notech_ao4 i_106854920(.A(n_32186), .B(n_33273), .C(n_248736166), .D(nbus_11271
		[27]), .Z(n_180969844));
	notech_ao4 i_107054918(.A(n_57370), .B(\nbus_11290[27] ), .C(n_57325), .D
		(n_5711), .Z(n_180769842));
	notech_and4 i_107754911(.A(n_180469839), .B(n_180269837), .C(n_159269630
		), .D(n_159569633), .Z(n_180669841));
	notech_ao4 i_107354915(.A(n_60454), .B(n_31535), .C(n_385264383), .D(n_31503
		), .Z(n_180469839));
	notech_ao4 i_107554913(.A(n_58100), .B(n_284131522), .C(n_172669762), .D
		(n_242836107), .Z(n_180269837));
	notech_and4 i_109154897(.A(n_58055), .B(n_179969834), .C(n_179669832), .D
		(n_160069638), .Z(n_180169836));
	notech_ao4 i_108754901(.A(n_32186), .B(n_33274), .C(n_248736166), .D(nbus_11271
		[29]), .Z(n_179969834));
	notech_ao4 i_108954899(.A(n_57370), .B(\nbus_11290[29] ), .C(n_4428), .D
		(n_57325), .Z(n_179669832));
	notech_and4 i_109654892(.A(n_179369829), .B(n_179169827), .C(n_160369641
		), .D(n_160669644), .Z(n_179569831));
	notech_ao4 i_109254896(.A(n_60454), .B(n_31537), .C(n_385264383), .D(n_31505
		), .Z(n_179369829));
	notech_ao4 i_109454894(.A(n_4387), .B(n_58100), .C(n_94229643), .D(n_242836107
		), .Z(n_179169827));
	notech_and4 i_128154709(.A(n_178869824), .B(n_178769823), .C(n_178569821
		), .D(n_178469820), .Z(n_179069826));
	notech_ao4 i_127554715(.A(n_178776847), .B(n_325760885), .C(n_178676846)
		, .D(n_325660884), .Z(n_178869824));
	notech_ao4 i_127654714(.A(n_178576845), .B(n_325460882), .C(n_178476844)
		, .D(n_325560883), .Z(n_178769823));
	notech_ao4 i_127854712(.A(n_31160), .B(n_56896), .C(n_200977065), .D(n_325360881
		), .Z(n_178569821));
	notech_ao4 i_127954711(.A(n_200877064), .B(n_325260880), .C(n_197877035)
		, .D(\nbus_11290[6] ), .Z(n_178469820));
	notech_ao4 i_128254708(.A(n_178376843), .B(n_324960877), .C(n_57289), .D
		(n_100542446), .Z(n_178169817));
	notech_ao4 i_128354707(.A(n_57432), .B(n_325160879), .C(n_58019), .D(n_31479
		), .Z(n_178069816));
	notech_and3 i_128854702(.A(n_177669812), .B(n_177869814), .C(n_162369661
		), .Z(n_177969815));
	notech_ao4 i_128554705(.A(n_245877510), .B(n_31514), .C(n_204977105), .D
		(n_33166), .Z(n_177869814));
	notech_ao4 i_128654704(.A(n_57157), .B(n_325060878), .C(n_57426), .D(n_156169599
		), .Z(n_177669812));
	notech_and4 i_172854268(.A(n_177369809), .B(n_177169807), .C(n_162669664
		), .D(n_162969667), .Z(n_177569811));
	notech_ao4 i_172454272(.A(n_309971082), .B(\nbus_11283[26] ), .C(n_310671088
		), .D(\nbus_11290[26] ), .Z(n_177369809));
	notech_ao4 i_172654270(.A(n_311771098), .B(n_33198), .C(n_56992), .D(n_31534
		), .Z(n_177169807));
	notech_and4 i_173354263(.A(n_176869804), .B(n_176669802), .C(n_163269670
		), .D(n_163569673), .Z(n_177069806));
	notech_ao4 i_172954267(.A(n_311471096), .B(n_31502), .C(n_61097), .D(n_30887
		), .Z(n_176869804));
	notech_ao4 i_173154265(.A(n_284231523), .B(n_311571097), .C(n_175169787)
		, .D(n_311271094), .Z(n_176669802));
	notech_ao4 i_173454262(.A(n_57117), .B(n_31797), .C(n_57609), .D(n_33275
		), .Z(n_176369799));
	notech_ao4 i_173554261(.A(n_57136), .B(n_31765), .C(n_57157), .D(n_33276
		), .Z(n_176269798));
	notech_and2 i_173954257(.A(n_176069796), .B(n_175969795), .Z(n_176169797
		));
	notech_ao4 i_173754259(.A(n_57168), .B(n_31861), .C(n_57178), .D(n_32022
		), .Z(n_176069796));
	notech_ao4 i_173854258(.A(n_57192), .B(n_31733), .C(n_30679), .D(n_31958
		), .Z(n_175969795));
	notech_and4 i_174754249(.A(n_175669792), .B(n_175569791), .C(n_175369789
		), .D(n_175269788), .Z(n_175869794));
	notech_ao4 i_174154255(.A(n_57062), .B(n_31701), .C(n_57072), .D(n_31829
		), .Z(n_175669792));
	notech_ao4 i_174254254(.A(n_57086), .B(n_31893), .C(n_57103), .D(n_31598
		), .Z(n_175569791));
	notech_ao4 i_174454252(.A(n_58701), .B(n_31990), .C(n_59100), .D(n_31925
		), .Z(n_175369789));
	notech_ao4 i_174554251(.A(n_57218), .B(n_31434), .C(n_57230), .D(n_31669
		), .Z(n_175269788));
	notech_nand2 i_1755925(.A(n_63792), .B(opc_10[26]), .Z(n_175169787));
	notech_and4 i_175254244(.A(n_174869784), .B(n_174669782), .C(n_165469692
		), .D(n_165769695), .Z(n_175069786));
	notech_ao4 i_174854248(.A(n_309971082), .B(\nbus_11283[27] ), .C(n_310671088
		), .D(\nbus_11290[27] ), .Z(n_174869784));
	notech_ao4 i_175054246(.A(n_311771098), .B(n_33195), .C(n_56992), .D(n_31535
		), .Z(n_174669782));
	notech_and4 i_175754239(.A(n_174369779), .B(n_174169777), .C(n_166069698
		), .D(n_166369701), .Z(n_174569781));
	notech_ao4 i_175354243(.A(n_311471096), .B(n_31503), .C(n_61097), .D(n_30888
		), .Z(n_174369779));
	notech_ao4 i_175554241(.A(n_284131522), .B(n_311571097), .C(n_172669762)
		, .D(n_311271094), .Z(n_174169777));
	notech_ao4 i_175854238(.A(n_57117), .B(n_31798), .C(n_57609), .D(n_33277
		), .Z(n_173869774));
	notech_ao4 i_175954237(.A(n_57136), .B(n_31766), .C(n_57157), .D(n_33278
		), .Z(n_173769773));
	notech_and2 i_176454233(.A(n_173569771), .B(n_173469770), .Z(n_173669772
		));
	notech_ao4 i_176254235(.A(n_57168), .B(n_31862), .C(n_57178), .D(n_32023
		), .Z(n_173569771));
	notech_ao4 i_176354234(.A(n_57192), .B(n_31734), .C(n_30679), .D(n_31959
		), .Z(n_173469770));
	notech_and4 i_177254225(.A(n_173169767), .B(n_173069766), .C(n_172869764
		), .D(n_172769763), .Z(n_173369769));
	notech_ao4 i_176654231(.A(n_57062), .B(n_31702), .C(n_57072), .D(n_31830
		), .Z(n_173169767));
	notech_ao4 i_176754230(.A(n_57086), .B(n_31894), .C(n_57103), .D(n_31599
		), .Z(n_173069766));
	notech_ao4 i_176954228(.A(n_58701), .B(n_31991), .C(n_59100), .D(n_31926
		), .Z(n_172869764));
	notech_ao4 i_177054227(.A(n_57218), .B(n_31435), .C(n_57230), .D(n_31670
		), .Z(n_172769763));
	notech_nand2 i_1855924(.A(opc_10[27]), .B(n_63760), .Z(n_172669762));
	notech_and4 i_177754220(.A(n_172369759), .B(n_172169757), .C(n_168269720
		), .D(n_168569723), .Z(n_172569761));
	notech_ao4 i_177354224(.A(n_309971082), .B(\nbus_11283[28] ), .C(n_310671088
		), .D(\nbus_11290[28] ), .Z(n_172369759));
	notech_ao4 i_177554222(.A(n_311771098), .B(n_33196), .C(n_56992), .D(n_31536
		), .Z(n_172169757));
	notech_and4 i_178254215(.A(n_171669754), .B(n_171469752), .C(n_168869726
		), .D(n_169169729), .Z(n_171869756));
	notech_ao4 i_177854219(.A(n_311471096), .B(n_31504), .C(n_61097), .D(n_30889
		), .Z(n_171669754));
	notech_ao4 i_178054217(.A(n_440082450), .B(n_311571097), .C(n_7636), .D(n_311271094
		), .Z(n_171469752));
	notech_and4 i_180154196(.A(n_171169749), .B(n_170969747), .C(n_169469732
		), .D(n_169769735), .Z(n_171369751));
	notech_ao4 i_179754200(.A(n_309971082), .B(\nbus_11283[29] ), .C(n_310671088
		), .D(\nbus_11290[29] ), .Z(n_171169749));
	notech_ao4 i_179954198(.A(n_311771098), .B(n_33197), .C(n_56992), .D(n_31537
		), .Z(n_170969747));
	notech_and4 i_180654191(.A(n_170669744), .B(n_170469742), .C(n_170069738
		), .D(n_170369741), .Z(n_170869746));
	notech_ao4 i_180254195(.A(n_311471096), .B(n_31505), .C(n_61097), .D(n_30892
		), .Z(n_170669744));
	notech_ao4 i_180454193(.A(n_4387), .B(n_311571097), .C(n_94229643), .D(n_311271094
		), .Z(n_170469742));
	notech_nand2 i_94255038(.A(\add_len_pc[29] ), .B(n_5680), .Z(n_170369741
		));
	notech_nand3 i_94555035(.A(n_2026), .B(n_6790), .C(n_32388), .Z(n_170069738
		));
	notech_or2 i_94855032(.A(n_4428), .B(n_311871099), .Z(n_169769735));
	notech_or2 i_95155029(.A(n_319071161), .B(nbus_11271[29]), .Z(n_169469732
		));
	notech_nand2 i_91455066(.A(\add_len_pc[28] ), .B(n_5680), .Z(n_169169729
		));
	notech_nand3 i_91755063(.A(n_2026), .B(n_6789), .C(n_32388), .Z(n_168869726
		));
	notech_or2 i_92055060(.A(n_4427), .B(n_311871099), .Z(n_168569723));
	notech_or2 i_92355057(.A(n_319071161), .B(nbus_11271[28]), .Z(n_168269720
		));
	notech_nand2 i_88455094(.A(\add_len_pc[27] ), .B(n_5680), .Z(n_166369701
		));
	notech_nand3 i_88755091(.A(n_2026), .B(n_6788), .C(n_32388), .Z(n_166069698
		));
	notech_or2 i_89055088(.A(n_5711), .B(n_311871099), .Z(n_165769695));
	notech_or2 i_89355085(.A(n_319071161), .B(nbus_11271[27]), .Z(n_165469692
		));
	notech_nand2 i_85055122(.A(\add_len_pc[26] ), .B(n_5680), .Z(n_163569673
		));
	notech_nand3 i_85355119(.A(n_6787), .B(n_2026), .C(n_32388), .Z(n_163269670
		));
	notech_or2 i_85655116(.A(n_5720), .B(n_311871099), .Z(n_162969667));
	notech_or2 i_85955113(.A(n_319071161), .B(nbus_11271[26]), .Z(n_162669664
		));
	notech_nand2 i_42255535(.A(n_4386), .B(opa[6]), .Z(n_162369661));
	notech_and2 i_42271558(.A(n_61286), .B(n_56734), .Z(n_116176227));
	notech_or4 i_49031(.A(n_124545737), .B(n_30312), .C(n_30311), .D(n_116176227
		), .Z(\nbus_11304[16] ));
	notech_nand3 i_8442(.A(n_19655), .B(n_30524), .C(n_61625), .Z(n_11335)
		);
	notech_or2 i_128466154(.A(n_57439), .B(n_27378), .Z(n_116576231));
	notech_nand2 i_1966137(.A(n_83839558), .B(n_328360911), .Z(n_116676232)
		);
	notech_or4 i_2966127(.A(n_338661014), .B(n_318160809), .C(n_285763759), 
		.D(n_192576983), .Z(n_116776233));
	notech_nor2 i_3066126(.A(n_376064291), .B(n_192576983), .Z(n_116876234)
		);
	notech_nand3 i_3166125(.A(n_61097), .B(n_61621), .C(read_data[0]), .Z(n_116976235
		));
	notech_ao3 i_6566091(.A(n_57027), .B(n_57213), .C(n_323878247), .Z(n_117076236
		));
	notech_and3 i_6666090(.A(n_57036), .B(n_323678245), .C(n_57217), .Z(n_117176237
		));
	notech_ao4 i_5866098(.A(n_32697), .B(n_31363), .C(n_30275), .D(n_220495876
		), .Z(n_117276238));
	notech_and2 i_5966097(.A(n_330060928), .B(n_329160919), .Z(n_117376239)
		);
	notech_mux2 i_5766099(.S(n_32243), .A(n_117876244), .B(n_117676242), .Z(n_117476240
		));
	notech_ao4 i_4166115(.A(n_60170), .B(n_59005), .C(n_30920), .D(n_27378),
		 .Z(n_117676242));
	notech_ao4 i_4066116(.A(n_60170), .B(nbus_11273[1]), .C(n_30919), .D(n_27378
		), .Z(n_117876244));
	notech_ao3 i_5566101(.A(n_279677807), .B(n_303378043), .C(n_192876986), 
		.Z(n_118176247));
	notech_and3 i_5666100(.A(n_279877809), .B(n_201077066), .C(n_280077811),
		 .Z(n_118276248));
	notech_nand3 i_60665562(.A(n_61099), .B(n_61621), .C(read_data[2]), .Z(n_118376249
		));
	notech_nand3 i_62265546(.A(n_61097), .B(n_61621), .C(read_data[4]), .Z(n_118476250
		));
	notech_nand3 i_63865530(.A(n_61099), .B(n_61621), .C(read_data[5]), .Z(n_118576251
		));
	notech_nand3 i_67065498(.A(n_61099), .B(n_61621), .C(read_data[7]), .Z(n_118676252
		));
	notech_ao3 i_5066106(.A(n_192676984), .B(n_57201), .C(n_116876234), .Z(n_118776253
		));
	notech_and3 i_5166105(.A(n_323278241), .B(n_116776233), .C(n_57200), .Z(n_118876254
		));
	notech_nao3 i_9366063(.A(n_63792), .B(opc_10[14]), .C(n_333978345), .Z(n_118976255
		));
	notech_or2 i_8866068(.A(n_58030), .B(n_31487), .Z(n_119676262));
	notech_or2 i_31065851(.A(n_336760995), .B(n_328760915), .Z(n_120176267)
		);
	notech_nao3 i_30765854(.A(n_1640), .B(n_2640), .C(n_163296016), .Z(n_120476270
		));
	notech_or4 i_30465857(.A(n_27379), .B(n_61935), .C(n_31611), .D(n_30549)
		, .Z(n_120776273));
	notech_nand2 i_34565816(.A(sav_esi[2]), .B(n_61866), .Z(n_122276288));
	notech_nand2 i_36065801(.A(sav_esi[4]), .B(n_61866), .Z(n_123776303));
	notech_nand2 i_37565786(.A(sav_esi[5]), .B(n_61866), .Z(n_125276318));
	notech_nand2 i_40865756(.A(sav_esi[7]), .B(n_61870), .Z(n_126776333));
	notech_or2 i_42265742(.A(n_336660994), .B(n_328860916), .Z(n_128476350)
		);
	notech_nand2 i_41565749(.A(opb[9]), .B(n_57129), .Z(n_129176357));
	notech_or2 i_50765660(.A(n_337561003), .B(nbus_11271[30]), .Z(n_129876364
		));
	notech_or2 i_50365663(.A(n_124726574), .B(n_33194), .Z(n_130176367));
	notech_or2 i_50065666(.A(n_328660914), .B(n_31506), .Z(n_130476370));
	notech_nand2 i_49665669(.A(sav_esi[30]), .B(n_61870), .Z(n_130776373));
	notech_or2 i_54565623(.A(n_58053), .B(n_31487), .Z(n_131676382));
	notech_ao3 i_56565603(.A(n_57392), .B(opd[30]), .C(n_57157), .Z(n_132576391
		));
	notech_or4 i_62165547(.A(n_28551), .B(n_30441), .C(n_61935), .D(n_31615)
		, .Z(n_132676392));
	notech_or4 i_63765531(.A(n_28551), .B(n_30441), .C(n_61935), .D(n_31616)
		, .Z(n_134176407));
	notech_or2 i_66965499(.A(n_331660944), .B(n_336060988), .Z(n_135676422)
		);
	notech_or4 i_86965299(.A(n_61935), .B(n_31624), .C(n_30319), .D(n_323578244
		), .Z(n_137576441));
	notech_nao3 i_86665302(.A(n_30300), .B(\opa_12[13] ), .C(n_376064291), .Z
		(n_137876444));
	notech_or4 i_86365305(.A(n_63698), .B(n_57387), .C(n_63782), .D(nbus_11273
		[13]), .Z(n_138176447));
	notech_nor2 i_88065288(.A(n_279977810), .B(nbus_11271[14]), .Z(n_138276448
		));
	notech_and4 i_87965289(.A(n_63774), .B(opc_10[14]), .C(n_29214), .D(n_30300
		), .Z(n_138576451));
	notech_nor2 i_87465294(.A(n_58029), .B(n_31487), .Z(n_139076456));
	notech_or2 i_766149(.A(n_27379), .B(n_30549), .Z(n_139176457));
	notech_or2 i_266150(.A(n_57439), .B(n_30549), .Z(n_139276458));
	notech_or4 i_1166145(.A(n_2383), .B(n_57439), .C(instrc[120]), .D(n_32161
		), .Z(n_139376459));
	notech_or2 i_1466142(.A(n_57439), .B(n_32243), .Z(n_139476460));
	notech_or4 i_1266144(.A(n_2383), .B(n_116576231), .C(instrc[120]), .D(n_32161
		), .Z(n_139576461));
	notech_nao3 i_1366143(.A(n_30549), .B(n_57461), .C(n_57439), .Z(n_139676462
		));
	notech_or4 i_2566131(.A(n_338661014), .B(n_169676762), .C(instrc[122]), 
		.D(n_32159), .Z(n_139876464));
	notech_nao3 i_2166135(.A(n_30319), .B(n_57627), .C(n_57666), .Z(n_139976465
		));
	notech_or2 i_2066136(.A(n_57666), .B(n_32252), .Z(n_140076466));
	notech_or4 i_2466132(.A(n_338661014), .B(n_57666), .C(instrc[122]), .D(n_32159
		), .Z(n_140176467));
	notech_ao4 i_175964433(.A(\nbus_11290[14] ), .B(n_118876254), .C(nbus_11273
		[14]), .D(n_118776253), .Z(n_140576471));
	notech_ao4 i_175864434(.A(n_323478243), .B(n_33215), .C(n_57609), .D(n_377064301
		), .Z(n_140776473));
	notech_ao4 i_175564437(.A(n_377164302), .B(n_334378349), .C(n_97342414),
		 .D(n_323378242), .Z(n_140976475));
	notech_or4 i_175764435(.A(n_138276448), .B(n_30558), .C(n_138576451), .D
		(n_30281), .Z(n_141276478));
	notech_ao4 i_175164441(.A(n_30474), .B(n_57609), .C(n_58029), .D(n_31486
		), .Z(n_141376479));
	notech_ao4 i_174964443(.A(\nbus_11290[13] ), .B(n_57238), .C(nbus_11273[
		13]), .D(n_57237), .Z(n_141576481));
	notech_and4 i_175364439(.A(n_141576481), .B(n_141376479), .C(n_137876444
		), .D(n_138176447), .Z(n_141776483));
	notech_ao4 i_174664446(.A(n_31497), .B(n_334378349), .C(n_375064281), .D
		(n_323378242), .Z(n_141876484));
	notech_ao4 i_174464448(.A(n_279977810), .B(nbus_11271[13]), .C(n_31498),
		 .D(n_334478350), .Z(n_142076486));
	notech_and4 i_174864444(.A(n_142076486), .B(n_141876484), .C(n_30468), .D
		(n_137576441), .Z(n_142276488));
	notech_ao4 i_156664626(.A(n_28259), .B(n_324760875), .C(n_28256), .D(n_324260870
		), .Z(n_142376489));
	notech_ao4 i_156564627(.A(n_28255), .B(n_324360871), .C(n_28258), .D(n_324460872
		), .Z(n_142476490));
	notech_ao4 i_156364629(.A(n_61099), .B(n_30841), .C(n_28260), .D(n_324160869
		), .Z(n_142676492));
	notech_ao4 i_156264630(.A(n_439367977), .B(n_324060868), .C(n_439467978)
		, .D(n_31480), .Z(n_142776493));
	notech_and4 i_156864624(.A(n_142776493), .B(n_142676492), .C(n_142476490
		), .D(n_142376489), .Z(n_142976495));
	notech_ao4 i_155964633(.A(n_439667980), .B(n_100242443), .C(n_439567979)
		, .D(n_33165), .Z(n_143076496));
	notech_ao4 i_155864634(.A(n_28252), .B(n_324660874), .C(n_28251), .D(n_324560873
		), .Z(n_143176497));
	notech_ao4 i_155664636(.A(n_333260960), .B(n_33435), .C(n_333360961), .D
		(n_33434), .Z(n_143376499));
	notech_and4 i_155764635(.A(n_28238), .B(n_143376499), .C(n_118676252), .D
		(n_135676422), .Z(n_143676502));
	notech_ao4 i_153864654(.A(n_28259), .B(n_31126), .C(n_28256), .D(n_31122
		), .Z(n_143876504));
	notech_ao4 i_153764655(.A(n_31125), .B(n_28255), .C(n_31123), .D(n_28258
		), .Z(n_143976505));
	notech_ao4 i_153564657(.A(n_61097), .B(n_30838), .C(n_28260), .D(n_31099
		), .Z(n_144176507));
	notech_ao4 i_153364658(.A(n_333260960), .B(n_33433), .C(n_333360961), .D
		(n_33432), .Z(n_144276508));
	notech_and4 i_154064652(.A(n_144276508), .B(n_144176507), .C(n_143976505
		), .D(n_143876504), .Z(n_144476510));
	notech_ao4 i_153064661(.A(n_331660944), .B(n_334960977), .C(n_439467978)
		, .D(n_31478), .Z(n_144576511));
	notech_ao4 i_152964662(.A(n_439567979), .B(n_33135), .C(n_439367977), .D
		(n_31098), .Z(n_144676512));
	notech_ao4 i_152664664(.A(n_31118), .B(n_28251), .C(n_439667980), .D(n_334860976
		), .Z(n_144876514));
	notech_and4 i_152864663(.A(n_28206), .B(n_144876514), .C(n_118576251), .D
		(n_134176407), .Z(n_145176517));
	notech_ao4 i_152264668(.A(n_28259), .B(n_31075), .C(n_28256), .D(n_31071
		), .Z(n_145376519));
	notech_ao4 i_152164669(.A(n_28255), .B(n_31074), .C(n_28258), .D(n_31072
		), .Z(n_145476520));
	notech_ao4 i_151964671(.A(n_61097), .B(n_30837), .C(n_28260), .D(n_31048
		), .Z(n_145676522));
	notech_ao4 i_151864672(.A(n_333260960), .B(n_33431), .C(n_333360961), .D
		(n_33430), .Z(n_145776523));
	notech_and4 i_152464666(.A(n_145776523), .B(n_145676522), .C(n_145476520
		), .D(n_145376519), .Z(n_145976525));
	notech_ao4 i_151564675(.A(n_331660944), .B(n_334760975), .C(n_439467978)
		, .D(n_31477), .Z(n_146076526));
	notech_ao4 i_151464676(.A(n_439567979), .B(n_33104), .C(n_439367977), .D
		(n_31047), .Z(n_146176527));
	notech_ao4 i_151264678(.A(n_28251), .B(n_31067), .C(n_439667980), .D(n_334660974
		), .Z(n_146376529));
	notech_and4 i_151364677(.A(n_28190), .B(n_146376529), .C(n_118476250), .D
		(n_132676392), .Z(n_146676532));
	notech_ao4 i_148164709(.A(n_5750), .B(n_302878038), .C(n_245877510), .D(n_31538
		), .Z(n_146976535));
	notech_ao4 i_148064710(.A(n_324678255), .B(\nbus_11283[30] ), .C(n_324578254
		), .D(\nbus_11290[30] ), .Z(n_147176537));
	notech_ao3 i_148364707(.A(n_146976535), .B(n_147176537), .C(n_132576391)
		, .Z(n_147276538));
	notech_ao4 i_147864712(.A(n_5758), .B(n_324478253), .C(n_324378252), .D(n_33194
		), .Z(n_147376539));
	notech_ao4 i_147764713(.A(n_302978039), .B(nbus_11271[30]), .C(n_318771158
		), .D(n_303078040), .Z(n_147476540));
	notech_ao4 i_146364727(.A(\nbus_11290[14] ), .B(n_118276248), .C(nbus_11273
		[14]), .D(n_118176247), .Z(n_147876544));
	notech_ao4 i_146264728(.A(n_57252), .B(n_33215), .C(n_57157), .D(n_377064301
		), .Z(n_148076546));
	notech_and3 i_146564725(.A(n_147876544), .B(n_148076546), .C(n_131676382
		), .Z(n_148176547));
	notech_ao4 i_146064730(.A(n_377164302), .B(n_200677062), .C(n_97342414),
		 .D(n_57317), .Z(n_148276548));
	notech_ao4 i_145964731(.A(n_245877510), .B(n_31522), .C(n_377264303), .D
		(n_200577061), .Z(n_148376549));
	notech_ao4 i_142864762(.A(n_330460932), .B(n_33429), .C(n_330560933), .D
		(n_33428), .Z(n_148576551));
	notech_ao4 i_142664764(.A(n_5750), .B(n_124126568), .C(n_57006), .D(n_31538
		), .Z(n_148776553));
	notech_and4 i_143064760(.A(n_148776553), .B(n_148576551), .C(n_130776373
		), .D(n_130476370), .Z(n_148976555));
	notech_ao4 i_142364767(.A(n_124626573), .B(\nbus_11283[30] ), .C(n_124526572
		), .D(\nbus_11290[30] ), .Z(n_149076556));
	notech_ao4 i_142164769(.A(n_318771158), .B(n_337661004), .C(n_5758), .D(n_124826575
		), .Z(n_149276558));
	notech_and4 i_142564765(.A(n_149276558), .B(n_149076556), .C(n_129876364
		), .D(n_130176367), .Z(n_149476560));
	notech_ao4 i_135864832(.A(n_330460932), .B(n_33427), .C(n_330560933), .D
		(n_33426), .Z(n_149576561));
	notech_ao4 i_135764833(.A(n_31482), .B(n_58025), .C(n_61097), .D(n_30814
		), .Z(n_149676562));
	notech_ao4 i_135564835(.A(n_57128), .B(nbus_11273[9]), .C(n_327060898), 
		.D(n_57394), .Z(n_149876564));
	notech_and4 i_136064830(.A(n_149876564), .B(n_149676562), .C(n_149576561
		), .D(n_129176357), .Z(n_150076566));
	notech_ao4 i_135264838(.A(n_99942440), .B(n_57275), .C(n_57274), .D(n_33168
		), .Z(n_150176567));
	notech_ao4 i_135164839(.A(n_334178347), .B(n_327260900), .C(n_327160899)
		, .D(n_334078346), .Z(n_150276568));
	notech_ao4 i_134964841(.A(n_57006), .B(n_31517), .C(n_327360901), .D(n_334278348
		), .Z(n_150476570));
	notech_and4 i_135464836(.A(n_150476570), .B(n_150276568), .C(n_150176567
		), .D(n_128476350), .Z(n_150676572));
	notech_ao4 i_134664844(.A(n_324760875), .B(n_139676462), .C(n_324260870)
		, .D(n_139476460), .Z(n_150776573));
	notech_ao4 i_134564845(.A(n_324460872), .B(n_139376459), .C(n_324360871)
		, .D(n_139576461), .Z(n_150876574));
	notech_ao4 i_134364847(.A(n_324560873), .B(n_139276458), .C(n_324660874)
		, .D(n_139176457), .Z(n_151076576));
	notech_ao4 i_134264848(.A(n_330560933), .B(n_33425), .C(n_324160869), .D
		(n_116576231), .Z(n_151176577));
	notech_and4 i_134864842(.A(n_151176577), .B(n_151076576), .C(n_150876574
		), .D(n_150776573), .Z(n_151376579));
	notech_ao4 i_133964851(.A(n_100242443), .B(n_57276), .C(n_330460932), .D
		(n_33424), .Z(n_151476580));
	notech_ao4 i_133864852(.A(n_324060868), .B(n_57439), .C(n_57277), .D(n_33165
		), .Z(n_151576581));
	notech_ao4 i_133664854(.A(n_58040), .B(n_31480), .C(n_336060988), .D(n_328760915
		), .Z(n_151776583));
	notech_and4 i_133764853(.A(n_28238), .B(n_118676252), .C(n_151776583), .D
		(n_126776333), .Z(n_151976585));
	notech_ao4 i_131864872(.A(n_31126), .B(n_139676462), .C(n_31122), .D(n_139476460
		), .Z(n_152176587));
	notech_ao4 i_131764873(.A(n_31123), .B(n_139376459), .C(n_31125), .D(n_139576461
		), .Z(n_152276588));
	notech_ao4 i_131564875(.A(n_31118), .B(n_139276458), .C(n_31119), .D(n_139176457
		), .Z(n_152476590));
	notech_ao4 i_131464876(.A(n_330560933), .B(n_33423), .C(n_31099), .D(n_116576231
		), .Z(n_152576591));
	notech_and4 i_132064870(.A(n_152576591), .B(n_152476590), .C(n_152276588
		), .D(n_152176587), .Z(n_152776593));
	notech_ao4 i_130964879(.A(n_334860976), .B(n_57276), .C(n_330460932), .D
		(n_33422), .Z(n_152876594));
	notech_ao4 i_130864880(.A(n_31098), .B(n_57439), .C(n_57277), .D(n_33135
		), .Z(n_152976595));
	notech_ao4 i_130664882(.A(n_58040), .B(n_31478), .C(n_334960977), .D(n_328760915
		), .Z(n_153176597));
	notech_and4 i_130764881(.A(n_28206), .B(n_118576251), .C(n_153176597), .D
		(n_125276318), .Z(n_153376599));
	notech_ao4 i_130264886(.A(n_31075), .B(n_139676462), .C(n_31071), .D(n_139476460
		), .Z(n_153576601));
	notech_ao4 i_130164887(.A(n_31072), .B(n_139376459), .C(n_31074), .D(n_139576461
		), .Z(n_153676602));
	notech_ao4 i_129964889(.A(n_31067), .B(n_139276458), .C(n_31068), .D(n_139176457
		), .Z(n_153876604));
	notech_ao4 i_129864890(.A(n_330560933), .B(n_33421), .C(n_31048), .D(n_116576231
		), .Z(n_153976605));
	notech_and4 i_130464884(.A(n_153976605), .B(n_153876604), .C(n_153676602
		), .D(n_153576601), .Z(n_154176607));
	notech_ao4 i_129564893(.A(n_334660974), .B(n_57276), .C(n_330460932), .D
		(n_33420), .Z(n_154276608));
	notech_ao4 i_129464894(.A(n_31047), .B(n_57439), .C(n_57277), .D(n_33104
		), .Z(n_154376609));
	notech_ao4 i_129264896(.A(n_58040), .B(n_31477), .C(n_334760975), .D(n_328760915
		), .Z(n_154576611));
	notech_and4 i_129364895(.A(n_28190), .B(n_118476250), .C(n_154576611), .D
		(n_123776303), .Z(n_154776613));
	notech_ao4 i_128864900(.A(n_326460892), .B(n_139676462), .C(n_326660894)
		, .D(n_139476460), .Z(n_154976615));
	notech_ao4 i_128764901(.A(n_326760895), .B(n_139376459), .C(n_326560893)
		, .D(n_139576461), .Z(n_155076616));
	notech_ao4 i_128364903(.A(n_326360891), .B(n_139276458), .C(n_326260890)
		, .D(n_139176457), .Z(n_155276618));
	notech_ao4 i_128264904(.A(n_330560933), .B(n_33419), .C(n_325960887), .D
		(n_116576231), .Z(n_155376619));
	notech_and4 i_129064898(.A(n_155376619), .B(n_155276618), .C(n_155076616
		), .D(n_154976615), .Z(n_155576621));
	notech_ao4 i_127964907(.A(n_100842449), .B(n_57276), .C(n_330460932), .D
		(n_33418), .Z(n_155676622));
	notech_ao4 i_127864908(.A(n_326160889), .B(n_57439), .C(n_57277), .D(n_33167
		), .Z(n_155776623));
	notech_ao4 i_127664910(.A(n_58040), .B(n_31474), .C(n_336160989), .D(n_328760915
		), .Z(n_155976625));
	notech_and4 i_127764909(.A(n_28158), .B(n_118376249), .C(n_155976625), .D
		(n_122276288), .Z(n_156176627));
	notech_ao4 i_127264914(.A(n_30916), .B(n_139176457), .C(n_83739557), .D(n_117476240
		), .Z(n_156376629));
	notech_ao4 i_127164915(.A(n_30896), .B(n_116576231), .C(n_30914), .D(n_139276458
		), .Z(n_156476630));
	notech_ao4 i_126964917(.A(n_330460932), .B(n_33417), .C(n_55793), .D(n_33416
		), .Z(n_156676632));
	notech_ao4 i_126864918(.A(n_57277), .B(n_33103), .C(n_334360971), .D(n_57276
		), .Z(n_156776633));
	notech_and4 i_127464912(.A(n_156776633), .B(n_156676632), .C(n_156476630
		), .D(n_156376629), .Z(n_156976635));
	notech_ao4 i_126564921(.A(n_59005), .B(n_334778353), .C(n_58229), .D(n_334878354
		), .Z(n_157076636));
	notech_ao4 i_126464922(.A(n_334060968), .B(n_328760915), .C(n_30891), .D
		(n_57439), .Z(n_157176637));
	notech_ao4 i_126264924(.A(n_61097), .B(n_30811), .C(n_58040), .D(n_31473
		), .Z(n_157376639));
	notech_and3 i_126364923(.A(n_169484150), .B(n_157376639), .C(n_142483880
		), .Z(n_157476640));
	notech_ao4 i_125964927(.A(\nbus_11290[0] ), .B(n_117376239), .C(nbus_11273
		[0]), .D(n_30277), .Z(n_157676642));
	notech_ao4 i_125764929(.A(n_55793), .B(n_33415), .C(n_327660904), .D(n_139276458
		), .Z(n_157876644));
	notech_and4 i_126164925(.A(n_157876644), .B(n_157676642), .C(n_120476270
		), .D(n_120776273), .Z(n_158076646));
	notech_ao4 i_125464932(.A(n_57277), .B(n_33169), .C(n_101142452), .D(n_57276
		), .Z(n_158176647));
	notech_ao4 i_125264934(.A(n_61097), .B(n_30810), .C(n_58040), .D(n_31472
		), .Z(n_158376649));
	notech_and3 i_125364933(.A(n_116976235), .B(n_169576761), .C(n_158376649
		), .Z(n_158476650));
	notech_ao4 i_105165117(.A(\nbus_11290[14] ), .B(n_117176237), .C(nbus_11273
		[14]), .D(n_117076236), .Z(n_158676652));
	notech_ao4 i_105065118(.A(n_323978248), .B(n_33215), .C(n_57072), .D(n_377064301
		), .Z(n_158876654));
	notech_ao4 i_104865120(.A(n_377164302), .B(n_333778343), .C(n_97342414),
		 .D(n_323778246), .Z(n_159076656));
	notech_and3 i_104965119(.A(n_186576923), .B(n_159076656), .C(n_118976255
		), .Z(n_159276658));
	notech_and2 i_15463205(.A(n_56615), .B(n_178076840), .Z(n_159576661));
	notech_and2 i_15563204(.A(n_56640), .B(n_178176841), .Z(n_159676662));
	notech_mux2 i_15063209(.S(n_32263), .A(n_160176667), .B(n_159976665), .Z
		(n_159776663));
	notech_ao4 i_11363244(.A(n_60170), .B(n_59005), .C(n_30920), .D(n_26063)
		, .Z(n_159976665));
	notech_ao4 i_11263245(.A(n_60170), .B(n_58229), .C(n_30919), .D(n_26063)
		, .Z(n_160176667));
	notech_nor2 i_14563214(.A(n_171976781), .B(n_329860926), .Z(n_160476670)
		);
	notech_and3 i_14663213(.A(n_330060928), .B(n_167376739), .C(n_329760925)
		, .Z(n_160576671));
	notech_mux2 i_14163218(.S(n_32252), .A(n_161076676), .B(n_160876674), .Z
		(n_160676672));
	notech_ao4 i_10563252(.A(n_60170), .B(n_59005), .C(n_30920), .D(n_29214)
		, .Z(n_160876674));
	notech_ao4 i_10463253(.A(n_60175), .B(n_58229), .C(n_30919), .D(n_29214)
		, .Z(n_161076676));
	notech_or4 i_25063110(.A(n_61870), .B(n_61679), .C(n_19680), .D(n_31508)
		, .Z(n_161776683));
	notech_or2 i_24763113(.A(n_381164342), .B(n_31472), .Z(n_162076686));
	notech_or4 i_46362914(.A(n_63698), .B(n_57438), .C(n_63760), .D(n_58229)
		, .Z(n_162576691));
	notech_nao3 i_46162915(.A(n_63774), .B(opc_10[1]), .C(n_150969547), .Z(n_162876694
		));
	notech_or2 i_45862918(.A(n_57027), .B(n_33103), .Z(n_163176697));
	notech_nao3 i_55862824(.A(opc_10[30]), .B(n_63760), .C(n_298922014), .Z(n_163876704
		));
	notech_or2 i_55362829(.A(n_57217), .B(\nbus_11290[30] ), .Z(n_164376709)
		);
	notech_nand2 i_59362790(.A(sav_esp[7]), .B(n_61870), .Z(n_165176717));
	notech_or2 i_58862795(.A(n_332460952), .B(n_100242443), .Z(n_165676722)
		);
	notech_nao3 i_58362800(.A(n_63774), .B(opc_10[7]), .C(n_26271), .Z(n_166176727
		));
	notech_or2 i_64262741(.A(n_57274), .B(n_33215), .Z(n_166676732));
	notech_or2 i_63962744(.A(n_58025), .B(n_31487), .Z(n_166976735));
	notech_nand2 i_63662747(.A(sav_esi[14]), .B(n_61866), .Z(n_167276738));
	notech_nao3 i_64662737(.A(n_32243), .B(n_30276), .C(n_163196017), .Z(n_167376739
		));
	notech_or4 i_72162662(.A(n_335478360), .B(n_61935), .C(n_31612), .D(n_30319
		), .Z(n_167976745));
	notech_or2 i_71862665(.A(n_192676984), .B(n_33103), .Z(n_168276748));
	notech_ao3 i_74862635(.A(opc_10[30]), .B(n_63760), .C(n_315725234), .Z(n_168776753
		));
	notech_or2 i_74362640(.A(n_57200), .B(\nbus_11290[30] ), .Z(n_169476760)
		);
	notech_ao4 i_31294(.A(n_331360941), .B(\nbus_11290[0] ), .C(n_28240), .D
		(nbus_11273[0]), .Z(n_169576761));
	notech_or2 i_12763232(.A(n_57666), .B(n_29214), .Z(n_169676762));
	notech_ao4 i_150761906(.A(n_324778256), .B(n_33194), .C(n_5758), .D(n_324878257
		), .Z(n_169776763));
	notech_ao4 i_150661907(.A(n_5750), .B(n_325325323), .C(\nbus_11283[30] )
		, .D(n_57201), .Z(n_169976765));
	notech_nand3 i_150961904(.A(n_169776763), .B(n_169976765), .C(n_169476760
		), .Z(n_170076766));
	notech_ao4 i_150461909(.A(n_324978258), .B(nbus_11271[30]), .C(n_58088),
		 .D(n_31506), .Z(n_170176767));
	notech_ao4 i_148861925(.A(n_30896), .B(n_169676762), .C(n_323578244), .D
		(n_160676672), .Z(n_170476770));
	notech_ao4 i_148761926(.A(n_323078239), .B(n_58229), .C(n_30280), .D(n_57616
		), .Z(n_170576771));
	notech_ao4 i_148561928(.A(n_334360971), .B(n_323278241), .C(n_323178240)
		, .D(n_59005), .Z(n_170776773));
	notech_and4 i_149061923(.A(n_170776773), .B(n_170576771), .C(n_170476770
		), .D(n_168276748), .Z(n_170976775));
	notech_ao4 i_148261931(.A(n_58044), .B(n_31473), .C(n_30914), .D(n_200477060
		), .Z(n_171076776));
	notech_ao4 i_148061933(.A(n_279977810), .B(nbus_11271[1]), .C(n_30891), 
		.D(n_57666), .Z(n_171276778));
	notech_and4 i_148461929(.A(n_30274), .B(n_171276778), .C(n_167976745), .D
		(n_171076776), .Z(n_171476780));
	notech_ao4 i_138562027(.A(n_32697), .B(n_31363), .C(n_30275), .D(n_30276
		), .Z(n_171976781));
	notech_ao4 i_138162031(.A(\nbus_11290[14] ), .B(n_160576671), .C(nbus_11273
		[14]), .D(n_160476670), .Z(n_172376783));
	notech_ao4 i_137962033(.A(n_55793), .B(n_33440), .C(n_330460932), .D(n_33439
		), .Z(n_172576785));
	notech_and4 i_138362029(.A(n_172576785), .B(n_172376783), .C(n_166976735
		), .D(n_167276738), .Z(n_172776787));
	notech_ao4 i_137662036(.A(n_97342414), .B(n_57275), .C(n_385364384), .D(n_328860916
		), .Z(n_172876788));
	notech_ao4 i_137362038(.A(n_377264303), .B(n_334178347), .C(n_377164302)
		, .D(n_334078346), .Z(n_173076790));
	notech_and3 i_137462037(.A(n_169684152), .B(n_160684062), .C(n_173076790
		), .Z(n_173176791));
	notech_ao4 i_134162070(.A(n_26268), .B(n_324560873), .C(n_26278), .D(n_324160869
		), .Z(n_173376793));
	notech_ao4 i_134062071(.A(n_26277), .B(n_324360871), .C(n_26272), .D(n_324760875
		), .Z(n_173576795));
	notech_and3 i_134362068(.A(n_173376793), .B(n_173576795), .C(n_166176727
		), .Z(n_173676796));
	notech_ao4 i_133762074(.A(n_26276), .B(n_324460872), .C(n_324260870), .D
		(n_26275), .Z(n_173776797));
	notech_ao4 i_133662075(.A(n_332160949), .B(n_324060868), .C(n_332260950)
		, .D(n_33165), .Z(n_173976799));
	notech_and4 i_134462067(.A(n_173776797), .B(n_173976799), .C(n_165676722
		), .D(n_173676796), .Z(n_174176801));
	notech_ao4 i_133262079(.A(n_331160939), .B(\nbus_11290[7] ), .C(n_331460942
		), .D(n_31480), .Z(n_174276802));
	notech_ao4 i_133162080(.A(n_125926586), .B(n_33438), .C(n_26603), .D(n_336060988
		), .Z(n_174476804));
	notech_and3 i_133462077(.A(n_174276802), .B(n_174476804), .C(n_165176717
		), .Z(n_174576805));
	notech_ao4 i_132962082(.A(n_26585), .B(n_30981), .C(n_126126588), .D(n_32066
		), .Z(n_174676806));
	notech_ao4 i_132862083(.A(n_28240), .B(nbus_11273[7]), .C(n_26600), .D(n_31515
		), .Z(n_174776807));
	notech_ao4 i_131362098(.A(n_324178250), .B(n_33194), .C(n_5758), .D(n_324278251
		), .Z(n_175076810));
	notech_ao4 i_131262099(.A(n_5750), .B(n_301522040), .C(\nbus_11283[30] )
		, .D(n_57213), .Z(n_175276812));
	notech_ao4 i_130962102(.A(nbus_11271[30]), .B(n_301822043), .C(n_58083),
		 .D(n_31506), .Z(n_175476814));
	notech_and4 i_131162100(.A(n_5774), .B(n_175476814), .C(n_30502), .D(n_163876704
		), .Z(n_175776817));
	notech_ao4 i_122362180(.A(n_30280), .B(n_30473), .C(n_324078249), .D(n_159776663
		), .Z(n_175876818));
	notech_ao4 i_122262181(.A(n_58229), .B(n_322878237), .C(n_143769475), .D
		(n_30896), .Z(n_175976819));
	notech_ao4 i_122062183(.A(n_57036), .B(n_334360971), .C(n_59005), .D(n_322978238
		), .Z(n_176176821));
	notech_and4 i_122662178(.A(n_176176821), .B(n_175976819), .C(n_175876818
		), .D(n_163176697), .Z(n_176376823));
	notech_ao4 i_121762186(.A(n_5783), .B(n_31473), .C(n_151069548), .D(n_30914
		), .Z(n_176476824));
	notech_and3 i_121662187(.A(n_30274), .B(n_5774), .C(n_162576691), .Z(n_176776827
		));
	notech_ao4 i_103662361(.A(\nbus_11290[0] ), .B(n_159676662), .C(nbus_11273
		[0]), .D(n_159576661), .Z(n_176976829));
	notech_ao4 i_103562362(.A(n_24424), .B(n_327660904), .C(n_24421), .D(n_327760905
		), .Z(n_177076830));
	notech_ao4 i_103362364(.A(n_381064341), .B(n_33169), .C(n_380964340), .D
		(n_101142452), .Z(n_177276832));
	notech_and4 i_103862359(.A(n_177276832), .B(n_177076830), .C(n_176976829
		), .D(n_162076686), .Z(n_177476834));
	notech_ao4 i_102962367(.A(n_336760995), .B(n_24717), .C(n_61097), .D(n_30760
		), .Z(n_177576835));
	notech_ao4 i_102762369(.A(n_24528), .B(n_33437), .C(n_24527), .D(n_33436
		), .Z(n_177776837));
	notech_and4 i_103262365(.A(n_177776837), .B(n_169576761), .C(n_177576835
		), .D(n_161776683), .Z(n_177976839));
	notech_or2 i_108760723(.A(n_383164362), .B(n_186876926), .Z(n_178076840)
		);
	notech_or4 i_108860722(.A(n_32275), .B(n_318160809), .C(n_256763514), .D
		(n_186876926), .Z(n_178176841));
	notech_and2 i_25260703(.A(n_116742608), .B(n_180276862), .Z(n_178276842)
		);
	notech_or2 i_133460654(.A(n_57432), .B(n_30315), .Z(n_178376843));
	notech_or4 i_179260641(.A(n_2580), .B(n_178376843), .C(n_32159), .D(n_32161
		), .Z(n_178476844));
	notech_nao3 i_179460640(.A(n_58279), .B(n_57529), .C(n_57432), .Z(n_178576845
		));
	notech_or2 i_179760639(.A(n_57432), .B(n_32254), .Z(n_178676846));
	notech_or4 i_179860638(.A(n_2580), .B(n_57432), .C(n_32159), .D(n_32161)
		, .Z(n_178776847));
	notech_or4 i_184560637(.A(n_316160789), .B(n_61725), .C(n_61679), .D(n_19680
		), .Z(n_178876848));
	notech_and3 i_5160589(.A(n_57217), .B(n_323778246), .C(n_323678245), .Z(n_178976849
		));
	notech_ao3 i_5260588(.A(n_57213), .B(n_323978248), .C(n_323878247), .Z(n_179076850
		));
	notech_and2 i_4660594(.A(n_197877035), .B(n_192476982), .Z(n_179176851)
		);
	notech_mux2 i_4760593(.S(n_32254), .A(n_179776857), .B(n_179576855), .Z(n_179276852
		));
	notech_and2 i_4860592(.A(n_193076988), .B(n_30322), .Z(n_179376853));
	notech_ao4 i_4960591(.A(n_60175), .B(\nbus_11290[1] ), .C(n_30920), .D(n_30315
		), .Z(n_179576855));
	notech_ao4 i_5060590(.A(n_60175), .B(nbus_11273[1]), .C(n_30919), .D(n_30315
		), .Z(n_179776857));
	notech_ao3 i_71059995(.A(n_328560913), .B(n_186876926), .C(n_258063525),
		 .Z(n_180076860));
	notech_or4 i_76959936(.A(n_61889), .B(n_61725), .C(n_30306), .D(n_57657)
		, .Z(n_180176861));
	notech_or4 i_78959916(.A(n_61823), .B(n_30309), .C(n_30698), .D(n_32210)
		, .Z(n_180276862));
	notech_or2 i_44660231(.A(n_30473), .B(n_327560903), .Z(n_180976869));
	notech_nao3 i_44060236(.A(n_63774), .B(opc[0]), .C(n_151069548), .Z(n_181476874
		));
	notech_nand3 i_53560167(.A(n_30524), .B(n_61621), .C(n_30336), .Z(n_182376883
		));
	notech_or2 i_62760076(.A(n_31071), .B(n_140076466), .Z(n_185476912));
	notech_nand2 i_70759998(.A(n_61621), .B(read_data[4]), .Z(n_186376921)
		);
	notech_and2 i_33502(.A(n_5774), .B(n_377364304), .Z(n_186576923));
	notech_ao3 i_112660660(.A(n_328160909), .B(n_24733), .C(n_2579), .Z(n_186876926
		));
	notech_nao3 i_47860687(.A(n_32323), .B(n_32310), .C(n_334760975), .Z(n_187176929
		));
	notech_ao4 i_154259217(.A(n_30376), .B(n_33104), .C(n_30378), .D(nbus_11273
		[4]), .Z(n_187276930));
	notech_ao4 i_154159218(.A(n_30379), .B(n_334660974), .C(n_30373), .D(\nbus_11290[4] 
		), .Z(n_187476932));
	notech_and3 i_49260677(.A(n_187276930), .B(n_187476932), .C(n_186376921)
		, .Z(n_187576933));
	notech_ao4 i_146359284(.A(n_334660974), .B(n_323278241), .C(n_57616), .D
		(n_187176929), .Z(n_187676934));
	notech_ao4 i_146259285(.A(n_58044), .B(n_31477), .C(n_192676984), .D(n_33104
		), .Z(n_187776935));
	notech_ao4 i_146059287(.A(n_31048), .B(n_169676762), .C(n_31047), .D(n_57666
		), .Z(n_187976937));
	notech_and4 i_146659282(.A(n_187976937), .B(n_187776935), .C(n_187676934
		), .D(n_185476912), .Z(n_188176939));
	notech_ao4 i_145759290(.A(n_31072), .B(n_140176467), .C(n_31074), .D(n_139876464
		), .Z(n_188276940));
	notech_ao4 i_145659291(.A(n_31068), .B(n_200377059), .C(n_31067), .D(n_200477060
		), .Z(n_188376941));
	notech_ao4 i_145459293(.A(n_279977810), .B(nbus_11271[4]), .C(n_31075), 
		.D(n_139976465), .Z(n_188576943));
	notech_and4 i_145959288(.A(n_187576933), .B(n_188576943), .C(n_188376941
		), .D(n_188276940), .Z(n_188776945));
	notech_ao4 i_139859347(.A(n_31071), .B(n_178676846), .C(n_31072), .D(n_178776847
		), .Z(n_188876946));
	notech_ao4 i_139759348(.A(n_31074), .B(n_178476844), .C(n_31075), .D(n_178576845
		), .Z(n_188976947));
	notech_ao4 i_139559350(.A(n_57157), .B(n_187176929), .C(n_31048), .D(n_178376843
		), .Z(n_189176949));
	notech_ao4 i_139459351(.A(n_197877035), .B(\nbus_11290[4] ), .C(n_56608)
		, .D(nbus_11273[4]), .Z(n_189276950));
	notech_and4 i_140059345(.A(n_189276950), .B(n_189176949), .C(n_188976947
		), .D(n_188876946), .Z(n_189476952));
	notech_ao4 i_139159354(.A(n_334660974), .B(n_57289), .C(n_245877510), .D
		(n_31512), .Z(n_189576953));
	notech_ao4 i_139059355(.A(n_58019), .B(n_31477), .C(n_204977105), .D(n_33104
		), .Z(n_189676954));
	notech_ao4 i_138859357(.A(n_31067), .B(n_200977065), .C(n_31047), .D(n_57432
		), .Z(n_189876956));
	notech_ao4 i_138759358(.A(n_193576993), .B(n_30942), .C(n_200877064), .D
		(n_31068), .Z(n_189976957));
	notech_and4 i_139359352(.A(n_189976957), .B(n_189876956), .C(n_189676954
		), .D(n_189576953), .Z(n_190176959));
	notech_ao4 i_136159379(.A(n_192776985), .B(n_179276852), .C(n_179176851)
		, .D(\nbus_11290[1] ), .Z(n_190276960));
	notech_ao4 i_136059380(.A(n_178876848), .B(n_31509), .C(nbus_11273[1]), 
		.D(n_179376853), .Z(n_190376961));
	notech_ao4 i_135859382(.A(n_57010), .B(n_33103), .C(n_30896), .D(n_178376843
		), .Z(n_190576963));
	notech_and4 i_136359377(.A(n_190576963), .B(n_190376961), .C(n_190276960
		), .D(n_182376883), .Z(n_190776965));
	notech_ao4 i_135559385(.A(n_30280), .B(n_57158), .C(n_58019), .D(n_31473
		), .Z(n_190876966));
	notech_ao4 i_135459386(.A(n_334360971), .B(n_57289), .C(n_30891), .D(n_57432
		), .Z(n_190976967));
	notech_ao4 i_135259388(.A(n_30914), .B(n_200977065), .C(n_30916), .D(n_200877064
		), .Z(n_191176969));
	notech_and4 i_135759383(.A(n_56896), .B(n_191176969), .C(n_190976967), .D
		(n_190876966), .Z(n_191376971));
	notech_ao4 i_118259541(.A(nbus_11273[0]), .B(n_179076850), .C(\nbus_11290[0] 
		), .D(n_178976849), .Z(n_191676974));
	notech_ao4 i_117959542(.A(n_57027), .B(n_33169), .C(n_150969547), .D(n_327760905
		), .Z(n_191876976));
	notech_ao4 i_117659545(.A(n_5783), .B(n_31472), .C(n_57036), .D(n_101142452
		), .Z(n_192076978));
	notech_and4 i_117859543(.A(n_5774), .B(n_327860906), .C(n_180976869), .D
		(n_192076978), .Z(n_192376981));
	notech_nao3 i_119158179(.A(n_201477070), .B(n_32254), .C(n_193276990), .Z
		(n_192476982));
	notech_and2 i_25358156(.A(n_116742608), .B(n_195877016), .Z(n_192576983)
		);
	notech_or2 i_88958154(.A(n_376064291), .B(n_335478360), .Z(n_192676984)
		);
	notech_ao4 i_30558151(.A(n_57679), .B(n_32314), .C(n_30719), .D(n_32223)
		, .Z(n_192776985));
	notech_ao4 i_46358138(.A(n_30317), .B(n_30420), .C(n_32317), .D(n_30528)
		, .Z(n_192876986));
	notech_nao3 i_119058182(.A(n_57529), .B(n_201477070), .C(n_193276990), .Z
		(n_193076988));
	notech_or4 i_162958117(.A(n_61917), .B(n_61901), .C(n_61889), .D(eval_flag
		), .Z(n_193176989));
	notech_ao4 i_125158122(.A(n_63774), .B(n_61958), .C(n_61056), .D(n_30315
		), .Z(n_193276990));
	notech_and4 i_3658085(.A(n_56720), .B(n_279677807), .C(n_56608), .D(n_198077037
		), .Z(n_193376991));
	notech_and4 i_3758084(.A(n_197877035), .B(n_303178041), .C(n_279877809),
		 .D(n_197977036), .Z(n_193476992));
	notech_and2 i_53758160(.A(n_57426), .B(n_56896), .Z(n_193576993));
	notech_and2 i_30258141(.A(n_116742608), .B(n_195677014), .Z(n_193676994)
		);
	notech_ao4 i_3458087(.A(n_32697), .B(n_30732), .C(n_201377069), .D(n_30300
		), .Z(n_193776995));
	notech_and2 i_3558086(.A(n_323378242), .B(n_323178240), .Z(n_193876996)
		);
	notech_ao4 i_2058101(.A(n_61056), .B(n_3452), .C(n_57194), .D(n_30936), 
		.Z(n_194176999));
	notech_nao3 i_75957404(.A(n_57529), .B(n_30318), .C(n_195177009), .Z(n_194377001
		));
	notech_and2 i_181058159(.A(n_58058), .B(n_342578429), .Z(n_194577003));
	notech_and2 i_121558123(.A(n_196377020), .B(n_58058), .Z(n_194777005));
	notech_or4 i_76757396(.A(n_2382), .B(n_2580), .C(n_193276990), .D(n_195177009
		), .Z(n_195077008));
	notech_ao4 i_30458140(.A(n_57566), .B(n_57657), .C(n_30723), .D(n_32223)
		, .Z(n_195177009));
	notech_or4 i_76857395(.A(n_1850), .B(n_57679), .C(n_61621), .D(eval_flag
		), .Z(n_195277010));
	notech_or4 i_77157392(.A(n_32574), .B(n_60170), .C(n_32394), .D(n_61621)
		, .Z(n_195577013));
	notech_or4 i_77257391(.A(n_61823), .B(n_30309), .C(n_30698), .D(n_32223)
		, .Z(n_195677014));
	notech_or4 i_77557388(.A(n_61823), .B(n_30309), .C(n_30698), .D(n_32227)
		, .Z(n_195877016));
	notech_nao3 i_77657387(.A(instrc[112]), .B(n_115942600), .C(n_2821), .Z(n_196077017
		));
	notech_nand2 i_77757386(.A(n_115942600), .B(n_32227), .Z(n_196177018));
	notech_nao3 i_77857385(.A(instrc[112]), .B(n_115442595), .C(n_2821), .Z(n_196277019
		));
	notech_or4 i_77957384(.A(n_32394), .B(n_60194), .C(n_193176989), .D(n_32574
		), .Z(n_196377020));
	notech_or2 i_69257471(.A(n_204977105), .B(n_33169), .Z(n_197277029));
	notech_or2 i_68757476(.A(n_57158), .B(n_327560903), .Z(n_197777034));
	notech_or2 i_161758157(.A(n_30373), .B(eval_flag), .Z(n_197877035));
	notech_or4 i_69657467(.A(n_2382), .B(n_2580), .C(n_193276990), .D(n_193676994
		), .Z(n_197977036));
	notech_or2 i_69557468(.A(n_56766), .B(n_193676994), .Z(n_198077037));
	notech_or2 i_71057453(.A(n_58053), .B(n_31482), .Z(n_198377040));
	notech_or2 i_70757456(.A(n_57252), .B(n_33168), .Z(n_198677043));
	notech_nand2 i_70457459(.A(ie), .B(n_30595), .Z(n_198977046));
	notech_or4 i_70157462(.A(n_192776985), .B(n_61935), .C(n_31620), .D(n_58279
		), .Z(n_199277049));
	notech_or2 i_73757426(.A(n_279977810), .B(nbus_11271[0]), .Z(n_199377050
		));
	notech_or2 i_73657427(.A(n_58044), .B(n_31472), .Z(n_199677053));
	notech_or4 i_73157432(.A(instrc[113]), .B(instrc[114]), .C(n_339561023),
		 .D(n_327560903), .Z(n_200277058));
	notech_nao3 i_30413(.A(n_33173), .B(n_286063762), .C(n_335478360), .Z(n_200377059
		));
	notech_or2 i_30409(.A(n_57666), .B(n_30319), .Z(n_200477060));
	notech_or2 i_31769(.A(n_192776985), .B(n_58279), .Z(n_200577061));
	notech_or2 i_31762(.A(n_57388), .B(n_58279), .Z(n_200677062));
	notech_or2 i_31765(.A(n_57388), .B(n_30315), .Z(n_200777063));
	notech_or2 i_31900(.A(n_195177009), .B(n_58279), .Z(n_200877064));
	notech_or2 i_31898(.A(n_57432), .B(n_58279), .Z(n_200977065));
	notech_or2 i_11431(.A(n_30496), .B(eval_flag), .Z(n_201077066));
	notech_nand3 i_81558153(.A(n_116742608), .B(n_195877016), .C(n_280977820
		), .Z(n_201377069));
	notech_nand3 i_106158124(.A(n_116742608), .B(n_195677014), .C(n_280377814
		), .Z(n_201477070));
	notech_ao4 i_142856766(.A(n_32254), .B(n_193276990), .C(n_60194), .D(n_30315
		), .Z(n_201777073));
	notech_ao4 i_134256847(.A(\nbus_11290[0] ), .B(n_193876996), .C(nbus_11273
		[0]), .D(n_30288), .Z(n_201977075));
	notech_ao4 i_134156848(.A(n_327760905), .B(n_200377059), .C(n_192676984)
		, .D(n_33169), .Z(n_202177077));
	notech_ao4 i_133856851(.A(n_101142452), .B(n_323278241), .C(n_200477060)
		, .D(n_327660904), .Z(n_202377079));
	notech_and4 i_134056849(.A(n_327860906), .B(n_202377079), .C(n_199377050
		), .D(n_199677053), .Z(n_202677082));
	notech_ao4 i_128756902(.A(n_57158), .B(n_326960897), .C(n_245877510), .D
		(n_31517), .Z(n_202777083));
	notech_ao4 i_128556904(.A(n_200777063), .B(n_327360901), .C(n_327160899)
		, .D(n_200677062), .Z(n_202977085));
	notech_and4 i_128956900(.A(n_202977085), .B(n_202777083), .C(n_198977046
		), .D(n_199277049), .Z(n_203177087));
	notech_ao4 i_128256907(.A(n_57133), .B(\nbus_11290[9] ), .C(n_57110), .D
		(nbus_11273[9]), .Z(n_203277088));
	notech_ao4 i_128056909(.A(n_327060898), .B(n_57388), .C(n_99942440), .D(n_57317
		), .Z(n_203477090));
	notech_and4 i_128456905(.A(n_203477090), .B(n_203277088), .C(n_198377040
		), .D(n_198677043), .Z(n_203677092));
	notech_ao4 i_126856921(.A(n_193476992), .B(\nbus_11290[0] ), .C(nbus_11273
		[0]), .D(n_193376991), .Z(n_204177097));
	notech_ao4 i_126756922(.A(n_193576993), .B(n_30939), .C(n_31508), .D(n_245877510
		), .Z(n_204377099));
	notech_and3 i_127056919(.A(n_204177097), .B(n_204377099), .C(n_197777034
		), .Z(n_204477100));
	notech_ao4 i_126456925(.A(n_327660904), .B(n_200977065), .C(n_327760905)
		, .D(n_200877064), .Z(n_204577101));
	notech_ao4 i_126356926(.A(n_58019), .B(n_31472), .C(n_101142452), .D(n_57289
		), .Z(n_204777103));
	notech_ao4 i_122758184(.A(n_56766), .B(n_195177009), .C(n_57657), .D(n_194777005
		), .Z(n_204977105));
	notech_or2 i_19755751(.A(n_57369), .B(\nbus_11283[28] ), .Z(n_205477110)
		);
	notech_or2 i_19455754(.A(n_57326), .B(n_33196), .Z(n_205777113));
	notech_nand2 i_19155757(.A(sav_ecx[28]), .B(n_61866), .Z(n_206077116));
	notech_or2 i_25555694(.A(n_301822043), .B(nbus_11271[26]), .Z(n_206477119
		));
	notech_nao3 i_24955699(.A(n_57392), .B(opd[26]), .C(n_30473), .Z(n_206977124
		));
	notech_nor2 i_26555686(.A(n_301822043), .B(nbus_11271[27]), .Z(n_207077125
		));
	notech_nao3 i_25855691(.A(n_57392), .B(opd[27]), .C(n_30473), .Z(n_207777132
		));
	notech_or2 i_27555678(.A(n_301822043), .B(nbus_11271[28]), .Z(n_208077135
		));
	notech_nand3 i_26855683(.A(n_57392), .B(n_32210), .C(opd[28]), .Z(n_208677140
		));
	notech_or2 i_28555670(.A(n_301822043), .B(nbus_11271[29]), .Z(n_208977143
		));
	notech_nand3 i_27855675(.A(n_57395), .B(n_32210), .C(opd[29]), .Z(n_209477148
		));
	notech_nao3 i_38155574(.A(n_164196010), .B(n_2691), .C(n_163296016), .Z(n_209777151
		));
	notech_or2 i_37855577(.A(n_124626573), .B(\nbus_11283[26] ), .Z(n_210077154
		));
	notech_or2 i_37555580(.A(n_124726574), .B(n_33198), .Z(n_210377157));
	notech_nand2 i_37255583(.A(sav_esi[26]), .B(n_61870), .Z(n_210677160));
	notech_nao3 i_39555562(.A(n_164196010), .B(n_2693), .C(n_163296016), .Z(n_210977163
		));
	notech_or2 i_39255565(.A(n_124626573), .B(\nbus_11283[27] ), .Z(n_211277166
		));
	notech_or2 i_38755568(.A(n_124726574), .B(n_33195), .Z(n_211577169));
	notech_nand2 i_38455571(.A(sav_esi[27]), .B(n_61866), .Z(n_211877172));
	notech_nao3 i_40755550(.A(n_164196010), .B(n_2695), .C(n_163296016), .Z(n_212177175
		));
	notech_or2 i_40455553(.A(n_124626573), .B(\nbus_11283[28] ), .Z(n_212477178
		));
	notech_or2 i_40155556(.A(n_124726574), .B(n_33196), .Z(n_212777181));
	notech_nand2 i_39855559(.A(sav_esi[28]), .B(n_61871), .Z(n_213077184));
	notech_nao3 i_41955538(.A(n_164196010), .B(n_2697), .C(n_163296016), .Z(n_213377187
		));
	notech_or2 i_41655541(.A(n_124626573), .B(\nbus_11283[29] ), .Z(n_213677190
		));
	notech_or2 i_41355544(.A(n_124726574), .B(n_33197), .Z(n_213977193));
	notech_nand2 i_41055547(.A(sav_esi[29]), .B(n_61873), .Z(n_214277196));
	notech_ao3 i_44155518(.A(n_57395), .B(opd[26]), .C(n_57158), .Z(n_215377205
		));
	notech_ao3 i_45055509(.A(n_57392), .B(opd[27]), .C(n_57158), .Z(n_216277214
		));
	notech_ao3 i_45955500(.A(n_57392), .B(opd[28]), .C(n_57158), .Z(n_217177223
		));
	notech_nao3 i_46855491(.A(n_57392), .B(opd[29]), .C(n_57158), .Z(n_218077232
		));
	notech_nor2 i_62755339(.A(n_324978258), .B(nbus_11271[26]), .Z(n_218177233
		));
	notech_nao3 i_62255344(.A(n_57392), .B(opd[26]), .C(n_57616), .Z(n_218877240
		));
	notech_nor2 i_63555331(.A(n_324978258), .B(nbus_11271[27]), .Z(n_218977241
		));
	notech_nao3 i_63055336(.A(n_57386), .B(opd[27]), .C(n_57616), .Z(n_219677248
		));
	notech_nor2 i_64355323(.A(n_324978258), .B(nbus_11271[28]), .Z(n_219777249
		));
	notech_nand3 i_63855328(.A(n_57386), .B(n_32227), .C(opd[28]), .Z(n_220477256
		));
	notech_or2 i_65155315(.A(n_324978258), .B(nbus_11271[29]), .Z(n_220577257
		));
	notech_nand3 i_64655320(.A(n_57386), .B(n_32227), .C(opd[29]), .Z(n_221277264
		));
	notech_or2 i_84655126(.A(n_30693), .B(\nbus_11290[29] ), .Z(n_221677268)
		);
	notech_ao4 i_172254274(.A(n_30689), .B(n_4428), .C(n_30697), .D(n_33197)
		, .Z(n_221777269));
	notech_ao4 i_172154275(.A(n_31537), .B(n_61679), .C(n_30695), .D(\nbus_11283[29] 
		), .Z(n_221977271));
	notech_and3 i_52155918(.A(n_221777269), .B(n_221977271), .C(n_221677268)
		, .Z(n_222077272));
	notech_ao4 i_147054520(.A(n_4387), .B(n_325325323), .C(n_94229643), .D(n_315725234
		), .Z(n_222177273));
	notech_ao4 i_146954521(.A(n_4428), .B(n_324878257), .C(n_324778256), .D(n_33197
		), .Z(n_222377275));
	notech_and3 i_147254518(.A(n_222177273), .B(n_222377275), .C(n_221277264
		), .Z(n_222477276));
	notech_ao4 i_146754523(.A(n_57201), .B(\nbus_11283[29] ), .C(n_57200), .D
		(\nbus_11290[29] ), .Z(n_222577277));
	notech_ao4 i_146354527(.A(n_440082450), .B(n_325325323), .C(n_7636), .D(n_315725234
		), .Z(n_222877280));
	notech_ao4 i_146254528(.A(n_4427), .B(n_324878257), .C(n_324778256), .D(n_33196
		), .Z(n_223077282));
	notech_nand3 i_146554525(.A(n_222877280), .B(n_223077282), .C(n_220477256
		), .Z(n_223177283));
	notech_ao4 i_146054530(.A(n_57201), .B(\nbus_11283[28] ), .C(n_57200), .D
		(\nbus_11290[28] ), .Z(n_223277284));
	notech_ao4 i_145654534(.A(n_284131522), .B(n_325325323), .C(n_172669762)
		, .D(n_315725234), .Z(n_223577287));
	notech_ao4 i_145554535(.A(n_5711), .B(n_324878257), .C(n_324778256), .D(n_33195
		), .Z(n_223777289));
	notech_nand3 i_145854532(.A(n_223577287), .B(n_223777289), .C(n_219677248
		), .Z(n_223877290));
	notech_ao4 i_145354537(.A(n_57201), .B(\nbus_11283[27] ), .C(n_57200), .D
		(\nbus_11290[27] ), .Z(n_223977291));
	notech_ao4 i_144954541(.A(n_284231523), .B(n_325325323), .C(n_175169787)
		, .D(n_315725234), .Z(n_224277294));
	notech_ao4 i_144854542(.A(n_5720), .B(n_324878257), .C(n_33198), .D(n_324778256
		), .Z(n_224477296));
	notech_nand3 i_145154539(.A(n_224277294), .B(n_224477296), .C(n_218877240
		), .Z(n_224577297));
	notech_ao4 i_144654544(.A(n_57201), .B(\nbus_11283[26] ), .C(n_57200), .D
		(\nbus_11290[26] ), .Z(n_224677298));
	notech_ao4 i_131554675(.A(n_4387), .B(n_302878038), .C(n_94229643), .D(n_303078040
		), .Z(n_224977301));
	notech_ao4 i_131454676(.A(n_324378252), .B(n_33197), .C(n_245877510), .D
		(n_31537), .Z(n_225177303));
	notech_and3 i_131754673(.A(n_224977301), .B(n_225177303), .C(n_218077232
		), .Z(n_225277304));
	notech_ao4 i_131254678(.A(n_324578254), .B(\nbus_11290[29] ), .C(n_4428)
		, .D(n_324478253), .Z(n_225377305));
	notech_ao4 i_131154679(.A(n_302978039), .B(nbus_11271[29]), .C(n_324678255
		), .D(\nbus_11283[29] ), .Z(n_225477306));
	notech_ao4 i_130854682(.A(n_440082450), .B(n_302878038), .C(n_7636), .D(n_303078040
		), .Z(n_225677308));
	notech_ao4 i_130754683(.A(n_324378252), .B(n_33196), .C(n_245877510), .D
		(n_31536), .Z(n_225877310));
	notech_ao3 i_131054680(.A(n_225677308), .B(n_225877310), .C(n_217177223)
		, .Z(n_225977311));
	notech_ao4 i_130554685(.A(n_324578254), .B(\nbus_11290[28] ), .C(n_4427)
		, .D(n_324478253), .Z(n_226077312));
	notech_ao4 i_130454686(.A(n_302978039), .B(nbus_11271[28]), .C(n_324678255
		), .D(\nbus_11283[28] ), .Z(n_226177313));
	notech_ao4 i_130154689(.A(n_284131522), .B(n_302878038), .C(n_172669762)
		, .D(n_303078040), .Z(n_226377315));
	notech_ao4 i_130054690(.A(n_324378252), .B(n_33195), .C(n_245877510), .D
		(n_31535), .Z(n_226577317));
	notech_ao3 i_130354687(.A(n_226377315), .B(n_226577317), .C(n_216277214)
		, .Z(n_226677318));
	notech_ao4 i_129854692(.A(n_324578254), .B(\nbus_11290[27] ), .C(n_5711)
		, .D(n_324478253), .Z(n_226777319));
	notech_ao4 i_129754693(.A(n_302978039), .B(nbus_11271[27]), .C(n_324678255
		), .D(\nbus_11283[27] ), .Z(n_226877320));
	notech_ao4 i_129454696(.A(n_284231523), .B(n_302878038), .C(n_175169787)
		, .D(n_303078040), .Z(n_227077322));
	notech_ao4 i_129354697(.A(n_324378252), .B(n_33198), .C(n_245877510), .D
		(n_31534), .Z(n_227277324));
	notech_ao3 i_129654694(.A(n_227077322), .B(n_227277324), .C(n_215377205)
		, .Z(n_227377325));
	notech_ao4 i_129154699(.A(n_324578254), .B(\nbus_11290[26] ), .C(n_5720)
		, .D(n_324478253), .Z(n_227477326));
	notech_ao4 i_129054700(.A(n_302978039), .B(nbus_11271[26]), .C(n_324678255
		), .D(\nbus_11283[26] ), .Z(n_227577327));
	notech_ao4 i_127254718(.A(n_4387), .B(n_124126568), .C(n_94229643), .D(n_337661004
		), .Z(n_227777329));
	notech_ao4 i_127054720(.A(n_57006), .B(n_31537), .C(n_328660914), .D(n_31505
		), .Z(n_227977331));
	notech_and4 i_127454716(.A(n_227977331), .B(n_227777329), .C(n_213977193
		), .D(n_214277196), .Z(n_228177333));
	notech_ao4 i_126754723(.A(n_124526572), .B(\nbus_11290[29] ), .C(n_4428)
		, .D(n_124826575), .Z(n_228277334));
	notech_ao4 i_126554725(.A(n_330460932), .B(n_33445), .C(n_337561003), .D
		(nbus_11271[29]), .Z(n_228477336));
	notech_and4 i_126954721(.A(n_228477336), .B(n_228277334), .C(n_213377187
		), .D(n_213677190), .Z(n_228677338));
	notech_ao4 i_126254728(.A(n_440082450), .B(n_124126568), .C(n_7636), .D(n_337661004
		), .Z(n_228777339));
	notech_ao4 i_126054730(.A(n_57006), .B(n_31536), .C(n_328660914), .D(n_31504
		), .Z(n_228977341));
	notech_and4 i_126454726(.A(n_228977341), .B(n_228777339), .C(n_212777181
		), .D(n_213077184), .Z(n_229177343));
	notech_ao4 i_125754733(.A(n_124526572), .B(\nbus_11290[28] ), .C(n_4427)
		, .D(n_124826575), .Z(n_229277344));
	notech_ao4 i_125554735(.A(n_330460932), .B(n_33444), .C(n_337561003), .D
		(nbus_11271[28]), .Z(n_229477346));
	notech_and4 i_125954731(.A(n_229477346), .B(n_229277344), .C(n_212177175
		), .D(n_212477178), .Z(n_229677348));
	notech_ao4 i_125254738(.A(n_284131522), .B(n_124126568), .C(n_172669762)
		, .D(n_337661004), .Z(n_229777349));
	notech_ao4 i_125054740(.A(n_57012), .B(n_31535), .C(n_328660914), .D(n_31503
		), .Z(n_229977351));
	notech_and4 i_125454736(.A(n_229977351), .B(n_229777349), .C(n_211577169
		), .D(n_211877172), .Z(n_230177353));
	notech_ao4 i_124754743(.A(n_124526572), .B(\nbus_11290[27] ), .C(n_5711)
		, .D(n_124826575), .Z(n_230277354));
	notech_ao4 i_124554745(.A(n_330460932), .B(n_33443), .C(n_337561003), .D
		(nbus_11271[27]), .Z(n_230477356));
	notech_and4 i_124954741(.A(n_230477356), .B(n_230277354), .C(n_210977163
		), .D(n_211277166), .Z(n_230677358));
	notech_ao4 i_124254748(.A(n_284231523), .B(n_124126568), .C(n_175169787)
		, .D(n_337661004), .Z(n_230777359));
	notech_ao4 i_124054750(.A(n_57012), .B(n_31534), .C(n_328660914), .D(n_31502
		), .Z(n_230977361));
	notech_and4 i_124454746(.A(n_230977361), .B(n_230777359), .C(n_210377157
		), .D(n_210677160), .Z(n_231177363));
	notech_ao4 i_123754753(.A(n_124526572), .B(\nbus_11290[26] ), .C(n_5720)
		, .D(n_124826575), .Z(n_231277364));
	notech_ao4 i_123554755(.A(n_55913), .B(n_33442), .C(n_337561003), .D(nbus_11271
		[26]), .Z(n_231477366));
	notech_and4 i_123954751(.A(n_231477366), .B(n_231277364), .C(n_209777151
		), .D(n_210077154), .Z(n_231677368));
	notech_ao4 i_115854830(.A(n_4387), .B(n_301522040), .C(n_94229643), .D(n_298922014
		), .Z(n_231777369));
	notech_ao4 i_115754831(.A(n_4428), .B(n_324278251), .C(n_324178250), .D(n_33197
		), .Z(n_231977371));
	notech_ao4 i_115454834(.A(n_57213), .B(\nbus_11283[29] ), .C(n_57217), .D
		(\nbus_11290[29] ), .Z(n_232177373));
	notech_and4 i_115654832(.A(n_5774), .B(n_232177373), .C(n_222077272), .D
		(n_208977143), .Z(n_232477376));
	notech_ao4 i_115054838(.A(n_440082450), .B(n_301522040), .C(n_7636), .D(n_298922014
		), .Z(n_232577377));
	notech_ao4 i_114954839(.A(n_4427), .B(n_324278251), .C(n_324178250), .D(n_33196
		), .Z(n_232777379));
	notech_ao4 i_114654842(.A(n_57213), .B(\nbus_11283[28] ), .C(n_57217), .D
		(\nbus_11290[28] ), .Z(n_232977381));
	notech_and4 i_114854840(.A(n_5774), .B(n_232977381), .C(n_30506), .D(n_208077135
		), .Z(n_233277384));
	notech_ao4 i_114254846(.A(n_284131522), .B(n_301522040), .C(n_172669762)
		, .D(n_298922014), .Z(n_233377385));
	notech_ao4 i_114154847(.A(n_5711), .B(n_324278251), .C(n_324178250), .D(n_33195
		), .Z(n_233577387));
	notech_nand3 i_114454844(.A(n_233377385), .B(n_233577387), .C(n_207777132
		), .Z(n_233677388));
	notech_ao4 i_113954849(.A(n_57213), .B(\nbus_11283[27] ), .C(n_57217), .D
		(\nbus_11290[27] ), .Z(n_233777389));
	notech_ao4 i_113554853(.A(n_284231523), .B(n_301522040), .C(n_175169787)
		, .D(n_298922014), .Z(n_234077392));
	notech_ao4 i_113454854(.A(n_5720), .B(n_324278251), .C(n_324178250), .D(n_33198
		), .Z(n_234277394));
	notech_ao4 i_113154857(.A(n_57213), .B(\nbus_11283[26] ), .C(n_57217), .D
		(\nbus_11290[26] ), .Z(n_234477396));
	notech_and4 i_113354855(.A(n_5774), .B(n_234477396), .C(n_65029351), .D(n_206477119
		), .Z(n_234777399));
	notech_ao4 i_108454904(.A(n_440082450), .B(n_58100), .C(n_7636), .D(n_242836107
		), .Z(n_234877400));
	notech_ao4 i_108254906(.A(n_60454), .B(n_31536), .C(n_385264383), .D(n_31504
		), .Z(n_235077402));
	notech_and4 i_108654902(.A(n_235077402), .B(n_234877400), .C(n_205777113
		), .D(n_206077116), .Z(n_235277404));
	notech_ao4 i_107954909(.A(n_57370), .B(\nbus_11290[28] ), .C(n_4427), .D
		(n_57325), .Z(n_235377405));
	notech_ao4 i_107854910(.A(n_32186), .B(n_33441), .C(n_248736166), .D(nbus_11271
		[28]), .Z(n_235577407));
	notech_nor2 i_49852577(.A(n_363350926), .B(n_442968013), .Z(n_235777409)
		);
	notech_ao3 i_49952576(.A(n_63774), .B(opc_10[25]), .C(n_442768011), .Z(n_236477416
		));
	notech_or4 i_2620760(.A(n_353367697), .B(n_257777629), .C(n_236477416), 
		.D(n_235777409), .Z(n_19718));
	notech_or4 i_56552515(.A(n_339561023), .B(n_2829), .C(n_444168025), .D(n_3464
		), .Z(n_236577417));
	notech_nao3 i_56652514(.A(opc_10[22]), .B(n_63758), .C(n_442768011), .Z(n_237277424
		));
	notech_nand3 i_2320757(.A(n_258577637), .B(n_237277424), .C(n_236577417)
		, .Z(n_19700));
	notech_nor2 i_70852373(.A(n_363350926), .B(n_443968023), .Z(n_237377425)
		);
	notech_ao3 i_70952372(.A(n_63774), .B(opc_10[25]), .C(n_444068024), .Z(n_238077432
		));
	notech_or4 i_2620984(.A(n_353367697), .B(n_259177643), .C(n_238077432), 
		.D(n_237377425), .Z(n_19022));
	notech_nor2 i_72452357(.A(n_364628688), .B(n_443968023), .Z(n_238177433)
		);
	notech_or2 i_71852363(.A(n_443668020), .B(nbus_11271[24]), .Z(n_238277434
		));
	notech_ao3 i_72352358(.A(n_57386), .B(opd[24]), .C(n_57141), .Z(n_238777439
		));
	notech_ao3 i_72552356(.A(n_63774), .B(opc_10[24]), .C(n_444068024), .Z(n_238877440
		));
	notech_or4 i_2520983(.A(n_259877650), .B(n_259577647), .C(n_238877440), 
		.D(n_238177433), .Z(n_19016));
	notech_nor2 i_90452181(.A(n_325325323), .B(n_363350926), .Z(n_238977441)
		);
	notech_ao3 i_90552180(.A(n_63774), .B(opc_10[25]), .C(n_315725234), .Z(n_239677448
		));
	notech_or4 i_2621080(.A(n_353367697), .B(n_260577657), .C(n_239677448), 
		.D(n_238977441), .Z(n_16373));
	notech_nor2 i_92052165(.A(n_325325323), .B(n_364628688), .Z(n_239777449)
		);
	notech_or2 i_91452171(.A(n_324978258), .B(nbus_11271[24]), .Z(n_239877450
		));
	notech_ao3 i_91952166(.A(n_57386), .B(opd[24]), .C(n_57616), .Z(n_240377455
		));
	notech_ao3 i_92152164(.A(n_63774), .B(opc_10[24]), .C(n_315725234), .Z(n_240477456
		));
	notech_or4 i_2521079(.A(n_261277664), .B(n_260977661), .C(n_240477456), 
		.D(n_239777449), .Z(n_16367));
	notech_or4 i_95252133(.A(n_340361031), .B(n_339561023), .C(n_444168025),
		 .D(n_3464), .Z(n_240577457));
	notech_nao3 i_95352132(.A(opc_10[22]), .B(n_63758), .C(n_315725234), .Z(n_241277464
		));
	notech_nand3 i_2321077(.A(n_262077672), .B(n_240577457), .C(n_241277464)
		, .Z(n_16355));
	notech_or2 i_124051850(.A(n_302878038), .B(n_363350926), .Z(n_241377465)
		);
	notech_nao3 i_123951851(.A(n_57386), .B(opd[25]), .C(n_57158), .Z(n_242077472
		));
	notech_nao3 i_124151849(.A(n_63774), .B(opc_10[25]), .C(n_303078040), .Z
		(n_242177473));
	notech_nand3 i_2621368(.A(n_262777679), .B(n_242177473), .C(n_241377465)
		, .Z(n_20534));
	notech_or2 i_125751833(.A(n_302878038), .B(n_364628688), .Z(n_242277474)
		);
	notech_nao3 i_125651834(.A(n_57392), .B(opd[24]), .C(n_57158), .Z(n_242977481
		));
	notech_nao3 i_125851832(.A(n_63774), .B(opc_10[24]), .C(n_303078040), .Z
		(n_243077482));
	notech_nand3 i_2521367(.A(n_263477686), .B(n_243077482), .C(n_242277474)
		, .Z(n_20528));
	notech_or2 i_127451816(.A(n_302878038), .B(n_363450925), .Z(n_243177483)
		);
	notech_nao3 i_127351817(.A(n_57392), .B(opd[23]), .C(n_57158), .Z(n_243877490
		));
	notech_nao3 i_127551815(.A(n_63774), .B(opc_10[23]), .C(n_303078040), .Z
		(n_243977491));
	notech_nand3 i_2421366(.A(n_265977693), .B(n_243977491), .C(n_243177483)
		, .Z(n_20522));
	notech_or2 i_129151799(.A(n_302878038), .B(n_3464), .Z(n_244077492));
	notech_nao3 i_129051800(.A(n_57392), .B(opd[22]), .C(n_57158), .Z(n_244777499
		));
	notech_ao3 i_129251798(.A(opc_10[22]), .B(n_63784), .C(n_303078040), .Z(n_244877500
		));
	notech_nao3 i_2321365(.A(n_266677700), .B(n_244077492), .C(n_244877500),
		 .Z(n_20516));
	notech_or2 i_130851782(.A(n_302878038), .B(n_3466), .Z(n_244977501));
	notech_nao3 i_130751783(.A(n_57386), .B(opd[21]), .C(n_57158), .Z(n_245677508
		));
	notech_nao3 i_130951781(.A(opc_10[21]), .B(n_63784), .C(n_303078040), .Z
		(n_245777509));
	notech_nand3 i_2221364(.A(n_268377707), .B(n_245777509), .C(n_244977501)
		, .Z(n_20510));
	notech_nand2 i_41758139(.A(n_30524), .B(n_61621), .Z(n_245877510));
	notech_or2 i_132551765(.A(n_346771358), .B(n_302878038), .Z(n_245977511)
		);
	notech_nao3 i_132451766(.A(n_57386), .B(opd[20]), .C(n_57158), .Z(n_246677518
		));
	notech_ao3 i_132651764(.A(opc_10[20]), .B(n_63784), .C(n_303078040), .Z(n_246777519
		));
	notech_nao3 i_2121363(.A(n_269077714), .B(n_245977511), .C(n_246777519),
		 .Z(n_20504));
	notech_nor2 i_149551595(.A(n_364628688), .B(n_387664407), .Z(n_246877520
		));
	notech_or2 i_148951601(.A(n_387564406), .B(nbus_11271[24]), .Z(n_246977521
		));
	notech_ao3 i_149451596(.A(n_57386), .B(opd[24]), .C(n_57086), .Z(n_247477526
		));
	notech_ao3 i_149651594(.A(n_63772), .B(opc_10[24]), .C(n_387764408), .Z(n_247577527
		));
	notech_or4 i_2521623(.A(n_270877720), .B(n_270577717), .C(n_247577527), 
		.D(n_246877520), .Z(n_13136));
	notech_or4 i_152751563(.A(n_2829), .B(n_2845), .C(n_444168025), .D(n_3464
		), .Z(n_247677528));
	notech_ao3 i_152851562(.A(opc_10[22]), .B(n_63754), .C(n_387764408), .Z(n_248377535
		));
	notech_nao3 i_2321621(.A(n_271777728), .B(n_247677528), .C(n_248377535),
		 .Z(n_13124));
	notech_nor2 i_172551365(.A(n_301522040), .B(n_363350926), .Z(n_248477536
		));
	notech_ao3 i_172651364(.A(n_63766), .B(opc_10[25]), .C(n_298922014), .Z(n_249177543
		));
	notech_or4 i_2621848(.A(n_353367697), .B(n_272377734), .C(n_249177543), 
		.D(n_248477536), .Z(n_12794));
	notech_or4 i_177551316(.A(n_340461032), .B(n_2845), .C(n_444168025), .D(n_3464
		), .Z(n_249277544));
	notech_nand3 i_177451317(.A(n_57395), .B(n_32210), .C(opd[22]), .Z(n_249877550
		));
	notech_nao3 i_177651315(.A(opc_10[22]), .B(n_63780), .C(n_298922014), .Z
		(n_249977551));
	notech_and4 i_2321845(.A(n_354467708), .B(n_273177742), .C(n_249977551),
		 .D(n_249277544), .Z(n_12776));
	notech_nor2 i_194151152(.A(n_58100), .B(n_363350926), .Z(n_250077552));
	notech_nand2 i_194051153(.A(sav_ecx[25]), .B(n_61873), .Z(n_250977561)
		);
	notech_ao3 i_194251151(.A(n_63766), .B(opc_10[25]), .C(n_242836107), .Z(n_251077562
		));
	notech_or4 i_2617016(.A(n_274077751), .B(n_273677747), .C(n_251077562), 
		.D(n_250077552), .Z(n_12085));
	notech_nor2 i_196251131(.A(n_58100), .B(n_364628688), .Z(n_251177563));
	notech_nand2 i_196151132(.A(sav_ecx[24]), .B(n_61873), .Z(n_252077572)
		);
	notech_ao3 i_196351130(.A(n_63766), .B(opc_10[24]), .C(n_242836107), .Z(n_252177573
		));
	notech_or4 i_2517015(.A(n_274977760), .B(n_274577756), .C(n_252177573), 
		.D(n_251177563), .Z(n_12079));
	notech_nor2 i_198451110(.A(n_58100), .B(n_363450925), .Z(n_252277574));
	notech_nand2 i_198351111(.A(sav_ecx[23]), .B(n_61873), .Z(n_253177583)
		);
	notech_ao3 i_198551109(.A(n_63766), .B(opc_10[23]), .C(n_242836107), .Z(n_253277584
		));
	notech_or4 i_2417014(.A(n_275877769), .B(n_275477765), .C(n_253277584), 
		.D(n_252277574), .Z(n_12073));
	notech_or2 i_202751067(.A(n_58100), .B(n_3466), .Z(n_253377585));
	notech_nao3 i_201851076(.A(\regs_1_0[21] ), .B(n_19680), .C(n_57012), .Z
		(n_253477586));
	notech_nao3 i_202851066(.A(opc_10[21]), .B(n_63784), .C(n_242836107), .Z
		(n_254377595));
	notech_nand3 i_2217012(.A(n_276977780), .B(n_254377595), .C(n_253377585)
		, .Z(n_12061));
	notech_nor2 i_204951045(.A(n_58100), .B(n_346771358), .Z(n_254477596));
	notech_nand2 i_204851046(.A(sav_ecx[20]), .B(n_61873), .Z(n_255377605)
		);
	notech_ao3 i_205051044(.A(opc_10[20]), .B(n_63784), .C(n_242836107), .Z(n_255477606
		));
	notech_or4 i_2117011(.A(n_277777788), .B(n_277377784), .C(n_255477606), 
		.D(n_254477596), .Z(n_12055));
	notech_nor2 i_206851026(.A(n_388064411), .B(n_363350926), .Z(n_255577607
		));
	notech_nao3 i_206751027(.A(n_57397), .B(opd[25]), .C(n_58701), .Z(n_256277614
		));
	notech_ao3 i_206951025(.A(n_63788), .B(opc_10[25]), .C(n_388164412), .Z(n_256377615
		));
	notech_or4 i_2617592(.A(n_353367697), .B(n_256377615), .C(n_255577607), 
		.D(n_30293), .Z(n_11716));
	notech_or4 i_210450990(.A(n_340361031), .B(n_2830), .C(n_444168025), .D(n_3464
		), .Z(n_256477616));
	notech_nao3 i_210350991(.A(n_57397), .B(opd[22]), .C(n_58701), .Z(n_257177623
		));
	notech_nao3 i_210550989(.A(opc_10[22]), .B(n_63784), .C(n_388164412), .Z
		(n_257277624));
	notech_and4 i_2317589(.A(n_279377804), .B(n_256477616), .C(n_354467708),
		 .D(n_257277624), .Z(n_11698));
	notech_ao4 i_50252573(.A(n_31501), .B(n_327960907), .C(n_117626503), .D(n_33172
		), .Z(n_257377625));
	notech_ao4 i_50052575(.A(n_442668010), .B(\nbus_11283[25] ), .C(n_442868012
		), .D(nbus_11271[25]), .Z(n_257477626));
	notech_ao4 i_50152574(.A(n_101026337), .B(n_117726504), .C(n_442568009),
		 .D(\nbus_11290[25] ), .Z(n_257577627));
	notech_nand3 i_50452571(.A(n_257577627), .B(n_257477626), .C(n_257377625
		), .Z(n_257777629));
	notech_ao4 i_56952511(.A(n_327960907), .B(n_31496), .C(n_117626503), .D(n_33284
		), .Z(n_258077632));
	notech_ao4 i_56752513(.A(n_442668010), .B(\nbus_11283[22] ), .C(n_442868012
		), .D(nbus_11271[22]), .Z(n_258177633));
	notech_ao4 i_56852512(.A(n_59464), .B(n_117726504), .C(n_442568009), .D(\nbus_11290[22] 
		), .Z(n_258277634));
	notech_and4 i_57252508(.A(n_258277634), .B(n_258177633), .C(n_258077632)
		, .D(n_354467708), .Z(n_258577637));
	notech_ao4 i_71252369(.A(n_31501), .B(n_379264323), .C(n_119226519), .D(n_33172
		), .Z(n_258777639));
	notech_ao4 i_71052371(.A(n_443768021), .B(\nbus_11283[25] ), .C(n_443668020
		), .D(nbus_11271[25]), .Z(n_258877640));
	notech_ao4 i_71152370(.A(n_101026337), .B(n_119326520), .C(n_443868022),
		 .D(\nbus_11290[25] ), .Z(n_258977641));
	notech_nand3 i_71452367(.A(n_258977641), .B(n_258877640), .C(n_258777639
		), .Z(n_259177643));
	notech_nao3 i_72952352(.A(n_238277434), .B(n_443068014), .C(n_238777439)
		, .Z(n_259577647));
	notech_ao4 i_72752354(.A(n_443868022), .B(\nbus_11290[24] ), .C(n_443768021
		), .D(\nbus_11283[24] ), .Z(n_259677648));
	notech_ao4 i_72852353(.A(n_119226519), .B(n_33171), .C(n_106826395), .D(n_119326520
		), .Z(n_259777649));
	notech_nand2 i_73052351(.A(n_259777649), .B(n_259677648), .Z(n_259877650
		));
	notech_ao4 i_90852177(.A(n_58088), .B(n_31501), .C(n_324778256), .D(n_33172
		), .Z(n_260177653));
	notech_ao4 i_90652179(.A(n_57201), .B(\nbus_11283[25] ), .C(n_324978258)
		, .D(nbus_11271[25]), .Z(n_260277654));
	notech_ao4 i_90752178(.A(n_324878257), .B(n_101026337), .C(n_57200), .D(\nbus_11290[25] 
		), .Z(n_260377655));
	notech_nand3 i_91052175(.A(n_260377655), .B(n_260277654), .C(n_260177653
		), .Z(n_260577657));
	notech_nao3 i_92552160(.A(n_443068014), .B(n_239877450), .C(n_240377455)
		, .Z(n_260977661));
	notech_ao4 i_92352162(.A(n_57200), .B(\nbus_11290[24] ), .C(n_57201), .D
		(\nbus_11283[24] ), .Z(n_261077662));
	notech_ao4 i_92452161(.A(n_324778256), .B(n_33171), .C(n_324878257), .D(n_106826395
		), .Z(n_261177663));
	notech_nand2 i_92652159(.A(n_261177663), .B(n_261077662), .Z(n_261277664
		));
	notech_ao4 i_95652129(.A(n_58088), .B(n_31496), .C(n_324778256), .D(n_33284
		), .Z(n_261577667));
	notech_ao4 i_95452131(.A(n_57201), .B(\nbus_11283[22] ), .C(n_324978258)
		, .D(nbus_11271[22]), .Z(n_261677668));
	notech_ao4 i_95552130(.A(n_324878257), .B(n_59464), .C(n_57200), .D(\nbus_11290[22] 
		), .Z(n_261777669));
	notech_and4 i_95952126(.A(n_261777669), .B(n_261677668), .C(n_261577667)
		, .D(n_354467708), .Z(n_262077672));
	notech_ao4 i_124251848(.A(n_324678255), .B(\nbus_11283[25] ), .C(n_302978039
		), .D(nbus_11271[25]), .Z(n_262277674));
	notech_ao4 i_124351847(.A(n_324478253), .B(n_101026337), .C(n_324578254)
		, .D(\nbus_11290[25] ), .Z(n_262477676));
	notech_ao4 i_124451846(.A(n_245877510), .B(n_31533), .C(n_324378252), .D
		(n_33172), .Z(n_262577677));
	notech_and4 i_124751843(.A(n_262577677), .B(n_262477676), .C(n_262277674
		), .D(n_242077472), .Z(n_262777679));
	notech_ao4 i_125951831(.A(n_324678255), .B(\nbus_11283[24] ), .C(n_302978039
		), .D(nbus_11271[24]), .Z(n_262977681));
	notech_ao4 i_126051830(.A(n_324478253), .B(n_106826395), .C(n_324578254)
		, .D(\nbus_11290[24] ), .Z(n_263177683));
	notech_ao4 i_126151829(.A(n_245877510), .B(n_31532), .C(n_324378252), .D
		(n_33171), .Z(n_263277684));
	notech_and4 i_126451826(.A(n_263277684), .B(n_263177683), .C(n_262977681
		), .D(n_242977481), .Z(n_263477686));
	notech_ao4 i_127651814(.A(n_324678255), .B(n_58420), .C(n_302978039), .D
		(n_60528), .Z(n_263677688));
	notech_ao4 i_127751813(.A(n_324478253), .B(n_109226419), .C(n_324578254)
		, .D(n_58902), .Z(n_263877690));
	notech_ao4 i_127851812(.A(n_245877510), .B(n_31531), .C(n_324378252), .D
		(n_33170), .Z(n_265177691));
	notech_and4 i_128151809(.A(n_265177691), .B(n_263877690), .C(n_263677688
		), .D(n_243877490), .Z(n_265977693));
	notech_ao4 i_129351797(.A(n_324678255), .B(\nbus_11283[22] ), .C(n_302978039
		), .D(nbus_11271[22]), .Z(n_266177695));
	notech_ao4 i_129451796(.A(n_324478253), .B(n_59464), .C(n_324578254), .D
		(\nbus_11290[22] ), .Z(n_266377697));
	notech_ao4 i_129551795(.A(n_245877510), .B(n_31530), .C(n_324378252), .D
		(n_33284), .Z(n_266477698));
	notech_and4 i_129851792(.A(n_266477698), .B(n_266377697), .C(n_266177695
		), .D(n_244777499), .Z(n_266677700));
	notech_ao4 i_131051780(.A(n_324678255), .B(n_58402), .C(n_302978039), .D
		(n_60546), .Z(n_267077702));
	notech_ao4 i_131151779(.A(n_324478253), .B(n_59465), .C(n_324578254), .D
		(n_58884), .Z(n_268077704));
	notech_ao4 i_131251778(.A(n_56783), .B(n_31529), .C(n_324378252), .D(n_33288
		), .Z(n_268177705));
	notech_and4 i_131551775(.A(n_268177705), .B(n_268077704), .C(n_267077702
		), .D(n_245677508), .Z(n_268377707));
	notech_ao4 i_132751763(.A(n_324678255), .B(n_58393), .C(n_302978039), .D
		(n_60555), .Z(n_268577709));
	notech_ao4 i_132851762(.A(n_324478253), .B(n_59466), .C(n_324578254), .D
		(n_58857), .Z(n_268777711));
	notech_ao4 i_132951761(.A(n_56783), .B(n_31528), .C(n_324378252), .D(n_33292
		), .Z(n_268877712));
	notech_and4 i_133251758(.A(n_268877712), .B(n_268777711), .C(n_268577709
		), .D(n_246677518), .Z(n_269077714));
	notech_nao3 i_150051590(.A(n_443068014), .B(n_246977521), .C(n_247477526
		), .Z(n_270577717));
	notech_ao4 i_149851592(.A(n_302844462), .B(\nbus_11290[24] ), .C(n_302744461
		), .D(\nbus_11283[24] ), .Z(n_270677718));
	notech_ao4 i_149951591(.A(n_125326580), .B(n_33171), .C(n_106826395), .D
		(n_125426581), .Z(n_270777719));
	notech_nand2 i_150151589(.A(n_270777719), .B(n_270677718), .Z(n_270877720
		));
	notech_ao4 i_153151559(.A(n_305644490), .B(n_31496), .C(n_125326580), .D
		(n_33284), .Z(n_271177723));
	notech_ao4 i_152951561(.A(n_302744461), .B(\nbus_11283[22] ), .C(n_387564406
		), .D(nbus_11271[22]), .Z(n_271277724));
	notech_ao4 i_153051560(.A(n_59464), .B(n_125426581), .C(n_302844462), .D
		(\nbus_11290[22] ), .Z(n_271377725));
	notech_and4 i_153451556(.A(n_271377725), .B(n_271277724), .C(n_271177723
		), .D(n_354467708), .Z(n_271777728));
	notech_ao4 i_172951361(.A(n_58083), .B(n_31501), .C(n_324178250), .D(n_33172
		), .Z(n_271977730));
	notech_ao4 i_172751363(.A(n_57213), .B(\nbus_11283[25] ), .C(n_301822043
		), .D(nbus_11271[25]), .Z(n_272077731));
	notech_ao4 i_172851362(.A(n_324278251), .B(n_101026337), .C(n_57217), .D
		(\nbus_11290[25] ), .Z(n_272177732));
	notech_nand3 i_173151359(.A(n_272177732), .B(n_272077731), .C(n_271977730
		), .Z(n_272377734));
	notech_ao4 i_177751314(.A(n_301822043), .B(nbus_11271[22]), .C(n_61621),
		 .D(n_383264363), .Z(n_272677737));
	notech_ao4 i_177851313(.A(n_57217), .B(n_58875), .C(n_57213), .D(\nbus_11283[22] 
		), .Z(n_272877739));
	notech_ao4 i_177951312(.A(n_324178250), .B(n_33284), .C(n_324278251), .D
		(n_59464), .Z(n_272977740));
	notech_and4 i_178251309(.A(n_272977740), .B(n_272877739), .C(n_272677737
		), .D(n_249877550), .Z(n_273177742));
	notech_ao4 i_194451149(.A(n_57370), .B(\nbus_11290[25] ), .C(n_57369), .D
		(\nbus_11283[25] ), .Z(n_273477745));
	notech_ao4 i_194551148(.A(n_57326), .B(n_33172), .C(n_57325), .D(n_101026337
		), .Z(n_273577746));
	notech_nand2 i_194851145(.A(n_273577746), .B(n_273477745), .Z(n_273677747
		));
	notech_ao4 i_194651147(.A(n_385264383), .B(n_31501), .C(n_60454), .D(n_31533
		), .Z(n_273777748));
	notech_ao4 i_194351150(.A(n_248736166), .B(nbus_11271[25]), .C(n_32186),
		 .D(n_33446), .Z(n_273877749));
	notech_nand3 i_194951144(.A(n_273877749), .B(n_273777748), .C(n_250977561
		), .Z(n_274077751));
	notech_ao4 i_196551128(.A(n_57370), .B(\nbus_11290[24] ), .C(n_57369), .D
		(\nbus_11283[24] ), .Z(n_274377754));
	notech_ao4 i_196651127(.A(n_57326), .B(n_33171), .C(n_57325), .D(n_106826395
		), .Z(n_274477755));
	notech_nand2 i_197051124(.A(n_274477755), .B(n_274377754), .Z(n_274577756
		));
	notech_ao4 i_196751126(.A(n_385264383), .B(n_31500), .C(n_60454), .D(n_31532
		), .Z(n_274677757));
	notech_ao4 i_196451129(.A(n_248736166), .B(nbus_11271[24]), .C(n_32186),
		 .D(n_33447), .Z(n_274777758));
	notech_nand3 i_197151123(.A(n_274777758), .B(n_274677757), .C(n_252077572
		), .Z(n_274977760));
	notech_ao4 i_198751107(.A(n_57370), .B(n_58902), .C(n_57369), .D(n_58420
		), .Z(n_275277763));
	notech_ao4 i_198851106(.A(n_57326), .B(n_33170), .C(n_57325), .D(n_109226419
		), .Z(n_275377764));
	notech_nand2 i_199151103(.A(n_275377764), .B(n_275277763), .Z(n_275477765
		));
	notech_ao4 i_198951105(.A(n_385264383), .B(n_31499), .C(n_60454), .D(n_31531
		), .Z(n_275577766));
	notech_ao4 i_198651108(.A(n_248736166), .B(n_60528), .C(n_32186), .D(n_33448
		), .Z(n_275677767));
	notech_nand3 i_199251102(.A(n_275677767), .B(n_275577766), .C(n_253177583
		), .Z(n_275877769));
	notech_ao4 i_203151063(.A(n_57325), .B(n_59465), .C(n_57370), .D(n_58884
		), .Z(n_276177772));
	notech_ao4 i_203251062(.A(n_60454), .B(n_31529), .C(n_57326), .D(n_33288
		), .Z(n_276277773));
	notech_ao4 i_203351061(.A(n_61106), .B(n_30773), .C(n_385264383), .D(n_31494
		), .Z(n_276477775));
	notech_ao4 i_203051064(.A(n_57369), .B(n_58402), .C(n_248736166), .D(n_60546
		), .Z(n_276677777));
	notech_and3 i_203451060(.A(n_58055), .B(n_276677777), .C(n_253477586), .Z
		(n_276777778));
	notech_and4 i_203751057(.A(n_276477775), .B(n_276277773), .C(n_276177772
		), .D(n_276777778), .Z(n_276977780));
	notech_ao4 i_205251042(.A(n_57370), .B(n_58857), .C(n_57369), .D(n_58393
		), .Z(n_277177782));
	notech_ao4 i_205351041(.A(n_57326), .B(n_33292), .C(n_57325), .D(n_59466
		), .Z(n_277277783));
	notech_nand2 i_205651038(.A(n_277277783), .B(n_277177782), .Z(n_277377784
		));
	notech_ao4 i_205451040(.A(n_385264383), .B(n_31493), .C(n_60454), .D(n_31528
		), .Z(n_277477785));
	notech_ao4 i_205151043(.A(n_248736166), .B(n_60555), .C(n_32186), .D(n_33449
		), .Z(n_277577786));
	notech_nand3 i_205751037(.A(n_277577786), .B(n_277477785), .C(n_255377605
		), .Z(n_277777788));
	notech_ao4 i_207051024(.A(n_131426641), .B(nbus_11271[25]), .C(n_56036),
		 .D(n_32552), .Z(n_278077791));
	notech_ao4 i_207151023(.A(n_387964410), .B(\nbus_11290[25] ), .C(n_387864409
		), .D(\nbus_11283[25] ), .Z(n_278277793));
	notech_ao4 i_207251022(.A(n_131526642), .B(n_33172), .C(n_131626643), .D
		(n_101026337), .Z(n_278377794));
	notech_and4 i_207551019(.A(n_278377794), .B(n_278277793), .C(n_278077791
		), .D(n_256277614), .Z(n_278577796));
	notech_ao4 i_210650988(.A(n_131426641), .B(nbus_11271[22]), .C(n_56036),
		 .D(n_32550), .Z(n_278877799));
	notech_ao4 i_210750987(.A(n_387964410), .B(n_58875), .C(n_387864409), .D
		(n_58411), .Z(n_279077801));
	notech_ao4 i_210850986(.A(n_131526642), .B(n_33284), .C(n_131626643), .D
		(n_59464), .Z(n_279177802));
	notech_and4 i_211150983(.A(n_279177802), .B(n_279077801), .C(n_278877799
		), .D(n_257177623), .Z(n_279377804));
	notech_or2 i_202458167(.A(n_56766), .B(n_280377814), .Z(n_279677807));
	notech_or4 i_199258168(.A(n_2382), .B(n_2580), .C(n_193276990), .D(n_280377814
		), .Z(n_279877809));
	notech_or4 i_40458203(.A(n_61912), .B(n_61901), .C(n_61889), .D(n_32181)
		, .Z(n_279977810));
	notech_or4 i_110266182(.A(n_2382), .B(n_2580), .C(n_193276990), .D(n_303978049
		), .Z(n_280077811));
	notech_or4 i_41658202(.A(n_61819), .B(n_30309), .C(n_57637), .D(n_57158)
		, .Z(n_280177812));
	notech_and4 i_349722(.A(n_116742608), .B(n_195877016), .C(n_335478360), 
		.D(n_323578244), .Z(n_280277813));
	notech_ao4 i_30358206(.A(n_32314), .B(n_57638), .C(n_30316), .D(n_32223)
		, .Z(n_280377814));
	notech_nand2 i_249723(.A(n_192776985), .B(n_303978049), .Z(n_280477815)
		);
	notech_and2 i_181558171(.A(n_194777005), .B(n_342578429), .Z(n_280777818
		));
	notech_ao4 i_26358209(.A(n_32314), .B(n_57638), .C(n_32227), .D(n_30316)
		, .Z(n_280977820));
	notech_or2 i_12249608(.A(n_57369), .B(\nbus_11283[17] ), .Z(n_281577826)
		);
	notech_or2 i_11949611(.A(n_57326), .B(n_33200), .Z(n_281877829));
	notech_nand2 i_11649614(.A(sav_ecx[17]), .B(n_61873), .Z(n_282177832));
	notech_or2 i_14449586(.A(n_57369), .B(\nbus_11283[19] ), .Z(n_282677837)
		);
	notech_or2 i_14149589(.A(n_57326), .B(n_33202), .Z(n_282977840));
	notech_nand2 i_13849592(.A(sav_ecx[19]), .B(n_61873), .Z(n_283277843));
	notech_nor2 i_21649514(.A(n_301822043), .B(nbus_11271[16]), .Z(n_283377844
		));
	notech_nand3 i_21149519(.A(n_57397), .B(n_32210), .C(opd[16]), .Z(n_284077851
		));
	notech_or2 i_22449506(.A(n_301822043), .B(nbus_11271[17]), .Z(n_284377854
		));
	notech_nand3 i_21949511(.A(n_57397), .B(n_32210), .C(opd[17]), .Z(n_284877859
		));
	notech_or2 i_23649498(.A(n_301822043), .B(nbus_11271[18]), .Z(n_285177862
		));
	notech_nand3 i_22749503(.A(n_57397), .B(n_32210), .C(opd[18]), .Z(n_285677867
		));
	notech_or2 i_24449490(.A(n_301822043), .B(nbus_11271[19]), .Z(n_285977870
		));
	notech_nand3 i_23949495(.A(n_57397), .B(n_32210), .C(opd[19]), .Z(n_286477875
		));
	notech_nao3 i_38649360(.A(n_164196010), .B(n_2645), .C(n_163296016), .Z(n_286577876
		));
	notech_nao3 i_39849348(.A(n_164196010), .B(n_2671), .C(n_163296016), .Z(n_288277893
		));
	notech_nand2 i_39549351(.A(sav_esi[16]), .B(n_61873), .Z(n_288577896));
	notech_or2 i_39249354(.A(n_124626573), .B(\nbus_11283[16] ), .Z(n_288877899
		));
	notech_or2 i_38949357(.A(n_320051171), .B(n_124126568), .Z(n_289177902)
		);
	notech_nao3 i_41049336(.A(n_164196010), .B(n_2673), .C(n_163296016), .Z(n_289477905
		));
	notech_nand2 i_40749339(.A(sav_esi[17]), .B(n_61873), .Z(n_289777908));
	notech_or2 i_40449342(.A(n_124626573), .B(\nbus_11283[17] ), .Z(n_290077911
		));
	notech_or2 i_40149345(.A(n_319951172), .B(n_124126568), .Z(n_290377914)
		);
	notech_nao3 i_42249324(.A(n_164196010), .B(n_2675), .C(n_163296016), .Z(n_290677917
		));
	notech_nand2 i_41949327(.A(sav_esi[18]), .B(n_61873), .Z(n_290977920));
	notech_or2 i_41649330(.A(n_124626573), .B(\nbus_11283[18] ), .Z(n_291277923
		));
	notech_or2 i_41349333(.A(n_319825274), .B(n_124126568), .Z(n_291577926)
		);
	notech_nao3 i_43449312(.A(n_164196010), .B(n_2677), .C(n_163296016), .Z(n_291877929
		));
	notech_nand2 i_43149315(.A(sav_esi[19]), .B(n_61873), .Z(n_292177932));
	notech_or2 i_42849318(.A(n_124626573), .B(\nbus_11283[19] ), .Z(n_292477935
		));
	notech_or2 i_42549321(.A(n_319725273), .B(n_124126568), .Z(n_292777938)
		);
	notech_nand2 i_44949297(.A(n_57950), .B(opa[3]), .Z(n_293077941));
	notech_or2 i_45249294(.A(n_267385090), .B(n_57158), .Z(n_295177962));
	notech_or2 i_46149285(.A(n_266585082), .B(n_57158), .Z(n_296077971));
	notech_or2 i_47049276(.A(n_265785074), .B(n_57158), .Z(n_296977980));
	notech_or2 i_48049267(.A(n_57157), .B(n_305478064), .Z(n_297877989));
	notech_nor2 i_62249130(.A(n_57201), .B(\nbus_11283[16] ), .Z(n_297977990
		));
	notech_or2 i_61749135(.A(n_5444), .B(n_324878257), .Z(n_298677997));
	notech_nor2 i_63049122(.A(n_57201), .B(\nbus_11283[17] ), .Z(n_298777998
		));
	notech_or2 i_62549127(.A(n_5397), .B(n_324878257), .Z(n_299478005));
	notech_nor2 i_63849114(.A(n_57201), .B(\nbus_11283[18] ), .Z(n_299578006
		));
	notech_or2 i_63349119(.A(n_5436), .B(n_324878257), .Z(n_300378013));
	notech_nor2 i_64649106(.A(n_57201), .B(\nbus_11283[19] ), .Z(n_300478014
		));
	notech_or2 i_64149111(.A(n_5356), .B(n_324878257), .Z(n_301178021));
	notech_or2 i_31653(.A(n_444168025), .B(n_57147), .Z(n_302878038));
	notech_nao3 i_2049705(.A(n_63788), .B(n_30315), .C(n_280377814), .Z(n_302978039
		));
	notech_nand2 i_2349702(.A(n_280477815), .B(n_30315), .Z(n_303078040));
	notech_or4 i_202858166(.A(n_2382), .B(n_2580), .C(n_193276990), .D(n_192776985
		), .Z(n_303178041));
	notech_or2 i_110166183(.A(n_56766), .B(n_303978049), .Z(n_303378043));
	notech_nor2 i_118948592(.A(n_280777818), .B(n_336360991), .Z(n_303578045
		));
	notech_ao4 i_223847555(.A(n_57679), .B(n_280777818), .C(n_56766), .D(n_303978049
		), .Z(n_303778047));
	notech_ao4 i_223747556(.A(n_30689), .B(eval_flag), .C(n_192776985), .D(n_56747
		), .Z(n_303878048));
	notech_and3 i_112566179(.A(n_116742608), .B(n_195677014), .C(n_195177009
		), .Z(n_303978049));
	notech_ao4 i_198147812(.A(n_242970425), .B(n_31125), .C(n_31123), .D(n_242870424
		), .Z(n_304078050));
	notech_ao4 i_198047813(.A(n_243270428), .B(n_31126), .C(n_243170427), .D
		(n_31122), .Z(n_304178051));
	notech_ao4 i_197847815(.A(n_262170616), .B(n_31099), .C(n_57441), .D(n_31098
		), .Z(n_304378053));
	notech_ao4 i_197747816(.A(n_31119), .B(n_249970494), .C(n_31118), .D(n_249870493
		), .Z(n_304478054));
	notech_and4 i_198347810(.A(n_304478054), .B(n_304378053), .C(n_304178051
		), .D(n_304078050), .Z(n_304678056));
	notech_ao4 i_197447819(.A(n_321271180), .B(n_334960977), .C(n_30326), .D
		(n_33458), .Z(n_304778057));
	notech_ao4 i_197347820(.A(n_57034), .B(n_33457), .C(n_61106), .D(n_30870
		), .Z(n_304878058));
	notech_ao4 i_197147822(.A(n_58042), .B(n_31478), .C(n_318971160), .D(n_31513
		), .Z(n_305078060));
	notech_ao4 i_197047823(.A(n_309771080), .B(n_33135), .C(n_309671079), .D
		(n_334860976), .Z(n_305178061));
	notech_and4 i_197647817(.A(n_305178061), .B(n_305078060), .C(n_304878058
		), .D(n_304778057), .Z(n_305378063));
	notech_or2 i_649719(.A(n_319725273), .B(n_444168025), .Z(n_305478064));
	notech_ao4 i_173948054(.A(n_57616), .B(n_305478064), .C(n_232870324), .D
		(n_315725234), .Z(n_305578065));
	notech_ao4 i_173848055(.A(n_324978258), .B(nbus_11271[19]), .C(n_324778256
		), .D(n_33202), .Z(n_305778067));
	notech_nand3 i_174148052(.A(n_305578065), .B(n_305778067), .C(n_301178021
		), .Z(n_305878068));
	notech_ao4 i_173648057(.A(n_57200), .B(\nbus_11290[19] ), .C(n_58088), .D
		(n_31492), .Z(n_305978069));
	notech_ao4 i_173248061(.A(n_265785074), .B(n_57616), .C(n_235370349), .D
		(n_315725234), .Z(n_306278072));
	notech_ao4 i_173148062(.A(n_324978258), .B(nbus_11271[18]), .C(n_324778256
		), .D(n_33201), .Z(n_306478074));
	notech_nand3 i_173448059(.A(n_306278072), .B(n_306478074), .C(n_300378013
		), .Z(n_306578075));
	notech_ao4 i_172948064(.A(n_57200), .B(\nbus_11290[18] ), .C(n_58088), .D
		(n_31491), .Z(n_306678076));
	notech_ao4 i_172548068(.A(n_266585082), .B(n_57616), .C(n_237870374), .D
		(n_315725234), .Z(n_306978079));
	notech_ao4 i_172448069(.A(n_324978258), .B(nbus_11271[17]), .C(n_324778256
		), .D(n_33200), .Z(n_307178081));
	notech_nand3 i_172748066(.A(n_306978079), .B(n_307178081), .C(n_299478005
		), .Z(n_307278082));
	notech_ao4 i_172248071(.A(n_57200), .B(\nbus_11290[17] ), .C(n_58088), .D
		(n_31490), .Z(n_307378083));
	notech_ao4 i_171848075(.A(n_267385090), .B(n_57616), .C(n_240370399), .D
		(n_315725234), .Z(n_307678086));
	notech_ao4 i_171748076(.A(n_324978258), .B(nbus_11271[16]), .C(n_324778256
		), .D(n_33199), .Z(n_307878088));
	notech_nand3 i_172048073(.A(n_307678086), .B(n_307878088), .C(n_298677997
		), .Z(n_307978089));
	notech_ao4 i_171548078(.A(n_57200), .B(\nbus_11290[16] ), .C(n_58088), .D
		(n_31489), .Z(n_308078090));
	notech_ao4 i_160648187(.A(n_302978039), .B(nbus_11271[19]), .C(n_232870324
		), .D(n_303078040), .Z(n_308378093));
	notech_ao4 i_160548188(.A(n_324378252), .B(n_33202), .C(n_5356), .D(n_324478253
		), .Z(n_308578095));
	notech_and3 i_160848185(.A(n_308378093), .B(n_308578095), .C(n_297877989
		), .Z(n_308678096));
	notech_ao4 i_160348190(.A(n_324678255), .B(\nbus_11283[19] ), .C(n_324578254
		), .D(\nbus_11290[19] ), .Z(n_308778097));
	notech_ao4 i_160248191(.A(n_56783), .B(n_31527), .C(n_31492), .D(n_280177812
		), .Z(n_308878098));
	notech_ao4 i_159948194(.A(n_302978039), .B(nbus_11271[18]), .C(n_235370349
		), .D(n_303078040), .Z(n_309078100));
	notech_ao4 i_159848195(.A(n_324378252), .B(n_33201), .C(n_5436), .D(n_324478253
		), .Z(n_309278102));
	notech_and3 i_160148192(.A(n_309078100), .B(n_309278102), .C(n_296977980
		), .Z(n_309378103));
	notech_ao4 i_159648197(.A(n_324678255), .B(\nbus_11283[18] ), .C(n_324578254
		), .D(\nbus_11290[18] ), .Z(n_309478104));
	notech_ao4 i_159548198(.A(n_56783), .B(n_31526), .C(n_280177812), .D(n_31491
		), .Z(n_309578105));
	notech_ao4 i_159248201(.A(n_302978039), .B(nbus_11271[17]), .C(n_237870374
		), .D(n_303078040), .Z(n_309778107));
	notech_ao4 i_159148202(.A(n_33200), .B(n_324378252), .C(n_5397), .D(n_324478253
		), .Z(n_309978109));
	notech_and3 i_159448199(.A(n_309778107), .B(n_309978109), .C(n_296077971
		), .Z(n_310078110));
	notech_ao4 i_158948204(.A(n_324678255), .B(\nbus_11283[17] ), .C(n_324578254
		), .D(\nbus_11290[17] ), .Z(n_310178111));
	notech_ao4 i_158848205(.A(n_56783), .B(n_31525), .C(n_280177812), .D(n_31490
		), .Z(n_310278112));
	notech_ao4 i_158548208(.A(n_302978039), .B(nbus_11271[16]), .C(n_240370399
		), .D(n_303078040), .Z(n_310478114));
	notech_ao4 i_158448209(.A(n_324378252), .B(n_33199), .C(n_5444), .D(n_324478253
		), .Z(n_310678116));
	notech_and3 i_158748206(.A(n_310478114), .B(n_310678116), .C(n_295177962
		), .Z(n_310778117));
	notech_ao4 i_158248211(.A(n_324678255), .B(\nbus_11283[16] ), .C(n_324578254
		), .D(\nbus_11290[16] ), .Z(n_310878118));
	notech_ao4 i_158148212(.A(n_56783), .B(n_31524), .C(n_280177812), .D(n_31489
		), .Z(n_310978119));
	notech_ao4 i_157848215(.A(n_74922852), .B(n_200977065), .C(n_66222765), 
		.D(n_57147), .Z(n_311178121));
	notech_ao4 i_157748216(.A(n_75322856), .B(n_178676846), .C(n_75222855), 
		.D(n_178576845), .Z(n_311278122));
	notech_ao4 i_157548218(.A(n_75522858), .B(n_178476844), .C(n_75622859), 
		.D(n_178776847), .Z(n_311478124));
	notech_ao4 i_157448219(.A(n_74622849), .B(n_57432), .C(n_74822851), .D(n_178376843
		), .Z(n_311578125));
	notech_and4 i_158048213(.A(n_311578125), .B(n_311478124), .C(n_311278122
		), .D(n_311178121), .Z(n_311778127));
	notech_ao4 i_157148222(.A(n_178876848), .B(n_31511), .C(n_74522848), .D(n_200877064
		), .Z(n_311878128));
	notech_ao4 i_157048223(.A(n_338361011), .B(n_57289), .C(n_31476), .D(n_58019
		), .Z(n_311978129));
	notech_ao4 i_156848225(.A(n_197877035), .B(\nbus_11290[3] ), .C(n_33118)
		, .D(n_57010), .Z(n_312178131));
	notech_and4 i_157348220(.A(n_312178131), .B(n_311978129), .C(n_311878128
		), .D(n_293077941), .Z(n_312378133));
	notech_ao4 i_156548228(.A(n_232870324), .B(n_337661004), .C(n_337561003)
		, .D(nbus_11271[19]), .Z(n_312478134));
	notech_ao4 i_156348230(.A(n_124726574), .B(n_33202), .C(n_5356), .D(n_124826575
		), .Z(n_312678136));
	notech_and4 i_156748226(.A(n_312678136), .B(n_312478134), .C(n_292477935
		), .D(n_292777938), .Z(n_312878138));
	notech_ao4 i_156048233(.A(n_328660914), .B(n_31492), .C(n_124526572), .D
		(\nbus_11290[19] ), .Z(n_312978139));
	notech_ao4 i_155848235(.A(n_55913), .B(n_33456), .C(n_57012), .D(n_31527
		), .Z(n_313178141));
	notech_and4 i_156248231(.A(n_313178141), .B(n_312978139), .C(n_291877929
		), .D(n_292177932), .Z(n_313378143));
	notech_ao4 i_155548238(.A(n_235370349), .B(n_337661004), .C(n_337561003)
		, .D(nbus_11271[18]), .Z(n_313478144));
	notech_ao4 i_155348240(.A(n_124726574), .B(n_33201), .C(n_5436), .D(n_124826575
		), .Z(n_313678146));
	notech_and4 i_155748236(.A(n_313678146), .B(n_313478144), .C(n_291277923
		), .D(n_291577926), .Z(n_313878148));
	notech_ao4 i_155048243(.A(n_328660914), .B(n_31491), .C(n_124526572), .D
		(\nbus_11290[18] ), .Z(n_313978149));
	notech_ao4 i_154848245(.A(n_55913), .B(n_33455), .C(n_57012), .D(n_31526
		), .Z(n_314178151));
	notech_and4 i_155248241(.A(n_314178151), .B(n_313978149), .C(n_290677917
		), .D(n_290977920), .Z(n_314378153));
	notech_ao4 i_154548248(.A(n_237870374), .B(n_337661004), .C(n_337561003)
		, .D(nbus_11271[17]), .Z(n_314478154));
	notech_ao4 i_154348250(.A(n_33200), .B(n_124726574), .C(n_5397), .D(n_124826575
		), .Z(n_314678156));
	notech_and4 i_154748246(.A(n_314678156), .B(n_314478154), .C(n_290077911
		), .D(n_290377914), .Z(n_314878158));
	notech_ao4 i_154048253(.A(n_328660914), .B(n_31490), .C(n_124526572), .D
		(\nbus_11290[17] ), .Z(n_314978159));
	notech_ao4 i_153848255(.A(n_55913), .B(n_33454), .C(n_57012), .D(n_31525
		), .Z(n_315178161));
	notech_and4 i_154248251(.A(n_315178161), .B(n_314978159), .C(n_289477905
		), .D(n_289777908), .Z(n_315378163));
	notech_ao4 i_153548258(.A(n_240370399), .B(n_337661004), .C(n_337561003)
		, .D(nbus_11271[16]), .Z(n_315478164));
	notech_ao4 i_153348260(.A(n_124726574), .B(n_33199), .C(n_5444), .D(n_124826575
		), .Z(n_315678166));
	notech_and4 i_153748256(.A(n_315678166), .B(n_315478164), .C(n_288877899
		), .D(n_289177902), .Z(n_315878168));
	notech_ao4 i_153048263(.A(n_328660914), .B(n_31489), .C(n_124526572), .D
		(\nbus_11290[16] ), .Z(n_315978169));
	notech_ao4 i_152848265(.A(n_55913), .B(n_33453), .C(n_57012), .D(n_31524
		), .Z(n_316178171));
	notech_and4 i_153248261(.A(n_316178171), .B(n_315978169), .C(n_288277893
		), .D(n_288577896), .Z(n_316378173));
	notech_ao4 i_152548268(.A(n_75222855), .B(n_139676462), .C(n_74922852), 
		.D(n_139276458), .Z(n_316478174));
	notech_ao4 i_152448269(.A(n_139376459), .B(n_75622859), .C(n_75322856), 
		.D(n_139476460), .Z(n_316578175));
	notech_ao4 i_152248271(.A(n_74822851), .B(n_116576231), .C(n_139576461),
		 .D(n_75522858), .Z(n_316778177));
	notech_ao4 i_152148272(.A(n_74522848), .B(n_139176457), .C(n_74622849), 
		.D(n_57439), .Z(n_316878178));
	notech_and4 i_152748266(.A(n_316878178), .B(n_316778177), .C(n_316578175
		), .D(n_316478174), .Z(n_317078180));
	notech_ao4 i_151848275(.A(n_61106), .B(n_30812), .C(n_338161009), .D(n_328760915
		), .Z(n_317178181));
	notech_ao4 i_151748276(.A(n_338361011), .B(n_57276), .C(n_31476), .D(n_58040
		), .Z(n_317278182));
	notech_ao4 i_151548278(.A(n_55913), .B(n_33452), .C(n_57277), .D(n_33118
		), .Z(n_317478184));
	notech_and4 i_151648277(.A(n_349581961), .B(n_246070456), .C(n_317478184
		), .D(n_286577876), .Z(n_317678186));
	notech_ao4 i_140548382(.A(n_319725273), .B(n_301522040), .C(n_232870324)
		, .D(n_298922014), .Z(n_317878188));
	notech_ao4 i_140448383(.A(n_5356), .B(n_324278251), .C(n_324178250), .D(n_33202
		), .Z(n_318078190));
	notech_ao4 i_140148386(.A(n_57213), .B(\nbus_11283[19] ), .C(n_57217), .D
		(\nbus_11290[19] ), .Z(n_318278192));
	notech_and4 i_140348384(.A(n_5774), .B(n_318278192), .C(n_285977870), .D
		(n_30510), .Z(n_318578195));
	notech_ao4 i_139748390(.A(n_319825274), .B(n_301522040), .C(n_235370349)
		, .D(n_298922014), .Z(n_318678196));
	notech_ao4 i_139648391(.A(n_5436), .B(n_324278251), .C(n_324178250), .D(n_33201
		), .Z(n_318878198));
	notech_ao4 i_139348394(.A(n_57213), .B(\nbus_11283[18] ), .C(n_57217), .D
		(\nbus_11290[18] ), .Z(n_319078200));
	notech_and4 i_139548392(.A(n_5774), .B(n_319078200), .C(n_285177862), .D
		(n_30511), .Z(n_319378203));
	notech_ao4 i_138948398(.A(n_319951172), .B(n_301522040), .C(n_237870374)
		, .D(n_298922014), .Z(n_319478204));
	notech_ao4 i_138848399(.A(n_5397), .B(n_324278251), .C(n_33200), .D(n_324178250
		), .Z(n_319678206));
	notech_ao4 i_138548402(.A(n_57213), .B(\nbus_11283[17] ), .C(n_57217), .D
		(\nbus_11290[17] ), .Z(n_319878208));
	notech_and4 i_138748400(.A(n_5774), .B(n_319878208), .C(n_284377854), .D
		(n_30512), .Z(n_320178211));
	notech_ao4 i_138148406(.A(n_320051171), .B(n_301522040), .C(n_240370399)
		, .D(n_298922014), .Z(n_320278212));
	notech_ao4 i_138048407(.A(n_5444), .B(n_324278251), .C(n_324178250), .D(n_33199
		), .Z(n_320478214));
	notech_nand3 i_138348404(.A(n_320278212), .B(n_320478214), .C(n_284077851
		), .Z(n_320578215));
	notech_ao4 i_137848409(.A(n_57213), .B(\nbus_11283[16] ), .C(n_57217), .D
		(\nbus_11290[16] ), .Z(n_320678216));
	notech_ao4 i_130948472(.A(n_319725273), .B(n_58100), .C(n_232870324), .D
		(n_242836107), .Z(n_320978219));
	notech_ao4 i_130748474(.A(n_60454), .B(n_31527), .C(n_385264383), .D(n_31492
		), .Z(n_321278221));
	notech_and4 i_131148470(.A(n_321278221), .B(n_320978219), .C(n_282977840
		), .D(n_283277843), .Z(n_321478223));
	notech_ao4 i_130448477(.A(n_57370), .B(\nbus_11290[19] ), .C(n_5356), .D
		(n_57325), .Z(n_321578224));
	notech_ao4 i_130348478(.A(n_32186), .B(n_33451), .C(n_248736166), .D(nbus_11271
		[19]), .Z(n_321778226));
	notech_ao4 i_129048491(.A(n_319951172), .B(n_58100), .C(n_237870374), .D
		(n_242836107), .Z(n_321978228));
	notech_ao4 i_128848493(.A(n_60454), .B(n_31525), .C(n_385264383), .D(n_31490
		), .Z(n_322178230));
	notech_and4 i_129248489(.A(n_322178230), .B(n_321978228), .C(n_281877829
		), .D(n_282177832), .Z(n_322378232));
	notech_ao4 i_128548496(.A(n_57370), .B(\nbus_11290[17] ), .C(n_5397), .D
		(n_57325), .Z(n_322478233));
	notech_ao4 i_128448497(.A(n_32186), .B(n_33450), .C(n_248736166), .D(nbus_11271
		[17]), .Z(n_322678235));
	notech_nao3 i_120763386(.A(n_58555), .B(n_30646), .C(n_57450), .Z(n_322878237
		));
	notech_or4 i_120663387(.A(n_256563512), .B(n_57450), .C(n_32159), .D(n_32269
		), .Z(n_322978238));
	notech_nao3 i_122563385(.A(n_201377069), .B(n_57627), .C(n_285763759), .Z
		(n_323078239));
	notech_nao3 i_122458185(.A(n_201377069), .B(n_32252), .C(n_285763759), .Z
		(n_323178240));
	notech_or4 i_89058194(.A(n_338661014), .B(n_318160809), .C(n_335478360),
		 .D(n_285763759), .Z(n_323278241));
	notech_or4 i_151358176(.A(n_338661014), .B(n_318160809), .C(n_285763759)
		, .D(n_323578244), .Z(n_323378242));
	notech_or2 i_151658175(.A(n_376064291), .B(n_323578244), .Z(n_323478243)
		);
	notech_ao4 i_28358207(.A(n_57679), .B(n_32314), .C(n_30719), .D(n_32227)
		, .Z(n_323578244));
	notech_or4 i_9763(.A(n_32269), .B(n_178276842), .C(n_32159), .D(n_256563512
		), .Z(n_323678245));
	notech_or4 i_146960745(.A(n_32269), .B(n_324078249), .C(n_32159), .D(n_256563512
		), .Z(n_323778246));
	notech_nor2 i_9765(.A(n_376364294), .B(n_178276842), .Z(n_323878247));
	notech_or2 i_147060744(.A(n_376364294), .B(n_324078249), .Z(n_323978248)
		);
	notech_ao4 i_28260786(.A(n_57679), .B(n_57566), .C(n_30719), .D(n_32210)
		, .Z(n_324078249));
	notech_ao3 i_114946490(.A(n_57027), .B(n_323978248), .C(n_323878247), .Z
		(n_324178250));
	notech_and3 i_115046491(.A(n_57036), .B(n_323678245), .C(n_323778246), .Z
		(n_324278251));
	notech_ao3 i_118249758(.A(n_303778047), .B(n_56720), .C(n_303578045), .Z
		(n_324378252));
	notech_and2 i_118349757(.A(n_280077811), .B(n_303878048), .Z(n_324478253
		));
	notech_ao4 i_113849776(.A(n_193176989), .B(n_30694), .C(n_280377814), .D
		(n_56747), .Z(n_324578254));
	notech_ao4 i_113749777(.A(n_57638), .B(n_194577003), .C(n_56766), .D(n_280377814
		), .Z(n_324678255));
	notech_ao3 i_115549768(.A(n_192676984), .B(n_323478243), .C(n_116876234)
		, .Z(n_324778256));
	notech_and3 i_115649767(.A(n_323278241), .B(n_116776233), .C(n_323378242
		), .Z(n_324878257));
	notech_ao4 i_113949775(.A(n_280977820), .B(n_375764288), .C(n_32181), .D
		(n_61621), .Z(n_324978258));
	notech_and4 i_88845566(.A(n_116742608), .B(n_180276862), .C(n_324078249)
		, .D(n_58208), .Z(n_325078259));
	notech_nand2 i_103945417(.A(n_115442595), .B(n_32227), .Z(n_325178260)
		);
	notech_nao3 i_104045416(.A(n_57627), .B(n_30642), .C(n_335478360), .Z(n_325278261
		));
	notech_nand2 i_104745410(.A(n_115442595), .B(n_32210), .Z(n_325578264)
		);
	notech_nao3 i_104845409(.A(n_58555), .B(n_30646), .C(n_58208), .Z(n_325678265
		));
	notech_or2 i_36546053(.A(n_57369), .B(\nbus_11283[31] ), .Z(n_326178270)
		);
	notech_or2 i_36246056(.A(n_57326), .B(n_33206), .Z(n_326478273));
	notech_nand2 i_35946059(.A(sav_ecx[31]), .B(n_61873), .Z(n_326778276));
	notech_or4 i_39846021(.A(n_256563512), .B(n_324078249), .C(n_5269), .D(n_58555
		), .Z(n_326878277));
	notech_or2 i_39746022(.A(n_323978248), .B(n_33253), .Z(n_327178280));
	notech_or2 i_39446025(.A(n_58030), .B(n_31481), .Z(n_327478283));
	notech_or4 i_39046028(.A(n_63698), .B(n_57393), .C(n_63784), .D(nbus_11273
		[8]), .Z(n_327778286));
	notech_nor2 i_40646013(.A(n_57213), .B(\nbus_11283[31] ), .Z(n_327878287
		));
	notech_or2 i_40146018(.A(n_301822043), .B(nbus_11271[31]), .Z(n_328578294
		));
	notech_nao3 i_47845953(.A(n_164196010), .B(n_2655), .C(n_163296016), .Z(n_328878297
		));
	notech_or2 i_47045960(.A(n_5269), .B(n_57275), .Z(n_329578304));
	notech_nao3 i_49145941(.A(n_164196010), .B(n_2701), .C(n_163296016), .Z(n_330278311
		));
	notech_or2 i_48845944(.A(n_124626573), .B(\nbus_11283[31] ), .Z(n_330578314
		));
	notech_or2 i_48545947(.A(n_124726574), .B(n_33206), .Z(n_331078317));
	notech_nand2 i_48145950(.A(sav_esi[31]), .B(n_61873), .Z(n_331378320));
	notech_ao3 i_50845924(.A(n_57397), .B(opd[31]), .C(n_57147), .Z(n_332278329
		));
	notech_nor2 i_59945835(.A(n_324978258), .B(nbus_11271[31]), .Z(n_332378330
		));
	notech_nand3 i_59445840(.A(n_57397), .B(n_32227), .C(opd[31]), .Z(n_333078337
		));
	notech_or2 i_66945768(.A(n_30496), .B(\nbus_11290[8] ), .Z(n_333678342)
		);
	notech_nao3 i_33484(.A(n_28557), .B(n_273263663), .C(n_57393), .Z(n_333778343
		));
	notech_or2 i_33483(.A(n_57393), .B(n_26063), .Z(n_333878344));
	notech_nao3 i_33481(.A(n_28557), .B(n_273263663), .C(n_324078249), .Z(n_333978345
		));
	notech_or2 i_32203(.A(n_57394), .B(n_30549), .Z(n_334078346));
	notech_or2 i_32201(.A(n_83739557), .B(n_30549), .Z(n_334178347));
	notech_or2 i_32200(.A(n_57394), .B(n_27378), .Z(n_334278348));
	notech_nao3 i_30319(.A(n_33173), .B(n_286063762), .C(n_57387), .Z(n_334378349
		));
	notech_or2 i_30318(.A(n_57387), .B(n_29214), .Z(n_334478350));
	notech_nand3 i_30317(.A(n_33173), .B(n_286063762), .C(n_30300), .Z(n_334578351
		));
	notech_nao3 i_120266177(.A(n_116676232), .B(n_32243), .C(n_163196017), .Z
		(n_334778353));
	notech_nao3 i_120366176(.A(n_57461), .B(n_116676232), .C(n_163196017), .Z
		(n_334878354));
	notech_nao3 i_104645411(.A(n_57461), .B(n_30911), .C(n_27379), .Z(n_334978355
		));
	notech_ao4 i_27358208(.A(n_57566), .B(n_57657), .C(n_30723), .D(n_32227)
		, .Z(n_335478360));
	notech_or2 i_47446424(.A(n_300722032), .B(n_30719), .Z(n_335678362));
	notech_ao4 i_173844775(.A(n_30499), .B(nbus_11273[8]), .C(n_31516), .D(n_61679
		), .Z(n_335778363));
	notech_ao4 i_173744776(.A(n_30501), .B(n_33253), .C(n_5269), .D(n_30503)
		, .Z(n_335978365));
	notech_and3 i_48246423(.A(n_335778363), .B(n_335978365), .C(n_333678342)
		, .Z(n_336078366));
	notech_ao4 i_167744836(.A(n_300822033), .B(n_325325323), .C(n_262470619)
		, .D(n_315725234), .Z(n_336278367));
	notech_ao4 i_167644837(.A(n_5243), .B(n_324878257), .C(n_324778256), .D(n_33206
		), .Z(n_336478369));
	notech_nand3 i_167944834(.A(n_336278367), .B(n_336478369), .C(n_333078337
		), .Z(n_336578370));
	notech_ao4 i_167444839(.A(n_57201), .B(\nbus_11283[31] ), .C(n_57200), .D
		(\nbus_11290[31] ), .Z(n_336678371));
	notech_ao4 i_154444964(.A(n_300822033), .B(n_302878038), .C(n_262470619)
		, .D(n_303078040), .Z(n_336978374));
	notech_ao4 i_154344965(.A(n_324378252), .B(n_33206), .C(n_56783), .D(n_31539
		), .Z(n_337178376));
	notech_ao3 i_154644962(.A(n_336978374), .B(n_337178376), .C(n_332278329)
		, .Z(n_337278377));
	notech_ao4 i_154144967(.A(n_324578254), .B(\nbus_11290[31] ), .C(n_5243)
		, .D(n_324478253), .Z(n_337378378));
	notech_ao4 i_154044968(.A(n_302978039), .B(nbus_11271[31]), .C(n_324678255
		), .D(\nbus_11283[31] ), .Z(n_337478379));
	notech_ao4 i_152644982(.A(n_300822033), .B(n_124126568), .C(n_262470619)
		, .D(n_337661004), .Z(n_337678381));
	notech_ao4 i_152444984(.A(n_57012), .B(n_31539), .C(n_328660914), .D(n_31507
		), .Z(n_337878383));
	notech_and4 i_152844980(.A(n_337878383), .B(n_337678381), .C(n_331078317
		), .D(n_331378320), .Z(n_338078385));
	notech_ao4 i_152144987(.A(n_124526572), .B(\nbus_11290[31] ), .C(n_5243)
		, .D(n_124826575), .Z(n_338178386));
	notech_ao4 i_151944989(.A(n_55913), .B(n_33461), .C(n_337561003), .D(nbus_11271
		[31]), .Z(n_338378388));
	notech_and4 i_152344985(.A(n_338378388), .B(n_338178386), .C(n_330278311
		), .D(n_330578314), .Z(n_338578390));
	notech_ao4 i_151644992(.A(n_266870661), .B(n_334278348), .C(n_266970662)
		, .D(n_334078346), .Z(n_338678391));
	notech_ao4 i_151544993(.A(n_267170664), .B(n_334178347), .C(n_267470667)
		, .D(n_57394), .Z(n_338778392));
	notech_ao4 i_151344995(.A(n_58025), .B(n_31481), .C(n_300722032), .D(n_328860916
		), .Z(n_338978394));
	notech_and4 i_151844990(.A(n_338978394), .B(n_338778392), .C(n_338678391
		), .D(n_329578304), .Z(n_339178396));
	notech_ao4 i_150944998(.A(\nbus_11290[8] ), .B(n_30320), .C(n_57274), .D
		(n_33253), .Z(n_339278397));
	notech_ao4 i_150844999(.A(n_61106), .B(n_30813), .C(nbus_11273[8]), .D(n_57128
		), .Z(n_339378398));
	notech_ao4 i_150645001(.A(n_55913), .B(n_33460), .C(n_57012), .D(n_31516
		), .Z(n_339578400));
	notech_and4 i_151244996(.A(n_339578400), .B(n_339378398), .C(n_339278397
		), .D(n_328878297), .Z(n_339778402));
	notech_ao4 i_146045044(.A(n_300822033), .B(n_301522040), .C(n_262470619)
		, .D(n_298922014), .Z(n_339978403));
	notech_ao4 i_145945045(.A(n_5243), .B(n_324278251), .C(n_324178250), .D(n_33206
		), .Z(n_340178405));
	notech_nand3 i_146245042(.A(n_339978403), .B(n_340178405), .C(n_328578294
		), .Z(n_340278406));
	notech_ao4 i_145745047(.A(n_57217), .B(\nbus_11290[31] ), .C(n_58083), .D
		(n_31507), .Z(n_340378407));
	notech_ao4 i_145345051(.A(n_266870661), .B(n_333878344), .C(n_266970662)
		, .D(n_333778343), .Z(n_340678410));
	notech_ao4 i_145145053(.A(n_267170664), .B(n_333978345), .C(n_30473), .D
		(n_335678362), .Z(n_340878412));
	notech_and4 i_145545049(.A(n_340878412), .B(n_340678410), .C(n_327478283
		), .D(n_327778286), .Z(n_341078414));
	notech_ao4 i_144845056(.A(n_57243), .B(nbus_11273[8]), .C(n_57244), .D(\nbus_11290[8] 
		), .Z(n_341178415));
	notech_and3 i_144745057(.A(n_336078366), .B(n_326878277), .C(n_5774), .Z
		(n_341478418));
	notech_ao4 i_141745079(.A(n_300822033), .B(n_58100), .C(n_262470619), .D
		(n_242836107), .Z(n_341678420));
	notech_ao4 i_141545081(.A(n_60449), .B(n_31539), .C(n_385264383), .D(n_31507
		), .Z(n_341878422));
	notech_and4 i_141945077(.A(n_341878422), .B(n_341678420), .C(n_326478273
		), .D(n_326778276), .Z(n_342078424));
	notech_ao4 i_141245084(.A(n_57370), .B(\nbus_11290[31] ), .C(n_5243), .D
		(n_57325), .Z(n_342178425));
	notech_ao4 i_141145085(.A(n_32186), .B(n_33459), .C(n_248736166), .D(nbus_11271
		[31]), .Z(n_342378427));
	notech_or4 i_203358164(.A(n_32383), .B(n_60157), .C(n_32394), .D(n_61621
		), .Z(n_342578429));
	notech_nand2 i_4640030(.A(n_56927), .B(n_343778441), .Z(n_342678430));
	notech_ao4 i_4540031(.A(n_100842449), .B(n_30380), .C(\nbus_11290[2] ), 
		.D(n_57742), .Z(n_342878432));
	notech_and3 i_4740029(.A(n_346478468), .B(n_346378467), .C(n_343978443),
		 .Z(n_342978433));
	notech_and2 i_4840028(.A(n_56608), .B(n_349778500), .Z(n_343078434));
	notech_ao3 i_103539071(.A(n_436867952), .B(n_32315), .C(n_343278436), .Z
		(n_343178435));
	notech_and4 i_5140025(.A(n_346778471), .B(n_326160889), .C(n_348678489),
		 .D(n_347078474), .Z(n_343278436));
	notech_and3 i_103639070(.A(n_32310), .B(n_32223), .C(opd[2]), .Z(n_343378437
		));
	notech_and2 i_5240024(.A(n_325960887), .B(n_348578488), .Z(n_343478438)
		);
	notech_or4 i_104539061(.A(n_61912), .B(n_61901), .C(n_61885), .D(n_336360991
		), .Z(n_343778441));
	notech_nand2 i_5040026(.A(n_344378447), .B(n_349278495), .Z(n_343878442)
		);
	notech_or2 i_104839058(.A(n_344078444), .B(n_33167), .Z(n_343978443));
	notech_ao4 i_4940027(.A(n_32386), .B(n_193176989), .C(n_57047), .D(n_342578429
		), .Z(n_344078444));
	notech_or4 i_105339053(.A(n_193276990), .B(n_100842449), .C(n_2382), .D(n_2580
		), .Z(n_344378447));
	notech_ao4 i_22506(.A(n_32323), .B(n_30904), .C(n_317960807), .D(n_317860806
		), .Z(n_344478448));
	notech_nand2 i_103439072(.A(nPF), .B(n_30595), .Z(n_345678460));
	notech_nao3 i_102839078(.A(n_348378486), .B(n_342678430), .C(n_57340), .Z
		(n_345978463));
	notech_ao4 i_102939077(.A(n_57656), .B(n_30904), .C(n_343378437), .D(n_343178435
		), .Z(n_346078464));
	notech_nao3 i_104639060(.A(n_436867952), .B(n_343878442), .C(n_30309), .Z
		(n_346378467));
	notech_or4 i_104739059(.A(n_30309), .B(n_336160989), .C(n_57147), .D(n_61819
		), .Z(n_346478468));
	notech_or4 i_104039066(.A(n_2580), .B(n_326760895), .C(n_32159), .D(n_32161
		), .Z(n_346778471));
	notech_nao3 i_103939067(.A(opa[2]), .B(n_57529), .C(n_60175), .Z(n_347078474
		));
	notech_nand3 i_108839019(.A(nbus_11273[2]), .B(opa[0]), .C(opa[1]), .Z(n_347478477
		));
	notech_or2 i_108939018(.A(n_316151269), .B(nbus_11273[2]), .Z(n_347578478
		));
	notech_nand3 i_22940093(.A(n_347578478), .B(n_347478477), .C(n_27833), .Z
		(n_347878481));
	notech_xor2 i_165740069(.A(opa[4]), .B(opa[3]), .Z(n_347978482));
	notech_xor2 i_38440092(.A(n_347978482), .B(n_347878481), .Z(n_348078483)
		);
	notech_xor2 i_129140080(.A(nbus_11273[7]), .B(opa[5]), .Z(n_348178484)
		);
	notech_xor2 i_166340068(.A(nbus_11273[6]), .B(n_348178484), .Z(n_348278485
		));
	notech_xor2 i_86740094(.A(n_348278485), .B(n_348078483), .Z(n_348378486)
		);
	notech_mux2 i_208038067(.S(n_32254), .A(n_326460892), .B(n_326560893), .Z
		(n_348578488));
	notech_mux2 i_207838069(.S(n_58279), .A(n_326360891), .B(n_343478438), .Z
		(n_348678489));
	notech_ao4 i_207338073(.A(n_56766), .B(n_33167), .C(n_326260890), .D(n_58279
		), .Z(n_349278495));
	notech_ao4 i_206538080(.A(n_57656), .B(n_342978433), .C(n_342878432), .D
		(n_193176989), .Z(n_349578498));
	notech_ao3 i_206738078(.A(n_349578498), .B(n_345978463), .C(n_346078464)
		, .Z(n_349678499));
	notech_ao4 i_206938077(.A(n_57679), .B(n_342578429), .C(n_344478448), .D
		(n_30421), .Z(n_349778500));
	notech_ao4 i_206338082(.A(n_56783), .B(n_31510), .C(nbus_11273[2]), .D(n_343078434
		), .Z(n_349878501));
	notech_nao3 i_159437480(.A(n_32514), .B(n_30377), .C(n_30336), .Z(n_350078503
		));
	notech_and2 i_19437332(.A(n_376464295), .B(n_350478507), .Z(n_350178504)
		);
	notech_ao4 i_19537331(.A(n_57218), .B(n_352678529), .C(n_350778510), .D(n_350678509
		), .Z(n_350278505));
	notech_and4 i_19737329(.A(n_351778520), .B(n_351678519), .C(n_351878521)
		, .D(n_354578548), .Z(n_350378506));
	notech_or4 i_59536988(.A(tcmp), .B(n_33162), .C(n_339061018), .D(n_59312350
		), .Z(n_350478507));
	notech_ao4 i_19637330(.A(tcmp), .B(n_57566), .C(n_352678529), .D(n_32204
		), .Z(n_350678509));
	notech_and4 i_19837328(.A(n_352478527), .B(n_24735), .C(n_352378526), .D
		(n_352578528), .Z(n_350778510));
	notech_or4 i_60836975(.A(n_322660854), .B(instrc[98]), .C(instrc[97]), .D
		(instrc[99]), .Z(n_351678519));
	notech_or4 i_60936974(.A(n_79112547), .B(n_30839), .C(instrc[127]), .D(n_33162
		), .Z(n_351778520));
	notech_or2 i_61036973(.A(n_30786), .B(n_24736), .Z(n_351878521));
	notech_or4 i_60636977(.A(n_375664287), .B(instrc[105]), .C(instrc[107]),
		 .D(n_30335), .Z(n_351978522));
	notech_or4 i_60736976(.A(instrc[102]), .B(instrc[101]), .C(instrc[103]),
		 .D(n_322060848), .Z(n_352078523));
	notech_or4 i_60436979(.A(instrc[90]), .B(n_78212538), .C(n_30334), .D(n_33160
		), .Z(n_352178524));
	notech_or4 i_60536978(.A(instrc[94]), .B(n_77812534), .C(n_321960847), .D
		(n_33163), .Z(n_352278525));
	notech_or4 i_60336980(.A(n_32323), .B(n_30904), .C(n_24736), .D(n_61935)
		, .Z(n_352378526));
	notech_or4 i_60136982(.A(n_59312350), .B(n_383164362), .C(n_32646), .D(n_33162
		), .Z(n_352478527));
	notech_nand3 i_60236981(.A(n_57637), .B(n_63784), .C(n_30314), .Z(n_352578528
		));
	notech_or4 i_69637530(.A(tcmp), .B(n_61819), .C(n_339461022), .D(n_61623
		), .Z(n_352678529));
	notech_ao4 i_125336415(.A(n_350278505), .B(n_61873), .C(n_61841), .D(n_350178504
		), .Z(n_353378536));
	notech_and4 i_125836410(.A(n_352078523), .B(n_351978522), .C(n_352278525
		), .D(n_352178524), .Z(n_354578548));
	notech_ao4 i_125236416(.A(n_56704), .B(n_30664), .C(n_350078503), .D(n_350378506
		), .Z(n_355078553));
	notech_ao3 i_186837757(.A(n_19680), .B(n_30650), .C(n_1836), .Z(n_56734)
		);
	notech_ao3 i_44066191(.A(n_328660914), .B(n_328860916), .C(n_330360931),
		 .Z(n_58040));
	notech_and3 i_106666188(.A(n_83839558), .B(n_328360911), .C(n_83739557),
		 .Z(n_57439));
	notech_ao4 i_123566173(.A(n_27379), .B(n_329060918), .C(n_61845), .D(n_2805
		), .Z(n_57277));
	notech_ao4 i_123666172(.A(n_27379), .B(n_27377), .C(n_61845), .D(n_30380
		), .Z(n_57276));
	notech_or2 i_131266171(.A(n_280977820), .B(n_376064291), .Z(n_57201));
	notech_or4 i_131366170(.A(n_338661014), .B(n_285763759), .C(n_280977820)
		, .D(n_318160809), .Z(n_57200));
	notech_or4 i_1521069(.A(n_141276478), .B(n_139076456), .C(n_30278), .D(n_30279
		), .Z(n_16307));
	notech_nand2 i_1421068(.A(n_142276488), .B(n_141776483), .Z(n_16301));
	notech_and4 i_821318(.A(n_143176497), .B(n_143076496), .C(n_143676502), 
		.D(n_142976495), .Z(n_15916));
	notech_and4 i_621316(.A(n_144676512), .B(n_144576511), .C(n_145176517), 
		.D(n_144476510), .Z(n_15904));
	notech_and4 i_521315(.A(n_146176527), .B(n_146076526), .C(n_146676532), 
		.D(n_145976525), .Z(n_15898));
	notech_nand3 i_3121373(.A(n_147476540), .B(n_147376539), .C(n_147276538)
		, .Z(n_20564));
	notech_nand3 i_1521357(.A(n_148376549), .B(n_148276548), .C(n_148176547)
		, .Z(n_20468));
	notech_nand2 i_3121533(.A(n_149476560), .B(n_148976555), .Z(n_15702));
	notech_nand2 i_1021512(.A(n_150676572), .B(n_150076566), .Z(n_15576));
	notech_and4 i_821510(.A(n_151576581), .B(n_151476580), .C(n_151976585), 
		.D(n_151376579), .Z(n_15564));
	notech_and4 i_621508(.A(n_152976595), .B(n_152876594), .C(n_153376599), 
		.D(n_152776593), .Z(n_15552));
	notech_and4 i_521507(.A(n_154376609), .B(n_154276608), .C(n_154776613), 
		.D(n_154176607), .Z(n_15546));
	notech_and4 i_321505(.A(n_155776623), .B(n_155676622), .C(n_156176627), 
		.D(n_155576621), .Z(n_15534));
	notech_and4 i_221504(.A(n_157176637), .B(n_157076636), .C(n_156976635), 
		.D(n_157476640), .Z(n_15528));
	notech_and4 i_121503(.A(n_158176647), .B(n_158076646), .C(n_120176267), 
		.D(n_158476650), .Z(n_15522));
	notech_and4 i_1521837(.A(n_158676652), .B(n_158876654), .C(n_159276658),
		 .D(n_119676262), .Z(n_12728));
	notech_nand2 i_20255746(.A(sav_ecx[29]), .B(n_61873), .Z(n_160669644));
	notech_or2 i_20555743(.A(n_57326), .B(n_33197), .Z(n_160369641));
	notech_or2 i_20855740(.A(n_57369), .B(\nbus_11283[29] ), .Z(n_160069638)
		);
	notech_or4 i_3121085(.A(n_170584161), .B(n_168776753), .C(n_170076766), 
		.D(n_30286), .Z(n_16403));
	notech_nand2 i_221056(.A(n_171476780), .B(n_170976775), .Z(n_16229));
	notech_and4 i_1521517(.A(n_172876788), .B(n_172776787), .C(n_166676732),
		 .D(n_173176791), .Z(n_15606));
	notech_and4 i_821766(.A(n_174776807), .B(n_174676806), .C(n_174176801), 
		.D(n_174576805), .Z(n_15212));
	notech_and4 i_3121853(.A(n_175076810), .B(n_175276812), .C(n_175776817),
		 .D(n_164376709), .Z(n_12824));
	notech_and4 i_221824(.A(n_162876694), .B(n_176476824), .C(n_176376823), 
		.D(n_176776827), .Z(n_12650));
	notech_nand2 i_116991(.A(n_177976839), .B(n_177476834), .Z(n_11935));
	notech_ao4 i_26260788(.A(n_57566), .B(n_57637), .C(n_32210), .D(n_30316)
		, .Z(n_58218));
	notech_ao4 i_27260787(.A(n_57566), .B(n_57656), .C(n_30723), .D(n_32210)
		, .Z(n_58208));
	notech_ao3 i_38060781(.A(n_24716), .B(n_24717), .C(n_2583), .Z(n_58100)
		);
	notech_or4 i_39760778(.A(n_61823), .B(n_30309), .C(n_57637), .D(n_30473)
		, .Z(n_58083));
	notech_ao4 i_53060768(.A(n_30317), .B(n_30420), .C(n_30904), .D(n_32317)
		, .Z(n_57950));
	notech_ao4 i_113560763(.A(n_61845), .B(n_30694), .C(n_385064381), .D(n_24735
		), .Z(n_57370));
	notech_ao4 i_113660762(.A(n_61845), .B(n_335360981), .C(n_385064381), .D
		(n_383164362), .Z(n_57369));
	notech_and3 i_118060761(.A(n_379464325), .B(n_335560983), .C(n_178076840
		), .Z(n_57326));
	notech_and3 i_118160760(.A(n_379564326), .B(n_335760985), .C(n_178176841
		), .Z(n_57325));
	notech_or4 i_129560752(.A(n_32269), .B(n_58218), .C(n_32159), .D(n_256563512
		), .Z(n_57217));
	notech_or2 i_129960751(.A(n_58218), .B(n_376364294), .Z(n_57213));
	notech_or4 i_150060741(.A(n_32269), .B(n_58208), .C(n_32159), .D(n_256563512
		), .Z(n_57036));
	notech_or2 i_151060740(.A(n_376364294), .B(n_58208), .Z(n_57027));
	notech_and2 i_153060739(.A(n_204977105), .B(n_180176861), .Z(n_57010));
	notech_nand2 i_18055768(.A(sav_ecx[27]), .B(n_61873), .Z(n_159569633));
	notech_nao3 i_31763(.A(n_61885), .B(n_316260790), .C(n_316160789), .Z(n_249536174
		));
	notech_nao3 i_199060732(.A(n_32241), .B(n_30647), .C(n_385064381), .Z(n_56640
		));
	notech_or2 i_202260729(.A(n_383164362), .B(n_385064381), .Z(n_56615));
	notech_nao3 i_34670(.A(n_30314), .B(n_63784), .C(n_385064381), .Z(n_248736166
		));
	notech_nand2 i_521059(.A(n_188776945), .B(n_188176939), .Z(n_16247));
	notech_nand2 i_521347(.A(n_190176959), .B(n_189476952), .Z(n_20408));
	notech_nand2 i_221344(.A(n_191376971), .B(n_190776965), .Z(n_20390));
	notech_and4 i_121823(.A(n_191676974), .B(n_191876976), .C(n_192376981), 
		.D(n_181476874), .Z(n_12644));
	notech_or2 i_132660655(.A(n_180076860), .B(n_24736), .Z(n_242836107));
	notech_or2 i_18355765(.A(n_57326), .B(n_33195), .Z(n_159269630));
	notech_or2 i_18655762(.A(n_57369), .B(\nbus_11283[27] ), .Z(n_158969627)
		);
	notech_nand2 i_16955779(.A(sav_ecx[26]), .B(n_61871), .Z(n_158469622));
	notech_or2 i_17255776(.A(n_57326), .B(n_33198), .Z(n_158169619));
	notech_or2 i_17555773(.A(n_57369), .B(\nbus_11283[26] ), .Z(n_157869616)
		);
	notech_or2 i_203058165(.A(n_331960947), .B(n_58058), .Z(n_56608));
	notech_nand3 i_11658217(.A(instrc[118]), .B(n_30727), .C(instrc[117]), .Z
		(n_58279));
	notech_or4 i_39258204(.A(n_61823), .B(n_30309), .C(n_57637), .D(n_57616)
		, .Z(n_58088));
	notech_or4 i_42258201(.A(n_32391), .B(n_32394), .C(n_61056), .D(n_193176989
		), .Z(n_58058));
	notech_and2 i_42758200(.A(n_280177812), .B(n_196277019), .Z(n_58053));
	notech_and2 i_43658199(.A(n_58088), .B(n_196177018), .Z(n_58044));
	notech_and2 i_46158198(.A(n_280177812), .B(n_196077017), .Z(n_58019));
	notech_nor2 i_81958197(.A(n_201377069), .B(n_30300), .Z(n_57666));
	notech_and4 i_107358191(.A(n_116742608), .B(n_195677014), .C(n_280377814
		), .D(n_192776985), .Z(n_57432));
	notech_and2 i_118958187(.A(n_303178041), .B(n_195277010), .Z(n_57317));
	notech_ao4 i_122358186(.A(n_195177009), .B(n_56747), .C(n_30380), .D(n_193176989
		), .Z(n_57289));
	notech_ao4 i_126058183(.A(n_192776985), .B(n_56766), .C(n_57679), .D(n_280777818
		), .Z(n_57252));
	notech_mux2 i_166858174(.S(n_61675), .A(n_30524), .B(n_194176999), .Z(n_56896
		));
	notech_and2 i_182758170(.A(n_201777073), .B(n_60157), .Z(n_56766));
	notech_or2 i_188558169(.A(n_56766), .B(n_192776985), .Z(n_56720));
	notech_and4 i_111758188(.A(n_280377814), .B(n_195177009), .C(n_116742608
		), .D(n_195677014), .Z(n_57388));
	notech_or4 i_185258152(.A(n_2580), .B(n_32159), .C(n_32161), .D(n_193276990
		), .Z(n_56747));
	notech_and4 i_121055(.A(n_200277058), .B(n_201977075), .C(n_202177077), 
		.D(n_202677082), .Z(n_16223));
	notech_nand2 i_1021352(.A(n_203677092), .B(n_203177087), .Z(n_20438));
	notech_and4 i_121343(.A(n_204577101), .B(n_204777103), .C(n_197277029), 
		.D(n_204477100), .Z(n_20384));
	notech_ao3 i_140358177(.A(n_193076988), .B(n_194377001), .C(n_192876986)
		, .Z(n_57110));
	notech_and3 i_138058178(.A(n_201077066), .B(n_195077008), .C(n_192476982
		), .Z(n_57133));
	notech_and2 i_107958189(.A(n_342578429), .B(n_195577013), .Z(n_57426));
	notech_or4 i_163055968(.A(n_61912), .B(n_61901), .C(n_61885), .D(n_27843
		), .Z(n_56927));
	notech_and4 i_3021084(.A(n_222077272), .B(n_222577277), .C(n_220577257),
		 .D(n_222477276), .Z(n_16397));
	notech_or4 i_2921083(.A(n_216384583), .B(n_219777249), .C(n_223177283), 
		.D(n_30289), .Z(n_16391));
	notech_or4 i_2821082(.A(n_217484594), .B(n_218977241), .C(n_223877290), 
		.D(n_30290), .Z(n_16385));
	notech_or4 i_2721081(.A(n_30574), .B(n_218177233), .C(n_224577297), .D(n_30291
		), .Z(n_16379));
	notech_nand3 i_3021372(.A(n_225477306), .B(n_225377305), .C(n_225277304)
		, .Z(n_20558));
	notech_nand3 i_2921371(.A(n_226177313), .B(n_226077312), .C(n_225977311)
		, .Z(n_20552));
	notech_nand3 i_2821370(.A(n_226877320), .B(n_226777319), .C(n_226677318)
		, .Z(n_20546));
	notech_nand3 i_2721369(.A(n_227577327), .B(n_227477326), .C(n_227377325)
		, .Z(n_20540));
	notech_nand2 i_3021532(.A(n_228677338), .B(n_228177333), .Z(n_15696));
	notech_nand2 i_2921531(.A(n_229677348), .B(n_229177343), .Z(n_15690));
	notech_nand2 i_2821530(.A(n_230677358), .B(n_230177353), .Z(n_15684));
	notech_nand2 i_2721529(.A(n_231677368), .B(n_231177363), .Z(n_15678));
	notech_and4 i_3021852(.A(n_231777369), .B(n_231977371), .C(n_232477376),
		 .D(n_209477148), .Z(n_12818));
	notech_and4 i_2921851(.A(n_232577377), .B(n_232777379), .C(n_233277384),
		 .D(n_208677140), .Z(n_12812));
	notech_or4 i_2821850(.A(n_217484594), .B(n_207077125), .C(n_233677388), 
		.D(n_30292), .Z(n_12806));
	notech_and4 i_2721849(.A(n_234077392), .B(n_234277394), .C(n_234777399),
		 .D(n_206977124), .Z(n_12800));
	notech_and4 i_2917019(.A(n_235377405), .B(n_235577407), .C(n_235277404),
		 .D(n_205477110), .Z(n_12103));
	notech_ao4 i_96855012(.A(n_27798), .B(n_27843), .C(n_317960807), .D(n_317860806
		), .Z(n_156269600));
	notech_or4 i_30209(.A(instrc[113]), .B(instrc[114]), .C(n_339561023), .D
		(n_444168025), .Z(n_325325323));
	notech_mux2 i_611652(.S(n_61286), .A(n_523), .B(add_len_pc32[5]), .Z(\add_len_pc[5] 
		));
	notech_nand2 i_620676(.A(n_305378063), .B(n_304678056), .Z(n_19924));
	notech_or4 i_2021074(.A(n_261285029), .B(n_300478014), .C(n_305878068), 
		.D(n_30294), .Z(n_16337));
	notech_or4 i_1921073(.A(n_262385040), .B(n_299578006), .C(n_306578075), 
		.D(n_30295), .Z(n_16331));
	notech_or4 i_1821072(.A(n_263485051), .B(n_298777998), .C(n_307278082), 
		.D(n_30296), .Z(n_16325));
	notech_or4 i_1721071(.A(n_264585062), .B(n_297977990), .C(n_307978089), 
		.D(n_30297), .Z(n_16319));
	notech_nand3 i_2021362(.A(n_308878098), .B(n_308778097), .C(n_308678096)
		, .Z(n_20498));
	notech_nand3 i_1921361(.A(n_309578105), .B(n_309478104), .C(n_309378103)
		, .Z(n_20492));
	notech_nand3 i_1821360(.A(n_310278112), .B(n_310178111), .C(n_310078110)
		, .Z(n_20486));
	notech_nand3 i_1721359(.A(n_310978119), .B(n_310878118), .C(n_310778117)
		, .Z(n_20480));
	notech_nand2 i_421346(.A(n_312378133), .B(n_311778127), .Z(n_20402));
	notech_nand2 i_2021522(.A(n_313378143), .B(n_312878138), .Z(n_15636));
	notech_nand2 i_1921521(.A(n_314378153), .B(n_313878148), .Z(n_15630));
	notech_nand2 i_1821520(.A(n_315378163), .B(n_314878158), .Z(n_15624));
	notech_nand2 i_1721519(.A(n_316378173), .B(n_315878168), .Z(n_15618));
	notech_and4 i_421506(.A(n_317278182), .B(n_317178181), .C(n_317678186), 
		.D(n_317078180), .Z(n_15540));
	notech_and4 i_2021842(.A(n_317878188), .B(n_318078190), .C(n_318578195),
		 .D(n_286477875), .Z(n_12758));
	notech_and4 i_1921841(.A(n_318678196), .B(n_318878198), .C(n_319378203),
		 .D(n_285677867), .Z(n_12752));
	notech_and4 i_1821840(.A(n_319478204), .B(n_319678206), .C(n_320178211),
		 .D(n_284877859), .Z(n_12746));
	notech_or4 i_1721839(.A(n_264585062), .B(n_283377844), .C(n_320578215), 
		.D(n_30298), .Z(n_12740));
	notech_and4 i_2017010(.A(n_321578224), .B(n_321778226), .C(n_321478223),
		 .D(n_282677837), .Z(n_12049));
	notech_and4 i_1817008(.A(n_322478233), .B(n_322678235), .C(n_322378232),
		 .D(n_281577826), .Z(n_12037));
	notech_nao3 i_1649709(.A(n_33173), .B(n_286063762), .C(n_280277813), .Z(n_315725234
		));
	notech_and2 i_10555821(.A(n_40282), .B(n_56908), .Z(n_156169599));
	notech_and2 i_45046492(.A(n_58083), .B(n_325578264), .Z(n_58030));
	notech_and3 i_138546489(.A(n_334878354), .B(n_382164352), .C(n_334978355
		), .Z(n_57128));
	notech_nand3 i_138446488(.A(n_329760925), .B(n_334778353), .C(n_381964350
		), .Z(n_57129));
	notech_ao4 i_123846487(.A(n_335660984), .B(n_273463665), .C(n_83739557),
		 .D(n_329060918), .Z(n_57274));
	notech_ao4 i_123746486(.A(n_57679), .B(n_273363664), .C(n_83739557), .D(n_27377
		), .Z(n_57275));
	notech_and3 i_111146485(.A(n_83839558), .B(n_328360911), .C(n_27379), .Z
		(n_57394));
	notech_ao3 i_45546484(.A(n_328660914), .B(n_328760915), .C(n_330360931),
		 .Z(n_58025));
	notech_and2 i_127546475(.A(n_323078239), .B(n_325278261), .Z(n_57237));
	notech_and2 i_127446474(.A(n_323278241), .B(n_323178240), .Z(n_57238));
	notech_and4 i_111846473(.A(n_116742608), .B(n_335478360), .C(n_280977820
		), .D(n_195877016), .Z(n_57387));
	notech_and2 i_45146472(.A(n_58088), .B(n_325178260), .Z(n_58029));
	notech_and4 i_97259734(.A(n_58055), .B(n_155869596), .C(n_155669594), .D
		(n_151669554), .Z(n_156069598));
	notech_nao3 i_33345(.A(n_26063), .B(n_63794), .C(n_58218), .Z(n_301822043
		));
	notech_ao4 i_96859738(.A(n_60449), .B(n_31538), .C(n_32186), .D(n_33271)
		, .Z(n_155869596));
	notech_or2 i_33360(.A(n_57256), .B(n_30473), .Z(n_301522040));
	notech_and2 i_111246493(.A(n_57450), .B(n_58208), .Z(n_57393));
	notech_or4 i_3221086(.A(n_293885352), .B(n_332378330), .C(n_336578370), 
		.D(n_30301), .Z(n_16409));
	notech_nand3 i_3221374(.A(n_337478379), .B(n_337378378), .C(n_337278377)
		, .Z(n_20570));
	notech_nand2 i_3221534(.A(n_338578390), .B(n_338078385), .Z(n_15708));
	notech_nand2 i_921511(.A(n_339778402), .B(n_339178396), .Z(n_15570));
	notech_or4 i_3221854(.A(n_293885352), .B(n_327878287), .C(n_340278406), 
		.D(n_30302), .Z(n_12830));
	notech_and4 i_921831(.A(n_341178415), .B(n_341078414), .C(n_327178280), 
		.D(n_341478418), .Z(n_12692));
	notech_and4 i_3217022(.A(n_342178425), .B(n_342378427), .C(n_342078424),
		 .D(n_326178270), .Z(n_12121));
	notech_nao3 i_136446411(.A(n_28557), .B(n_273263663), .C(n_325078259), .Z
		(n_298922014));
	notech_and2 i_126846494(.A(n_57036), .B(n_322978238), .Z(n_57244));
	notech_and2 i_126946495(.A(n_322878237), .B(n_325678265), .Z(n_57243));
	notech_ao4 i_97059736(.A(n_58100), .B(n_5750), .C(n_57370), .D(\nbus_11290[30] 
		), .Z(n_155669594));
	notech_and4 i_97759729(.A(n_155369591), .B(n_155169589), .C(n_151969557)
		, .D(n_152269560), .Z(n_155569593));
	notech_ao4 i_97359733(.A(n_57326), .B(n_33194), .C(n_57325), .D(n_5758),
		 .Z(n_155369591));
	notech_ao4 i_97559731(.A(n_385264383), .B(n_31506), .C(n_318771158), .D(n_242836107
		), .Z(n_155169589));
	notech_and3 i_104359663(.A(n_5774), .B(n_154769585), .C(n_325860886), .Z
		(n_154969587));
	notech_ao4 i_104259664(.A(n_30590), .B(n_325060878), .C(n_25094), .D(\nbus_11290[6] 
		), .Z(n_154769585));
	notech_ao4 i_104459662(.A(n_58051), .B(n_31479), .C(n_188084307), .D(n_324960877
		), .Z(n_154569583));
	notech_nand3 i_321345(.A(n_349878501), .B(n_345678460), .C(n_349678499),
		 .Z(n_20396));
	notech_ao4 i_104559661(.A(n_57383), .B(n_325160879), .C(n_57260), .D(n_325360881
		), .Z(n_154469582));
	notech_and4 i_105659652(.A(n_154169579), .B(n_154069578), .C(n_153869576
		), .D(n_153769575), .Z(n_154369581));
	notech_ao4 i_190437728(.A(n_1850), .B(n_76712523), .C(n_30823), .D(n_350078503
		), .Z(n_56704));
	notech_ao4 i_104859658(.A(n_382664357), .B(n_100542446), .C(n_382864359)
		, .D(n_33166), .Z(n_154169579));
	notech_ao4 i_104959657(.A(n_383064361), .B(n_325260880), .C(n_56036), .D
		(n_32558), .Z(n_154069578));
	notech_ao4 i_105159655(.A(n_179284222), .B(n_325660884), .C(n_179384223)
		, .D(n_325760885), .Z(n_153869576));
	notech_ao4 i_105359654(.A(n_179484224), .B(n_325460882), .C(n_179584225)
		, .D(n_325560883), .Z(n_153769575));
	notech_or2 i_21460429(.A(n_248736166), .B(nbus_11271[30]), .Z(n_152269560
		));
	notech_or2 i_21760426(.A(n_57369), .B(\nbus_11283[30] ), .Z(n_151969557)
		);
	notech_nand2 i_22060423(.A(sav_ecx[30]), .B(n_61871), .Z(n_151669554));
	notech_nand2 i_79359912(.A(n_115942600), .B(n_32210), .Z(n_151169549));
	notech_nao3 i_156660650(.A(n_28557), .B(n_273263663), .C(n_57438), .Z(n_151069548
		));
	notech_nao3 i_153660651(.A(n_28557), .B(n_273263663), .C(n_58208), .Z(n_150969547
		));
	notech_and4 i_98462410(.A(n_150669544), .B(n_150469542), .C(n_150369541)
		, .D(n_325860886), .Z(n_150869546));
	notech_ao4 i_97962415(.A(n_25094), .B(nbus_11271[6]), .C(n_56035), .D(n_32534
		), .Z(n_150669544));
	notech_ao4 i_98162413(.A(n_23518), .B(n_325560883), .C(n_23517), .D(n_325460882
		), .Z(n_150469542));
	notech_ao4 i_98262412(.A(n_23514), .B(n_325660884), .C(n_23515), .D(n_325760885
		), .Z(n_150369541));
	notech_and4 i_99162403(.A(n_150069538), .B(n_149969537), .C(n_149769535)
		, .D(n_149669534), .Z(n_150269540));
	notech_ao4 i_98562409(.A(n_23510), .B(n_325360881), .C(n_23511), .D(n_325260880
		), .Z(n_150069538));
	notech_ao4 i_98662408(.A(n_391264443), .B(n_33166), .C(n_391164442), .D(n_100542446
		), .Z(n_149969537));
	notech_ao4 i_98862406(.A(n_23519), .B(n_324960877), .C(n_334560973), .D(n_325160879
		), .Z(n_149769535));
	notech_ao4 i_98962405(.A(n_58702), .B(n_325060878), .C(n_334460972), .D(n_31479
		), .Z(n_149669534));
	notech_and4 i_104562352(.A(n_169484150), .B(n_58055), .C(n_149269530), .D
		(n_149169529), .Z(n_149569533));
	notech_ao4 i_104062357(.A(n_24528), .B(n_33267), .C(n_24527), .D(n_33266
		), .Z(n_149269530));
	notech_and3 i_104462353(.A(n_138169419), .B(n_138069418), .C(n_149069528
		), .Z(n_149169529));
	notech_ao4 i_104262355(.A(n_60449), .B(n_31509), .C(n_24717), .D(n_334060968
		), .Z(n_149069528));
	notech_ao4 i_104662351(.A(n_61106), .B(n_30761), .C(n_381164342), .D(n_31473
		), .Z(n_148669524));
	notech_ao4 i_104762350(.A(n_380764338), .B(n_30891), .C(n_381064341), .D
		(n_33103), .Z(n_148569523));
	notech_and3 i_105262345(.A(n_139069428), .B(n_148169519), .C(n_148369521
		), .Z(n_148469522));
	notech_ao4 i_104962348(.A(n_380964340), .B(n_334360971), .C(n_30896), .D
		(n_24430), .Z(n_148369521));
	notech_ao4 i_105062347(.A(n_24421), .B(n_30916), .C(n_24733), .D(n_135369391
		), .Z(n_148169519));
	notech_and4 i_111262289(.A(n_58055), .B(n_143869476), .C(n_147769515), .D
		(n_147669514), .Z(n_148069518));
	notech_ao4 i_110662295(.A(n_24528), .B(n_33269), .C(n_24527), .D(n_33268
		), .Z(n_147769515));
	notech_and3 i_111162290(.A(n_147369511), .B(n_147569513), .C(n_139769435
		), .Z(n_147669514));
	notech_ao4 i_110862293(.A(n_60449), .B(n_31514), .C(n_24717), .D(n_337261000
		), .Z(n_147569513));
	notech_ao4 i_110962292(.A(n_381164342), .B(n_31479), .C(n_380764338), .D
		(n_325160879), .Z(n_147369511));
	notech_ao4 i_111362288(.A(n_381064341), .B(n_33166), .C(n_380964340), .D
		(n_100542446), .Z(n_147069508));
	notech_ao4 i_111462287(.A(n_24430), .B(n_324960877), .C(n_24424), .D(n_325360881
		), .Z(n_146969507));
	notech_and3 i_111962282(.A(n_140669444), .B(n_146569503), .C(n_146769505
		), .Z(n_146869506));
	notech_ao4 i_111662285(.A(n_24421), .B(n_325260880), .C(n_24431), .D(n_325660884
		), .Z(n_146769505));
	notech_ao4 i_111762284(.A(n_24429), .B(n_325460882), .C(n_24425), .D(n_325760885
		), .Z(n_146569503));
	notech_ao3 i_120062201(.A(n_169684152), .B(n_58055), .C(n_140769445), .Z
		(n_146369501));
	notech_ao4 i_120162200(.A(n_24527), .B(n_33270), .C(n_377264303), .D(n_24539
		), .Z(n_146069498));
	notech_ao4 i_120262199(.A(n_377164302), .B(n_24541), .C(n_381464345), .D
		(n_33215), .Z(n_145969497));
	notech_and4 i_121262191(.A(n_145669494), .B(n_145469492), .C(n_145369491
		), .D(n_141469452), .Z(n_145869496));
	notech_ao4 i_120562196(.A(n_385364384), .B(n_24716), .C(n_381264343), .D
		(n_31487), .Z(n_145669494));
	notech_ao4 i_120962194(.A(n_60449), .B(n_31522), .C(n_61106), .D(n_30771
		), .Z(n_145469492));
	notech_ao4 i_121062193(.A(\nbus_11290[14] ), .B(n_136169399), .C(nbus_11273
		[14]), .D(n_136069398), .Z(n_145369491));
	notech_and4 i_126162149(.A(n_144869486), .B(n_144669484), .C(n_144569483
		), .D(n_325860886), .Z(n_145069488));
	notech_ao4 i_125462154(.A(n_383264363), .B(n_61623), .C(n_151069548), .D
		(n_325360881), .Z(n_144869486));
	notech_ao4 i_125662152(.A(n_150969547), .B(n_325260880), .C(n_57027), .D
		(n_33166), .Z(n_144669484));
	notech_ao4 i_125762151(.A(n_100542446), .B(n_57036), .C(n_57438), .D(n_325160879
		), .Z(n_144569483));
	notech_and4 i_126762143(.A(n_144269480), .B(n_144069478), .C(n_143969477
		), .D(n_142869466), .Z(n_144469482));
	notech_ao4 i_126262148(.A(n_30473), .B(n_325060878), .C(n_143769475), .D
		(n_324960877), .Z(n_144269480));
	notech_ao4 i_126462146(.A(n_143469472), .B(n_325660884), .C(n_143569473)
		, .D(n_325460882), .Z(n_144069478));
	notech_ao4 i_126562145(.A(n_143669474), .B(n_325560883), .C(n_143369471)
		, .D(n_325760885), .Z(n_143969477));
	notech_ao4 i_31176(.A(n_331360941), .B(\nbus_11290[6] ), .C(n_28240), .D
		(nbus_11273[6]), .Z(n_143869476));
	notech_or2 i_4763310(.A(n_57438), .B(n_26063), .Z(n_143769475));
	notech_or4 i_8263275(.A(instrc[123]), .B(n_318060808), .C(n_143769475), 
		.D(n_32159), .Z(n_143669474));
	notech_or2 i_8163276(.A(n_143769475), .B(n_32263), .Z(n_143569473));
	notech_or2 i_8063277(.A(n_57438), .B(n_32263), .Z(n_143469472));
	notech_or4 i_8363274(.A(instrc[123]), .B(n_318060808), .C(n_57438), .D(n_32159
		), .Z(n_143369471));
	notech_or2 i_50162879(.A(n_5783), .B(n_31479), .Z(n_142869466));
	notech_or2 i_45062926(.A(n_87434558), .B(n_383164362), .Z(n_142069458)
		);
	notech_or4 i_45162925(.A(n_32275), .B(n_318160809), .C(n_87434558), .D(n_256763514
		), .Z(n_141969457));
	notech_or2 i_44462932(.A(n_97342414), .B(n_381364344), .Z(n_141469452)
		);
	notech_ao3 i_44962927(.A(n_3486), .B(n_61286), .C(n_32186), .Z(n_140769445
		));
	notech_or4 i_32963038(.A(n_24430), .B(n_61056), .C(n_30664), .D(\nbus_11290[6] 
		), .Z(n_140669444));
	notech_nand2 i_33863029(.A(sav_ecx[6]), .B(n_61871), .Z(n_139769435));
	notech_or4 i_25663105(.A(n_380764338), .B(n_24736), .C(n_61935), .D(nbus_11271
		[1]), .Z(n_139069428));
	notech_or4 i_26563097(.A(n_256763514), .B(n_32241), .C(n_256463511), .D(nbus_11273
		[1]), .Z(n_138169419));
	notech_or4 i_26463098(.A(n_256763514), .B(n_256463511), .C(n_30664), .D(\nbus_11290[1] 
		), .Z(n_138069418));
	notech_and3 i_15263207(.A(n_379564326), .B(n_56640), .C(n_141969457), .Z
		(n_136169399));
	notech_and3 i_15163208(.A(n_56615), .B(n_142069458), .C(n_379464325), .Z
		(n_136069398));
	notech_ao4 i_11463243(.A(n_60177), .B(nbus_11273[1]), .C(n_30919), .D(n_30314
		), .Z(n_135769395));
	notech_ao4 i_11563242(.A(n_60177), .B(\nbus_11290[1] ), .C(n_30920), .D(n_30314
		), .Z(n_135569393));
	notech_mux2 i_15363206(.S(n_32241), .A(n_135769395), .B(n_135569393), .Z
		(n_135369391));
	notech_ao4 i_113965040(.A(n_28240), .B(nbus_11273[6]), .C(n_26585), .D(n_30979
		), .Z(n_134869386));
	notech_ao4 i_114065039(.A(n_126126588), .B(n_32065), .C(n_125926586), .D
		(n_33261), .Z(n_134769385));
	notech_ao3 i_114565034(.A(n_134369381), .B(n_134569383), .C(n_121469252)
		, .Z(n_134669384));
	notech_ao4 i_114265037(.A(n_337261000), .B(n_26603), .C(n_26600), .D(n_31514
		), .Z(n_134569383));
	notech_ao4 i_114365036(.A(n_26277), .B(n_325560883), .C(n_26276), .D(n_325760885
		), .Z(n_134369381));
	notech_and4 i_115565024(.A(n_121969257), .B(n_133869376), .C(n_134069378
		), .D(n_133769375), .Z(n_134269380));
	notech_ao4 i_114765032(.A(n_26275), .B(n_325660884), .C(n_26271), .D(n_325260880
		), .Z(n_134069378));
	notech_ao4 i_114865031(.A(n_100542446), .B(n_332460952), .C(n_332260950)
		, .D(n_33166), .Z(n_133869376));
	notech_and3 i_115465025(.A(n_133469372), .B(n_133669374), .C(n_122469262
		), .Z(n_133769375));
	notech_ao4 i_115165028(.A(n_26278), .B(n_324960877), .C(n_332160949), .D
		(n_325160879), .Z(n_133669374));
	notech_ao4 i_115265027(.A(n_331160939), .B(\nbus_11290[6] ), .C(n_61104)
		, .D(n_30783), .Z(n_133469372));
	notech_and4 i_132364867(.A(n_143869476), .B(n_133069368), .C(n_120669244
		), .D(n_122569263), .Z(n_133269370));
	notech_ao4 i_132264868(.A(n_58040), .B(n_31479), .C(n_328760915), .D(n_337261000
		), .Z(n_133069368));
	notech_ao4 i_132464866(.A(n_57439), .B(n_325160879), .C(n_57277), .D(n_33166
		), .Z(n_132869366));
	notech_ao4 i_132564865(.A(n_57276), .B(n_100542446), .C(n_55913), .D(n_33262
		), .Z(n_132769365));
	notech_and4 i_133464856(.A(n_132469362), .B(n_132369361), .C(n_132169359
		), .D(n_132069358), .Z(n_132669364));
	notech_ao4 i_132864862(.A(n_55793), .B(n_33263), .C(n_116576231), .D(n_324960877
		), .Z(n_132469362));
	notech_ao4 i_132964861(.A(n_139276458), .B(n_325360881), .C(n_139176457)
		, .D(n_325260880), .Z(n_132369361));
	notech_ao4 i_133164859(.A(n_139376459), .B(n_325760885), .C(n_139576461)
		, .D(n_325560883), .Z(n_132169359));
	notech_ao4 i_133264858(.A(n_139676462), .B(n_325460882), .C(n_139476460)
		, .D(n_325660884), .Z(n_132069358));
	notech_and4 i_154364649(.A(n_120669244), .B(n_143869476), .C(n_131569353
		), .D(n_124069278), .Z(n_131869356));
	notech_ao4 i_154264650(.A(n_333260960), .B(n_33265), .C(n_333360961), .D
		(n_33264), .Z(n_131569353));
	notech_ao4 i_154464648(.A(n_28252), .B(n_325260880), .C(n_28251), .D(n_325360881
		), .Z(n_131369351));
	notech_ao4 i_154564647(.A(n_439667980), .B(n_100542446), .C(n_439567979)
		, .D(n_33166), .Z(n_131269350));
	notech_and4 i_155464638(.A(n_130969347), .B(n_130869346), .C(n_130669344
		), .D(n_130569343), .Z(n_131169349));
	notech_ao4 i_154864644(.A(n_439367977), .B(n_325160879), .C(n_439467978)
		, .D(n_31479), .Z(n_130969347));
	notech_ao4 i_154964643(.A(n_61104), .B(n_30840), .C(n_28260), .D(n_324960877
		), .Z(n_130869346));
	notech_ao4 i_155164641(.A(n_28255), .B(n_325560883), .C(n_28258), .D(n_325760885
		), .Z(n_130669344));
	notech_ao4 i_155264640(.A(n_28259), .B(n_325460882), .C(n_28256), .D(n_325660884
		), .Z(n_130569343));
	notech_and4 i_168564507(.A(n_130269340), .B(n_130069338), .C(n_129969337
		), .D(n_325860886), .Z(n_130469342));
	notech_ao4 i_168064512(.A(n_279977810), .B(nbus_11271[6]), .C(n_200377059
		), .D(n_325260880), .Z(n_130269340));
	notech_ao4 i_168264510(.A(n_200477060), .B(n_325360881), .C(n_323278241)
		, .D(n_100542446), .Z(n_130069338));
	notech_ao4 i_168364509(.A(n_192676984), .B(n_33166), .C(n_169676762), .D
		(n_324960877), .Z(n_129969337));
	notech_and4 i_169164501(.A(n_129669334), .B(n_129469332), .C(n_129369331
		), .D(n_126369301), .Z(n_129869336));
	notech_ao4 i_168664506(.A(n_57616), .B(n_325060878), .C(n_58044), .D(n_31479
		), .Z(n_129669334));
	notech_ao4 i_168864504(.A(n_140076466), .B(n_325660884), .C(n_139976465)
		, .D(n_325460882), .Z(n_129469332));
	notech_ao4 i_168964503(.A(n_140176467), .B(n_325760885), .C(n_139876464)
		, .D(n_325560883), .Z(n_129369331));
	notech_and4 i_178964403(.A(n_129069328), .B(n_128869326), .C(n_128769325
		), .D(n_325860886), .Z(n_129269330));
	notech_ao4 i_178464408(.A(n_29334), .B(n_325260880), .C(n_29333), .D(n_325360881
		), .Z(n_129069328));
	notech_ao4 i_178664406(.A(n_29540), .B(n_100542446), .C(n_29550), .D(n_33166
		), .Z(n_128869326));
	notech_ao4 i_178764405(.A(n_29342), .B(n_324960877), .C(n_378364314), .D
		(n_325160879), .Z(n_128769325));
	notech_and4 i_179564397(.A(n_128469322), .B(n_128269320), .C(n_128169319
		), .D(n_127669314), .Z(n_128669324));
	notech_ao4 i_179064402(.A(n_57062), .B(n_325060878), .C(n_29533), .D(\nbus_11290[6] 
		), .Z(n_128469322));
	notech_ao4 i_179264400(.A(n_29341), .B(n_325460882), .C(n_29338), .D(n_325760885
		), .Z(n_128269320));
	notech_ao4 i_179364399(.A(n_29337), .B(n_325660884), .C(n_29340), .D(n_325560883
		), .Z(n_128169319));
	notech_or2 i_91165257(.A(n_386464395), .B(n_31479), .Z(n_127669314));
	notech_or4 i_79765371(.A(n_63698), .B(n_57666), .C(n_63784), .D(nbus_11273
		[6]), .Z(n_126369301));
	notech_or2 i_65365515(.A(n_331660944), .B(n_337261000), .Z(n_124069278)
		);
	notech_nand2 i_39065771(.A(sav_esi[6]), .B(n_61871), .Z(n_122569263));
	notech_or2 i_18165976(.A(n_331460942), .B(n_31479), .Z(n_122469262));
	notech_or4 i_18665971(.A(n_332160949), .B(n_56003), .C(n_61933), .D(nbus_11271
		[6]), .Z(n_121969257));
	notech_nor2 i_19165966(.A(n_26272), .B(n_325460882), .Z(n_121469252));
	notech_nand3 i_65465514(.A(n_61104), .B(n_61623), .C(read_data[6]), .Z(n_120669244
		));
	notech_nand2 i_198286293(.A(n_1836), .B(n_19680), .Z(n_1835));
	notech_nand3 i_97686292(.A(reps[2]), .B(n_435767941), .C(n_435467938), .Z
		(n_1836));
	notech_and3 i_192137457(.A(n_33159), .B(instrc[98]), .C(n_33139), .Z(n_30864
		));
	notech_and3 i_192037458(.A(instrc[102]), .B(n_33161), .C(n_33142), .Z(n_30855
		));
	notech_or4 i_51802(.A(n_33176), .B(instrc[101]), .C(instrc[103]), .D(instrc
		[100]), .Z(n_447368057));
	notech_or4 i_51803(.A(instrc[97]), .B(n_33178), .C(instrc[99]), .D(instrc
		[96]), .Z(n_447268056));
	notech_nand2 i_1221354(.A(n_434967933), .B(n_434467928), .Z(n_447168055)
		);
	notech_ao4 i_166940130(.A(n_4448), .B(n_433867922), .C(n_431767901), .D(n_433767921
		), .Z(n_447068054));
	notech_or2 i_9413(.A(n_61816493), .B(n_3912), .Z(n_446968053));
	notech_and4 i_1216202(.A(n_429667880), .B(n_429567879), .C(n_430667890),
		 .D(n_429467878), .Z(n_446868052));
	notech_and4 i_1316203(.A(n_428067864), .B(n_427967863), .C(n_429067874),
		 .D(n_427867862), .Z(n_446768051));
	notech_or4 i_1616206(.A(n_30458), .B(n_427067854), .C(n_426567849), .D(n_426167845
		), .Z(n_446668050));
	notech_nand2 i_920839(.A(n_3906), .B(n_3902), .Z(n_446568049));
	notech_nand2 i_920743(.A(n_3897), .B(n_3889), .Z(n_446468048));
	notech_nand2 i_1220682(.A(n_3876), .B(n_3868), .Z(n_446368047));
	notech_nand2 i_1320683(.A(n_386167792), .B(n_3852), .Z(n_446268046));
	notech_nand2 i_1620686(.A(n_3846), .B(n_3840), .Z(n_446168045));
	notech_or2 i_87346440(.A(n_29888), .B(n_379364324), .Z(n_446068044));
	notech_nao3 i_86946441(.A(n_32259), .B(n_30658), .C(n_29888), .Z(n_445968043
		));
	notech_nao3 i_29323(.A(instrc[119]), .B(n_275560604), .C(n_72542166), .Z
		(n_30075));
	notech_nor2 i_29322(.A(n_72542166), .B(n_30212), .Z(n_30076));
	notech_nand3 i_29320(.A(instrc[119]), .B(n_275560604), .C(n_30428), .Z(n_30078
		));
	notech_nand3 i_28884(.A(n_339961027), .B(n_30727), .C(n_30429), .Z(n_445868042
		));
	notech_or2 i_28883(.A(n_91142352), .B(n_323660864), .Z(n_445768041));
	notech_nao3 i_28882(.A(n_339961027), .B(n_30727), .C(n_91142352), .Z(n_445668040
		));
	notech_mux2 i_1611662(.S(n_61286), .A(n_533), .B(add_len_pc32[15]), .Z(\add_len_pc[15] 
		));
	notech_mux2 i_1311659(.S(n_61286), .A(n_530), .B(add_len_pc32[12]), .Z(\add_len_pc[12] 
		));
	notech_mux2 i_1211658(.S(n_61286), .A(n_529), .B(add_len_pc32[11]), .Z(\add_len_pc[11] 
		));
	notech_and2 i_44846456(.A(n_305744491), .B(n_3619), .Z(n_4922));
	notech_nor2 i_82146457(.A(n_30077), .B(n_30483), .Z(n_72542166));
	notech_and2 i_84646458(.A(n_30196), .B(n_291167288), .Z(n_4924));
	notech_and2 i_84746459(.A(n_3606), .B(n_3620), .Z(n_72742168));
	notech_and2 i_45246468(.A(n_386864399), .B(n_3621), .Z(n_445268036));
	notech_nor2 i_82346469(.A(n_29419), .B(n_30283), .Z(n_445168035));
	notech_and2 i_84346470(.A(n_439767981), .B(n_3622), .Z(n_445068034));
	notech_and3 i_85846471(.A(n_29533), .B(n_29540), .C(n_442368007), .Z(n_444968033
		));
	notech_ao3 i_45646478(.A(n_331060938), .B(n_331660944), .C(n_333660964),
		 .Z(n_444868032));
	notech_and3 i_111546479(.A(n_28551), .B(n_330960937), .C(n_28552), .Z(n_444768031
		));
	notech_ao4 i_124346480(.A(n_57679), .B(n_273363664), .C(n_28558), .D(n_28554
		), .Z(n_444668030));
	notech_ao4 i_124446481(.A(n_335660984), .B(n_273463665), .C(n_28558), .D
		(n_323260860), .Z(n_444568029));
	notech_and3 i_138846482(.A(n_3754), .B(n_381964350), .C(n_436967953), .Z
		(n_444468028));
	notech_and3 i_138946483(.A(n_437067954), .B(n_382164352), .C(n_3755), .Z
		(n_444368027));
	notech_and3 i_84249786(.A(n_30721), .B(n_30719), .C(n_30723), .Z(n_444168025
		));
	notech_or4 i_23449789(.A(n_176660368), .B(n_32323), .C(n_30904), .D(n_61623
		), .Z(n_30695));
	notech_or4 i_23349790(.A(n_61912), .B(n_61901), .C(n_61885), .D(n_30694)
		, .Z(n_30693));
	notech_or4 i_23249791(.A(n_61892), .B(n_335660984), .C(n_61725), .D(n_32317
		), .Z(n_30697));
	notech_or4 i_23149792(.A(n_61892), .B(n_61725), .C(n_1850), .D(n_32317),
		 .Z(n_30689));
	notech_and3 i_115949764(.A(n_304744481), .B(n_30191), .C(n_3596), .Z(n_118426511
		));
	notech_and3 i_116049763(.A(n_304644480), .B(n_30196), .C(n_3595), .Z(n_118526512
		));
	notech_and3 i_115749766(.A(n_446068044), .B(n_376964300), .C(n_3598), .Z
		(n_119226519));
	notech_and3 i_115849765(.A(n_376864299), .B(n_445968043), .C(n_3597), .Z
		(n_119326520));
	notech_nao3 i_136249725(.A(instrc[117]), .B(n_286063762), .C(n_3593), .Z
		(n_444068024));
	notech_or2 i_29532(.A(n_57251), .B(n_57141), .Z(n_443968023));
	notech_nao3 i_3049699(.A(n_32259), .B(n_30658), .C(n_379064321), .Z(n_443868022
		));
	notech_or2 i_2249703(.A(n_379364324), .B(n_379064321), .Z(n_443768021)
		);
	notech_or4 i_1349712(.A(n_379064321), .B(n_33173), .C(n_30733), .D(n_61933
		), .Z(n_443668020));
	notech_nao3 i_133049726(.A(instrc[119]), .B(n_275560604), .C(n_3592), .Z
		(n_443568019));
	notech_or2 i_29212(.A(n_57251), .B(n_57117), .Z(n_443468018));
	notech_or4 i_2949700(.A(instrc[121]), .B(n_32305), .C(n_1481), .D(n_1486
		), .Z(n_443368017));
	notech_or2 i_2449701(.A(n_304344477), .B(n_1486), .Z(n_443268016));
	notech_nao3 i_1449711(.A(n_30212), .B(n_63784), .C(n_1486), .Z(n_443168015
		));
	notech_ao3 i_51666156(.A(n_265767048), .B(n_265967050), .C(n_265667047),
		 .Z(n_443068014));
	notech_nand2 i_3653038(.A(read_data[25]), .B(n_61623), .Z(n_350128600)
		);
	notech_nand2 i_3453040(.A(read_data[22]), .B(n_61623), .Z(n_350328602)
		);
	notech_or2 i_7355853(.A(n_57251), .B(n_57168), .Z(n_442968013));
	notech_nao3 i_7155855(.A(n_323660864), .B(n_63784), .C(n_323360861), .Z(n_442868012
		));
	notech_nao3 i_7055856(.A(n_339961027), .B(n_30727), .C(n_3339), .Z(n_442768011
		));
	notech_or2 i_6955857(.A(n_323360861), .B(n_337060998), .Z(n_442668010)
		);
	notech_or4 i_6855858(.A(n_338661014), .B(n_2382), .C(n_184660383), .D(n_323360861
		), .Z(n_442568009));
	notech_or4 i_12871(.A(n_32574), .B(n_32184), .C(n_61845), .D(n_340561033
		), .Z(n_442468008));
	notech_and3 i_116255971(.A(n_323860866), .B(n_442268006), .C(n_3355), .Z
		(n_117726504));
	notech_and3 i_116155972(.A(n_323960867), .B(n_442168005), .C(n_3356), .Z
		(n_117626503));
	notech_nao3 i_91355978(.A(n_29419), .B(n_32244), .C(n_286263764), .Z(n_442368007
		));
	notech_or4 i_88055979(.A(n_338661014), .B(n_2382), .C(n_184660383), .D(n_336860996
		), .Z(n_442268006));
	notech_or2 i_87155983(.A(n_337060998), .B(n_336860996), .Z(n_442168005)
		);
	notech_and4 i_53259(.A(n_442468008), .B(n_3423), .C(n_3422), .D(n_3357),
		 .Z(n_442068004));
	notech_and2 i_44460771(.A(n_382264353), .B(n_310667483), .Z(n_441968003)
		);
	notech_and2 i_125360755(.A(n_310567482), .B(n_383064361), .Z(n_441868002
		));
	notech_and2 i_126760753(.A(n_440567989), .B(n_310467481), .Z(n_441768001
		));
	notech_and2 i_138160749(.A(n_441567999), .B(n_382664357), .Z(n_441668000
		));
	notech_and2 i_1760623(.A(n_25094), .B(n_310367480), .Z(n_441567999));
	notech_nand2 i_1217578(.A(n_3338), .B(n_3331), .Z(n_441467998));
	notech_nand2 i_1317579(.A(n_3323), .B(n_3318), .Z(n_441367997));
	notech_nand2 i_1617582(.A(n_331167635), .B(n_3305), .Z(n_441267996));
	notech_nand2 i_1617006(.A(n_329867629), .B(n_329267623), .Z(n_441167995)
		);
	notech_nand2 i_321889(.A(n_328667617), .B(n_3280), .Z(n_441067994));
	notech_and4 i_1221898(.A(n_326767604), .B(n_3266), .C(n_318167544), .D(n_327067606
		), .Z(n_440967993));
	notech_nand2 i_1321899(.A(n_326067602), .B(n_3255), .Z(n_440867992));
	notech_and4 i_1621902(.A(n_324667593), .B(n_324567592), .C(n_320367565),
		 .D(n_324967596), .Z(n_440767991));
	notech_and4 i_137860750(.A(n_258463528), .B(n_116542606), .C(n_384864379
		), .D(n_382764358), .Z(n_440667990));
	notech_nao3 i_119960659(.A(n_58597), .B(n_244036119), .C(n_384764378), .Z
		(n_440567989));
	notech_and4 i_316993(.A(n_308767464), .B(n_308667463), .C(n_309767474), 
		.D(n_308567462), .Z(n_440467988));
	notech_nand2 i_1217002(.A(n_308167458), .B(n_307567452), .Z(n_440367987)
		);
	notech_nand2 i_1317003(.A(n_306967446), .B(n_306367440), .Z(n_440267986)
		);
	notech_nand2 i_321825(.A(n_305667433), .B(n_305067427), .Z(n_440167985)
		);
	notech_or4 i_1221834(.A(n_299367370), .B(n_304467421), .C(n_303967416), 
		.D(n_30509), .Z(n_440067984));
	notech_nand2 i_220832(.A(n_303567412), .B(n_303067407), .Z(n_439967983)
		);
	notech_and4 i_220736(.A(n_301867395), .B(n_302067397), .C(n_302567402), 
		.D(n_301367390), .Z(n_439867982));
	notech_nao3 i_82863399(.A(n_29419), .B(n_57472), .C(n_286263764), .Z(n_439767981
		));
	notech_ao4 i_124263381(.A(n_28551), .B(n_28554), .C(n_61846), .D(n_30380
		), .Z(n_439667980));
	notech_ao4 i_124163382(.A(n_28551), .B(n_323260860), .C(n_61846), .D(n_2805
		), .Z(n_439567979));
	notech_ao3 i_44263405(.A(n_331060938), .B(n_331760945), .C(n_333660964),
		 .Z(n_439467978));
	notech_and3 i_107063389(.A(n_28558), .B(n_330960937), .C(n_28552), .Z(n_439367977
		));
	notech_or4 i_1321835(.A(n_238466784), .B(n_30498), .C(n_290467281), .D(n_290267279
		), .Z(n_439267976));
	notech_or4 i_1621838(.A(n_239466794), .B(n_30497), .C(n_289567272), .D(n_289367270
		), .Z(n_439167975));
	notech_and4 i_321761(.A(n_288667263), .B(n_288567262), .C(n_288067257), 
		.D(n_288467261), .Z(n_439067974));
	notech_nand2 i_1221770(.A(n_287167248), .B(n_286567242), .Z(n_438967973)
		);
	notech_nand2 i_1321771(.A(n_285867235), .B(n_285267229), .Z(n_438867972)
		);
	notech_nand2 i_1621774(.A(n_284567222), .B(n_283967216), .Z(n_438767971)
		);
	notech_nand2 i_1221514(.A(n_283267209), .B(n_282667203), .Z(n_438667970)
		);
	notech_nand2 i_1321515(.A(n_282067197), .B(n_281467191), .Z(n_438567969)
		);
	notech_nand2 i_1621518(.A(n_280867185), .B(n_280267179), .Z(n_438467968)
		);
	notech_and4 i_1321355(.A(n_279367170), .B(n_279567172), .C(n_279267169),
		 .D(n_251666909), .Z(n_438367967));
	notech_and4 i_1621358(.A(n_278467161), .B(n_278667163), .C(n_278367160),
		 .D(n_252766920), .Z(n_438267966));
	notech_and4 i_321313(.A(n_277367150), .B(n_277267149), .C(n_277767154), 
		.D(n_277167148), .Z(n_438167965));
	notech_nand2 i_1221322(.A(n_276467141), .B(n_275867135), .Z(n_438067964)
		);
	notech_nand2 i_1321323(.A(n_275267129), .B(n_274667123), .Z(n_437967963)
		);
	notech_nand2 i_1621326(.A(n_274067118), .B(n_273467112), .Z(n_437867962)
		);
	notech_nand2 i_1221066(.A(n_272767106), .B(n_272167101), .Z(n_437767961)
		);
	notech_nand2 i_1321067(.A(n_271467096), .B(n_270867091), .Z(n_437667960)
		);
	notech_nand2 i_1621070(.A(n_270267087), .B(n_269767082), .Z(n_437567959)
		);
	notech_or4 i_1221002(.A(n_262367014), .B(n_30500), .C(n_269067075), .D(n_268867073
		), .Z(n_437467958));
	notech_or4 i_1321003(.A(n_263367024), .B(n_30498), .C(n_268167066), .D(n_267967064
		), .Z(n_437367957));
	notech_or4 i_1621006(.A(n_264367034), .B(n_30497), .C(n_267267057), .D(n_266867055
		), .Z(n_437267956));
	notech_nand2 i_204366167(.A(read_data[24]), .B(n_61623), .Z(n_437167955)
		);
	notech_nao3 i_121366174(.A(n_57417), .B(n_290767284), .C(n_165695997), .Z
		(n_437067954));
	notech_nao3 i_121266175(.A(n_290767284), .B(n_32544), .C(n_165695997), .Z
		(n_436967953));
	notech_or4 i_87869347(.A(instrc[121]), .B(n_32305), .C(n_1481), .D(n_30201
		), .Z(n_304644480));
	notech_or2 i_87269349(.A(n_304344477), .B(n_30201), .Z(n_304744481));
	notech_nao3 i_106040121(.A(instrc[112]), .B(n_63800), .C(n_2821), .Z(n_436867952
		));
	notech_and2 i_145237624(.A(n_33159), .B(instrc[98]), .Z(n_30865));
	notech_and2 i_67486267(.A(n_1835), .B(n_19655), .Z(n_30867));
	notech_ao3 i_187737464(.A(n_30332), .B(n_78412540), .C(instrc[96]), .Z(n_436767951
		));
	notech_or4 i_187537465(.A(n_80512561), .B(instrc[100]), .C(n_79512551), 
		.D(n_30855), .Z(n_436667950));
	notech_and2 i_110737501(.A(n_33162), .B(\opcode[0] ), .Z(n_436567949));
	notech_or4 i_2271942(.A(n_32394), .B(n_184666276), .C(n_32383), .D(n_60157
		), .Z(n_240546897));
	notech_ao3 i_071959(.A(n_178666218), .B(n_178366215), .C(n_178566217), .Z
		(n_242146913));
	notech_ao4 i_54417(.A(n_184166271), .B(n_179266224), .C(n_57147), .D(n_30800
		), .Z(n_250947001));
	notech_and3 i_11375(.A(n_61106), .B(n_61675), .C(n_179366225), .Z(n_251347005
		));
	notech_or4 i_29149(.A(n_322060848), .B(n_30618), .C(n_30343), .D(n_30550
		), .Z(n_30249));
	notech_nao3 i_28530(.A(n_61623), .B(n_32481), .C(n_32484), .Z(n_30868)
		);
	notech_nand2 i_28549(.A(instrc[101]), .B(instrc[103]), .Z(n_30849));
	notech_and2 i_145137623(.A(instrc[102]), .B(n_33161), .Z(n_436467948));
	notech_nand3 i_29150(.A(instrc[102]), .B(n_33161), .C(instrc[103]), .Z(n_30248
		));
	notech_nao3 i_6571899(.A(instrc[127]), .B(instrc[126]), .C(instrc[125]),
		 .Z(n_30266));
	notech_nand2 i_1617998(.A(n_168566129), .B(n_168466128), .Z(write_data_26
		[15]));
	notech_nand2 i_1317995(.A(n_168366127), .B(n_168266126), .Z(write_data_26
		[12]));
	notech_nand2 i_1217994(.A(n_168166125), .B(n_168066124), .Z(write_data_26
		[11]));
	notech_nand2 i_2617880(.A(n_167966123), .B(n_167866122), .Z(write_data_25
		[25]));
	notech_nao3 i_42386262(.A(reps[0]), .B(n_435667940), .C(first_rep), .Z(n_435767941
		));
	notech_xor2 i_9386261(.A(nZF), .B(reps[1]), .Z(n_435667940));
	notech_nand2 i_42086260(.A(reps[0]), .B(first_rep), .Z(n_435567939));
	notech_nand2 i_42286259(.A(n_435567939), .B(n_30313), .Z(n_435467938));
	notech_and4 i_208638061(.A(n_434767931), .B(n_434567929), .C(n_432267906
		), .D(n_432567909), .Z(n_434967933));
	notech_ao4 i_208238065(.A(n_200777063), .B(n_3753), .C(n_200677062), .D(n_3752
		), .Z(n_434767931));
	notech_ao4 i_208438063(.A(n_57133), .B(\nbus_11290[11] ), .C(n_431067894
		), .D(n_57317), .Z(n_434567929));
	notech_and4 i_209238055(.A(n_434267926), .B(n_434067924), .C(n_433967923
		), .D(n_432867912), .Z(n_434467928));
	notech_ao4 i_208738060(.A(n_58053), .B(n_31484), .C(n_56783), .D(n_31519
		), .Z(n_434267926));
	notech_ao4 i_208938058(.A(n_447068054), .B(n_57426), .C(n_57152), .D(n_433367917
		), .Z(n_434067924));
	notech_ao4 i_209038057(.A(n_430967893), .B(nbus_11273[11]), .C(n_430867892
		), .D(n_33258), .Z(n_433967923));
	notech_or2 i_212238027(.A(opbs), .B(opas), .Z(n_433867922));
	notech_nand2 i_212438025(.A(opbs), .B(opas), .Z(n_433767921));
	notech_ao4 i_212538024(.A(n_57679), .B(opa[7]), .C(opa[15]), .D(n_336360991
		), .Z(n_433667920));
	notech_or2 i_28952(.A(n_430767891), .B(n_30719), .Z(n_433367917));
	notech_or4 i_106339044(.A(n_63698), .B(n_57388), .C(n_63784), .D(nbus_11273
		[11]), .Z(n_432867912));
	notech_or4 i_106639041(.A(n_192776985), .B(n_58279), .C(n_61933), .D(n_31622
		), .Z(n_432567909));
	notech_nand2 i_106939038(.A(nOF), .B(n_30595), .Z(n_432267906));
	notech_or2 i_110139006(.A(n_27843), .B(opa[31]), .Z(n_431967903));
	notech_and2 i_2840048(.A(n_433667920), .B(n_431967903), .Z(n_431767901)
		);
	notech_ao4 i_107139036(.A(n_30528), .B(n_32317), .C(n_30317), .D(n_4443)
		, .Z(n_431367897));
	notech_and2 i_4140035(.A(n_194777005), .B(n_30421), .Z(n_431267896));
	notech_and4 i_92243368(.A(n_422767811), .B(n_422667810), .C(n_4222), .D(n_422567809
		), .Z(n_431067894));
	notech_ao3 i_4040036(.A(n_194377001), .B(n_193076988), .C(n_431367897), 
		.Z(n_430967893));
	notech_ao4 i_3940037(.A(n_57679), .B(n_431267896), .C(n_56766), .D(n_192776985
		), .Z(n_430867892));
	notech_and4 i_143446514(.A(n_3790), .B(n_3789), .C(n_3785), .D(n_3788), 
		.Z(n_430767891));
	notech_and4 i_144741898(.A(n_3967), .B(n_429967883), .C(n_430167885), .D
		(n_430567889), .Z(n_430667890));
	notech_and4 i_144241903(.A(n_446968053), .B(n_382982260), .C(n_430367887
		), .D(n_3914), .Z(n_430567889));
	notech_ao4 i_144141904(.A(n_56929), .B(\nbus_11290[27] ), .C(n_4437), .D
		(n_32168), .Z(n_430367887));
	notech_ao4 i_144341902(.A(n_60516480), .B(nbus_11273[11]), .C(n_431067894
		), .D(n_60216477), .Z(n_430167885));
	notech_ao4 i_144441901(.A(n_61116486), .B(n_33145), .C(n_60916484), .D(n_32209
		), .Z(n_429967883));
	notech_ao4 i_144841897(.A(n_61016485), .B(nbus_11271[11]), .C(n_40316278
		), .D(n_32714), .Z(n_429667880));
	notech_ao4 i_144941896(.A(n_40116276), .B(n_32876), .C(n_40216277), .D(n_31503
		), .Z(n_429567879));
	notech_and3 i_145441891(.A(n_429167875), .B(n_429367877), .C(n_3987), .Z
		(n_429467878));
	notech_ao4 i_145141894(.A(n_40616281), .B(n_32251), .C(n_443982453), .D(\nbus_11290[11] 
		), .Z(n_429367877));
	notech_ao4 i_145241893(.A(n_61716492), .B(n_32253), .C(n_4438), .D(n_31519
		), .Z(n_429167875));
	notech_and4 i_146341882(.A(n_4007), .B(n_428367867), .C(n_428567869), .D
		(n_428967873), .Z(n_429067874));
	notech_and4 i_145841887(.A(n_446968053), .B(n_382982260), .C(n_428767871
		), .D(n_398867796), .Z(n_428967873));
	notech_ao4 i_145741888(.A(n_56929), .B(\nbus_11290[28] ), .C(n_4437), .D
		(n_32169), .Z(n_428767871));
	notech_ao4 i_145941886(.A(n_60516480), .B(nbus_11273[12]), .C(n_3907), .D
		(n_60216477), .Z(n_428567869));
	notech_ao4 i_146041885(.A(n_61116486), .B(n_33149), .C(n_60916484), .D(n_32212
		), .Z(n_428367867));
	notech_ao4 i_146441881(.A(n_61016485), .B(nbus_11271[12]), .C(n_40316278
		), .D(n_32715), .Z(n_428067864));
	notech_ao4 i_146541880(.A(n_40116276), .B(n_32877), .C(n_40216277), .D(n_31504
		), .Z(n_427967863));
	notech_and3 i_147041875(.A(n_427567859), .B(n_427767861), .C(n_4052), .Z
		(n_427867862));
	notech_ao4 i_146741878(.A(n_40616281), .B(n_32248), .C(n_443982453), .D(\nbus_11290[12] 
		), .Z(n_427767861));
	notech_ao4 i_146841877(.A(n_61716492), .B(n_32255), .C(n_4438), .D(n_31520
		), .Z(n_427567859));
	notech_and4 i_150641839(.A(n_446968053), .B(n_427167855), .C(n_294388843
		), .D(n_322951208), .Z(n_427367857));
	notech_ao4 i_150541840(.A(n_25433), .B(nbus_11271[7]), .C(n_56929), .D(\nbus_11290[31] 
		), .Z(n_427167855));
	notech_nand3 i_151041835(.A(n_426767851), .B(n_426967853), .C(n_4066), .Z
		(n_427067854));
	notech_ao4 i_150741838(.A(n_4437), .B(n_32172), .C(n_60516480), .D(nbus_11273
		[15]), .Z(n_426967853));
	notech_ao4 i_150841837(.A(n_60316478), .B(n_31488), .C(n_33146), .D(n_61116486
		), .Z(n_426767851));
	notech_nand3 i_151541830(.A(n_426267846), .B(n_426467848), .C(n_4113), .Z
		(n_426567849));
	notech_ao4 i_151241833(.A(n_60916484), .B(n_32218), .C(n_61016485), .D(nbus_11271
		[15]), .Z(n_426467848));
	notech_ao4 i_151341832(.A(n_40116276), .B(n_32880), .C(n_40216277), .D(n_31507
		), .Z(n_426267846));
	notech_nao3 i_152041826(.A(n_425867842), .B(n_426067844), .C(n_4118), .Z
		(n_426167845));
	notech_ao4 i_151641829(.A(n_40616281), .B(n_32246), .C(n_4436), .D(n_32326
		), .Z(n_426067844));
	notech_ao4 i_151841828(.A(n_4438), .B(n_31523), .C(n_3909), .D(\nbus_11290[15] 
		), .Z(n_425867842));
	notech_ao4 i_195241423(.A(n_58597), .B(n_32011), .C(n_58566), .D(n_31979
		), .Z(n_425567839));
	notech_ao4 i_195341422(.A(n_30664), .B(n_31423), .C(n_57529), .D(n_33255
		), .Z(n_425467838));
	notech_and2 i_195741418(.A(n_425267836), .B(n_425167835), .Z(n_425367837
		));
	notech_ao4 i_195541420(.A(n_57449), .B(n_31587), .C(n_57435), .D(n_31947
		), .Z(n_425267836));
	notech_ao4 i_195641419(.A(n_57417), .B(n_31914), .C(n_57407), .D(n_31882
		), .Z(n_425167835));
	notech_and4 i_196641410(.A(n_424867832), .B(n_424767831), .C(n_424567829
		), .D(n_424467828), .Z(n_425067834));
	notech_ao4 i_195941416(.A(n_57517), .B(n_31850), .C(n_58555), .D(n_31818
		), .Z(n_424867832));
	notech_ao4 i_196141415(.A(n_57506), .B(n_31786), .C(n_57494), .D(n_31754
		), .Z(n_424767831));
	notech_ao4 i_196341413(.A(n_57627), .B(n_33254), .C(n_30363), .D(n_31722
		), .Z(n_424567829));
	notech_ao4 i_196441412(.A(n_57472), .B(n_31690), .C(n_57461), .D(n_31658
		), .Z(n_424467828));
	notech_ao4 i_198141395(.A(n_58597), .B(n_32008), .C(n_58566), .D(n_31976
		), .Z(n_424167825));
	notech_ao4 i_198241394(.A(n_30664), .B(n_31420), .C(n_57529), .D(n_33257
		), .Z(n_424067824));
	notech_and2 i_198641390(.A(n_423867822), .B(n_423767821), .Z(n_423967823
		));
	notech_ao4 i_198441392(.A(n_57449), .B(n_31584), .C(n_57435), .D(n_31944
		), .Z(n_423867822));
	notech_ao4 i_198541391(.A(n_57417), .B(n_31911), .C(n_57407), .D(n_31879
		), .Z(n_423767821));
	notech_and4 i_199441382(.A(n_423467818), .B(n_423367817), .C(n_423167815
		), .D(n_423067814), .Z(n_423667820));
	notech_ao4 i_198841388(.A(n_57517), .B(n_31847), .C(n_58555), .D(n_31815
		), .Z(n_423467818));
	notech_ao4 i_198941387(.A(n_57506), .B(n_31783), .C(n_57494), .D(n_31751
		), .Z(n_423367817));
	notech_ao4 i_199141385(.A(n_57627), .B(n_33256), .C(n_30363), .D(n_31719
		), .Z(n_423167815));
	notech_ao4 i_199241384(.A(n_57472), .B(n_31687), .C(n_57461), .D(n_31655
		), .Z(n_423067814));
	notech_ao4 i_214241238(.A(n_58597), .B(n_32007), .C(n_58566), .D(n_31975
		), .Z(n_422767811));
	notech_ao4 i_214341237(.A(n_30664), .B(n_31419), .C(n_57529), .D(n_33260
		), .Z(n_422667810));
	notech_and2 i_214741233(.A(n_4224), .B(n_4223), .Z(n_422567809));
	notech_ao4 i_214541235(.A(n_57449), .B(n_31583), .C(n_57435), .D(n_31943
		), .Z(n_4224));
	notech_ao4 i_214641234(.A(n_57417), .B(n_31910), .C(n_57407), .D(n_31878
		), .Z(n_4223));
	notech_and4 i_215541225(.A(n_422067808), .B(n_4218), .C(n_4214), .D(n_4212
		), .Z(n_4222));
	notech_ao4 i_214941231(.A(n_57517), .B(n_31846), .C(n_58555), .D(n_31814
		), .Z(n_422067808));
	notech_ao4 i_215041230(.A(n_57506), .B(n_31782), .C(n_57494), .D(n_31750
		), .Z(n_4218));
	notech_ao4 i_215241228(.A(n_57627), .B(n_33259), .C(n_30363), .D(n_31718
		), .Z(n_4214));
	notech_ao4 i_215341227(.A(n_57472), .B(n_31686), .C(n_57461), .D(n_31654
		), .Z(n_4212));
	notech_ao3 i_35742933(.A(imm[15]), .B(n_32243), .C(n_61816493), .Z(n_4118
		));
	notech_nao3 i_36242928(.A(nbus_136[15]), .B(n_30521), .C(n_59316468), .Z
		(n_4113));
	notech_or2 i_36742923(.A(n_3910), .B(n_60216477), .Z(n_4066));
	notech_nand2 i_30342987(.A(add_src[12]), .B(n_30416), .Z(n_4052));
	notech_or2 i_31242978(.A(n_60316478), .B(n_31485), .Z(n_4007));
	notech_or4 i_31742973(.A(n_28098), .B(n_340561033), .C(n_61623), .D(nbus_11271
		[4]), .Z(n_398867796));
	notech_nand2 i_28643004(.A(add_src[11]), .B(n_30416), .Z(n_3987));
	notech_or2 i_29542995(.A(n_60316478), .B(n_31484), .Z(n_3967));
	notech_or4 i_30042990(.A(n_28098), .B(n_340561033), .C(n_61621), .D(nbus_11271
		[3]), .Z(n_3914));
	notech_or4 i_2343254(.A(instrc[123]), .B(instrc[121]), .C(n_318160809), 
		.D(n_4432), .Z(n_3913));
	notech_and2 i_57142720(.A(n_4441), .B(n_3913), .Z(n_3912));
	notech_and4 i_92643350(.A(n_425567839), .B(n_425467838), .C(n_425067834)
		, .D(n_425367837), .Z(n_3910));
	notech_ao4 i_1843259(.A(n_26637), .B(n_27909), .C(n_25467), .D(n_61623),
		 .Z(n_3909));
	notech_and4 i_92329160(.A(n_424167825), .B(n_424067824), .C(n_423667820)
		, .D(n_423967823), .Z(n_3907));
	notech_and4 i_171544798(.A(n_3623), .B(n_336078366), .C(n_3903), .D(n_3626
		), .Z(n_3906));
	notech_ao4 i_171344800(.A(n_72742168), .B(nbus_11273[8]), .C(n_4924), .D
		(\nbus_11290[8] ), .Z(n_3903));
	notech_and4 i_172044793(.A(n_3900), .B(n_3898), .C(n_3629), .D(n_3632), 
		.Z(n_3902));
	notech_ao4 i_171644797(.A(n_267170664), .B(n_30078), .C(n_57117), .D(n_335678362
		), .Z(n_3900));
	notech_ao4 i_171844795(.A(n_266870661), .B(n_30426), .C(n_30075), .D(n_266970662
		), .Z(n_3898));
	notech_and4 i_173144782(.A(n_336078366), .B(n_3890), .C(n_3633), .D(n_3636
		), .Z(n_3897));
	notech_ao4 i_172944784(.A(n_91542356), .B(\nbus_11290[8] ), .C(n_91442355
		), .D(nbus_11273[8]), .Z(n_3890));
	notech_and4 i_173644777(.A(n_3884), .B(n_3877), .C(n_364067748), .D(n_3643
		), .Z(n_3889));
	notech_ao4 i_173244781(.A(n_267170664), .B(n_445868042), .C(n_57170), .D
		(n_335678362), .Z(n_3884));
	notech_ao4 i_173444779(.A(n_266870661), .B(n_445768041), .C(n_445668040)
		, .D(n_266970662), .Z(n_3877));
	notech_and4 i_182744686(.A(n_3873), .B(n_3870), .C(n_3869), .D(n_3646), 
		.Z(n_3876));
	notech_ao4 i_182244691(.A(n_57034), .B(n_33252), .C(n_310371085), .D(n_33258
		), .Z(n_3873));
	notech_ao4 i_182444689(.A(n_310771089), .B(n_431067894), .C(n_61104), .D
		(n_30876), .Z(n_3870));
	notech_ao4 i_182544688(.A(n_309871081), .B(n_430767891), .C(n_30326), .D
		(n_30433), .Z(n_3869));
	notech_and4 i_183344680(.A(n_3865), .B(n_3863), .C(n_3862), .D(n_365367754
		), .Z(n_3868));
	notech_ao4 i_182844685(.A(n_3750), .B(n_299422019), .C(n_265570648), .D(nbus_11273
		[11]), .Z(n_3865));
	notech_ao4 i_183044683(.A(n_299222017), .B(\nbus_11290[11] ), .C(n_265370646
		), .D(n_3751), .Z(n_3863));
	notech_ao4 i_183144682(.A(n_3752), .B(n_265070645), .C(n_3753), .D(n_264970644
		), .Z(n_3862));
	notech_and4 i_183944674(.A(n_3858), .B(n_3854), .C(n_3853), .D(n_366067761
		), .Z(n_386167792));
	notech_ao4 i_183444679(.A(n_57034), .B(n_33251), .C(n_310371085), .D(n_33250
		), .Z(n_3858));
	notech_ao4 i_183644677(.A(n_310771089), .B(n_3907), .C(n_61106), .D(n_30877
		), .Z(n_3854));
	notech_ao4 i_183744676(.A(n_309871081), .B(n_3609), .C(n_30326), .D(n_30432
		), .Z(n_3853));
	notech_and4 i_184544668(.A(n_3850), .B(n_3848), .C(n_3847), .D(n_366767768
		), .Z(n_3852));
	notech_ao4 i_184044673(.A(n_299422019), .B(n_368667786), .C(n_265570648)
		, .D(nbus_11273[12]), .Z(n_3850));
	notech_ao4 i_184244671(.A(n_299222017), .B(\nbus_11290[12] ), .C(n_265370646
		), .D(n_368767787), .Z(n_3848));
	notech_ao4 i_184344670(.A(n_265070645), .B(n_3688), .C(n_264970644), .D(n_3689
		), .Z(n_3847));
	notech_and4 i_187544638(.A(n_3844), .B(n_3842), .C(n_3841), .D(n_367467775
		), .Z(n_3846));
	notech_ao4 i_187044643(.A(n_57034), .B(n_33249), .C(n_310371085), .D(n_33248
		), .Z(n_3844));
	notech_ao4 i_187244641(.A(n_310771089), .B(n_3910), .C(n_61106), .D(n_30880
		), .Z(n_3842));
	notech_ao4 i_187344640(.A(n_309871081), .B(n_3610), .C(n_30326), .D(n_30430
		), .Z(n_3841));
	notech_and4 i_188144632(.A(n_3838), .B(n_3836), .C(n_3835), .D(n_3681), 
		.Z(n_3840));
	notech_ao4 i_187644637(.A(n_299422019), .B(n_3690), .C(n_265570648), .D(nbus_11273
		[15]), .Z(n_3838));
	notech_ao4 i_187844635(.A(n_299222017), .B(\nbus_11290[15] ), .C(n_265370646
		), .D(n_3691), .Z(n_3836));
	notech_ao4 i_187944634(.A(n_265070645), .B(n_3692), .C(n_264970644), .D(n_3693
		), .Z(n_3835));
	notech_ao4 i_197044543(.A(n_57117), .B(n_31786), .C(n_57616), .D(n_33254
		), .Z(n_3832));
	notech_ao4 i_197144542(.A(n_57141), .B(n_31754), .C(n_57147), .D(n_33255
		), .Z(n_3831));
	notech_and2 i_197544538(.A(n_3829), .B(n_3828), .Z(n_3830));
	notech_ao4 i_197344540(.A(n_57170), .B(n_31850), .C(n_30590), .D(n_32011
		), .Z(n_3829));
	notech_ao4 i_197444539(.A(n_57192), .B(n_31722), .C(n_30679), .D(n_31947
		), .Z(n_3828));
	notech_and4 i_198344530(.A(n_3825), .B(n_3824), .C(n_3822), .D(n_3821), 
		.Z(n_382767791));
	notech_ao4 i_197744536(.A(n_57064), .B(n_31690), .C(n_30473), .D(n_31818
		), .Z(n_3825));
	notech_ao4 i_197844535(.A(n_57086), .B(n_31882), .C(n_57103), .D(n_31587
		), .Z(n_3824));
	notech_ao4 i_198044533(.A(n_58702), .B(n_31979), .C(n_59100), .D(n_31914
		), .Z(n_3822));
	notech_ao4 i_198144532(.A(n_57218), .B(n_31423), .C(n_57230), .D(n_31658
		), .Z(n_3821));
	notech_ao4 i_200244511(.A(n_57122), .B(n_31783), .C(n_57616), .D(n_33256
		), .Z(n_3818));
	notech_ao4 i_200344510(.A(n_57141), .B(n_31751), .C(n_57147), .D(n_33257
		), .Z(n_3812));
	notech_and2 i_200744506(.A(n_3810), .B(n_3809), .Z(n_381167790));
	notech_ao4 i_200544508(.A(n_57170), .B(n_31847), .C(n_30590), .D(n_32008
		), .Z(n_3810));
	notech_ao4 i_200644507(.A(n_57192), .B(n_31719), .C(n_30679), .D(n_31944
		), .Z(n_3809));
	notech_and4 i_201644498(.A(n_3803), .B(n_3801), .C(n_3798), .D(n_3797), 
		.Z(n_380667789));
	notech_ao4 i_200944504(.A(n_57064), .B(n_31687), .C(n_30473), .D(n_31815
		), .Z(n_3803));
	notech_ao4 i_201044503(.A(n_57086), .B(n_31879), .C(n_57103), .D(n_31584
		), .Z(n_3801));
	notech_ao4 i_201344501(.A(n_58702), .B(n_31976), .C(n_59100), .D(n_31911
		), .Z(n_3798));
	notech_ao4 i_201444500(.A(n_57218), .B(n_31420), .C(n_57230), .D(n_31655
		), .Z(n_3797));
	notech_ao4 i_211044404(.A(n_57122), .B(n_31782), .C(n_57616), .D(n_33259
		), .Z(n_3790));
	notech_ao4 i_211144403(.A(n_57141), .B(n_31750), .C(n_57147), .D(n_33260
		), .Z(n_3789));
	notech_and2 i_211544399(.A(n_3787), .B(n_3786), .Z(n_3788));
	notech_ao4 i_211344401(.A(n_57170), .B(n_31846), .C(n_30590), .D(n_32007
		), .Z(n_3787));
	notech_ao4 i_211444400(.A(n_57195), .B(n_31718), .C(n_30679), .D(n_31943
		), .Z(n_3786));
	notech_and4 i_212344391(.A(n_3780), .B(n_3779), .C(n_3777), .D(n_3776), 
		.Z(n_3785));
	notech_ao4 i_211744397(.A(n_57064), .B(n_31686), .C(n_30473), .D(n_31814
		), .Z(n_3780));
	notech_ao4 i_211844396(.A(n_57091), .B(n_31878), .C(n_57103), .D(n_31583
		), .Z(n_3779));
	notech_ao4 i_212044394(.A(n_58702), .B(n_31975), .C(n_59100), .D(n_31910
		), .Z(n_3777));
	notech_ao4 i_212144393(.A(n_57218), .B(n_31419), .C(n_57230), .D(n_31654
		), .Z(n_3776));
	notech_nao3 i_104345414(.A(n_57417), .B(n_30910), .C(n_28551), .Z(n_3755
		));
	notech_or4 i_11986(.A(n_2382), .B(n_2383), .C(n_28551), .D(n_165695997),
		 .Z(n_3754));
	notech_nao3 i_27988(.A(n_63788), .B(opa[11]), .C(\opcode[1] ), .Z(n_3753
		));
	notech_nand2 i_27989(.A(n_63788), .B(opc[11]), .Z(n_3752));
	notech_nand2 i_27991(.A(n_63788), .B(opc_10[11]), .Z(n_3751));
	notech_nao3 i_28011(.A(n_61933), .B(opa[11]), .C(n_63712), .Z(n_3750));
	notech_nao3 i_27807(.A(n_63788), .B(opa[15]), .C(n_63712), .Z(n_3693));
	notech_nand2 i_27810(.A(n_63788), .B(opc[15]), .Z(n_3692));
	notech_nand2 i_27813(.A(n_63788), .B(opc_10[15]), .Z(n_3691));
	notech_nao3 i_27836(.A(n_61933), .B(opa[15]), .C(n_63712), .Z(n_3690));
	notech_nao3 i_27944(.A(n_63796), .B(opa[12]), .C(n_63712), .Z(n_3689));
	notech_nand2 i_27945(.A(n_63796), .B(opc[12]), .Z(n_3688));
	notech_nand2 i_27947(.A(n_63796), .B(opc_10[12]), .Z(n_368767787));
	notech_nao3 i_27967(.A(n_61933), .B(opa[12]), .C(n_63712), .Z(n_368667786
		));
	notech_nao3 i_29980(.A(instrc[117]), .B(n_290663806), .C(n_445168035), .Z
		(n_29418));
	notech_nor2 i_29981(.A(n_445168035), .B(n_29557), .Z(n_29417));
	notech_nand3 i_29982(.A(n_290663806), .B(instrc[117]), .C(n_30282), .Z(n_29416
		));
	notech_or2 i_31030(.A(n_444768031), .B(n_28555), .Z(n_28368));
	notech_or2 i_31031(.A(n_444768031), .B(n_30441), .Z(n_28367));
	notech_or2 i_31033(.A(n_28558), .B(n_30441), .Z(n_28365));
	notech_nand2 i_84145603(.A(opd[15]), .B(n_300322028), .Z(n_3681));
	notech_nao3 i_85545596(.A(n_19655), .B(read_data[15]), .C(n_60449), .Z(n_367467775
		));
	notech_nand2 i_79645643(.A(n_300322028), .B(opd[12]), .Z(n_366767768));
	notech_nao3 i_80345636(.A(n_19655), .B(read_data[12]), .C(n_60449), .Z(n_366067761
		));
	notech_nand2 i_78245657(.A(opd[11]), .B(n_300322028), .Z(n_365367754));
	notech_nao3 i_78945650(.A(n_19655), .B(read_data[11]), .C(n_60449), .Z(n_3646
		));
	notech_or4 i_65945778(.A(n_63718), .B(n_91142352), .C(n_63794), .D(nbus_11273
		[8]), .Z(n_3643));
	notech_or2 i_66245775(.A(n_90742348), .B(n_31481), .Z(n_364067748));
	notech_nao3 i_66545772(.A(n_30429), .B(\opa_12[8] ), .C(n_337060998), .Z
		(n_3636));
	notech_or2 i_66645771(.A(n_442268006), .B(n_5269), .Z(n_3633));
	notech_or4 i_64145796(.A(n_63718), .B(n_72542166), .C(n_63758), .D(nbus_11273
		[8]), .Z(n_3632));
	notech_or2 i_64445793(.A(n_4922), .B(n_31481), .Z(n_3629));
	notech_nao3 i_64745790(.A(n_30428), .B(\opa_12[8] ), .C(n_304344477), .Z
		(n_3626));
	notech_or4 i_64845789(.A(n_1481), .B(n_30201), .C(n_5269), .D(n_57506), 
		.Z(n_3623));
	notech_nao3 i_103845418(.A(n_57472), .B(n_30283), .C(n_286263764), .Z(n_3622
		));
	notech_nand2 i_103745419(.A(n_115442595), .B(n_32211), .Z(n_3621));
	notech_nao3 i_103045426(.A(n_57506), .B(n_30483), .C(n_1481), .Z(n_3620)
		);
	notech_nand2 i_102945427(.A(n_115442595), .B(n_125342694), .Z(n_3619));
	notech_nao3 i_102845428(.A(n_57517), .B(n_30484), .C(n_184660383), .Z(n_3618
		));
	notech_nand2 i_102745429(.A(n_115442595), .B(n_32220), .Z(n_3617));
	notech_and4 i_143829657(.A(n_3832), .B(n_3831), .C(n_382767791), .D(n_3830
		), .Z(n_3610));
	notech_and4 i_143546445(.A(n_3818), .B(n_3812), .C(n_380667789), .D(n_381167790
		), .Z(n_3609));
	notech_and2 i_84946455(.A(n_292067297), .B(n_323860866), .Z(n_91542356)
		);
	notech_and2 i_84846454(.A(n_3607), .B(n_3618), .Z(n_91442355));
	notech_and2 i_44746452(.A(n_327960907), .B(n_3617), .Z(n_90742348));
	notech_nor2 i_82446453(.A(n_3608), .B(n_30484), .Z(n_91142352));
	notech_nand3 i_82069352(.A(n_57544), .B(n_323360861), .C(n_184360381), .Z
		(n_3608));
	notech_nao3 i_83163396(.A(n_3608), .B(n_57517), .C(n_184660383), .Z(n_3607
		));
	notech_nao3 i_83063397(.A(n_30077), .B(n_57506), .C(n_1481), .Z(n_3606)
		);
	notech_or2 i_119348588(.A(n_379364324), .B(n_29887), .Z(n_3598));
	notech_nao3 i_119248589(.A(n_32259), .B(n_30658), .C(n_29887), .Z(n_3597
		));
	notech_or2 i_119148590(.A(n_304344477), .B(n_30200), .Z(n_3596));
	notech_or4 i_119048591(.A(instrc[121]), .B(n_32305), .C(n_1481), .D(n_30200
		), .Z(n_3595));
	notech_nand3 i_29520(.A(instrc[117]), .B(n_286063762), .C(n_63758), .Z(n_3594
		));
	notech_and4 i_117548598(.A(n_234763344), .B(n_57544), .C(n_29888), .D(n_379164322
		), .Z(n_3593));
	notech_and4 i_117448599(.A(n_57544), .B(n_1484), .C(n_30201), .D(n_305844492
		), .Z(n_3592));
	notech_and3 i_161651474(.A(n_358267744), .B(n_358167743), .C(n_3589), .Z
		(n_3590));
	notech_and4 i_161551475(.A(n_3587), .B(n_3586), .C(n_358467746), .D(n_352767691
		), .Z(n_3589));
	notech_ao4 i_160951481(.A(n_126826595), .B(\nbus_11290[24] ), .C(n_126726594
		), .D(\nbus_11283[24] ), .Z(n_3587));
	notech_ao4 i_160851482(.A(n_337761005), .B(nbus_11271[24]), .C(n_125926586
		), .D(n_33247), .Z(n_3586));
	notech_ao4 i_160751483(.A(n_126126588), .B(n_32083), .C(n_26585), .D(n_31016
		), .Z(n_358467746));
	notech_ao4 i_161151479(.A(n_337861006), .B(n_31500), .C(n_26600), .D(n_31532
		), .Z(n_358267744));
	notech_ao4 i_161051480(.A(n_126926596), .B(n_33171), .C(n_106826395), .D
		(n_127026597), .Z(n_358167743));
	notech_nand3 i_113451953(.A(n_357667738), .B(n_357567737), .C(n_357467736
		), .Z(n_357867740));
	notech_ao4 i_112651959(.A(n_122726554), .B(\nbus_11283[24] ), .C(n_337361001
		), .D(nbus_11271[24]), .Z(n_357667738));
	notech_ao4 i_112551960(.A(n_333360961), .B(n_33246), .C(n_333260960), .D
		(n_33245), .Z(n_357567737));
	notech_ao4 i_113151956(.A(n_61106), .B(n_30856), .C(n_57012), .D(n_31532
		), .Z(n_357467736));
	notech_nand2 i_113351954(.A(n_357267734), .B(n_357167733), .Z(n_357367735
		));
	notech_ao4 i_112851957(.A(n_31500), .B(n_331060938), .C(n_122826555), .D
		(n_33171), .Z(n_357267734));
	notech_ao4 i_112751958(.A(n_106826395), .B(n_122926556), .C(n_122626553)
		, .D(\nbus_11290[24] ), .Z(n_357167733));
	notech_nand3 i_110951976(.A(n_356567728), .B(n_356367727), .C(n_356267726
		), .Z(n_356867730));
	notech_ao4 i_110351982(.A(n_122726554), .B(\nbus_11283[25] ), .C(n_337361001
		), .D(nbus_11271[25]), .Z(n_356567728));
	notech_ao4 i_110251983(.A(n_333360961), .B(n_33244), .C(n_333260960), .D
		(n_33243), .Z(n_356367727));
	notech_ao4 i_110651979(.A(n_61106), .B(n_30857), .C(n_57012), .D(n_31533
		), .Z(n_356267726));
	notech_nand2 i_110851977(.A(n_356067724), .B(n_355967723), .Z(n_356167725
		));
	notech_ao4 i_110551980(.A(n_331060938), .B(n_31501), .C(n_122826555), .D
		(n_33172), .Z(n_356067724));
	notech_ao4 i_110451981(.A(n_101026337), .B(n_122926556), .C(n_122626553)
		, .D(\nbus_11290[25] ), .Z(n_355967723));
	notech_and4 i_76352318(.A(n_355467718), .B(n_355367717), .C(n_355267716)
		, .D(n_354467708), .Z(n_355767721));
	notech_ao4 i_75952322(.A(n_59464), .B(n_119326520), .C(n_443868022), .D(n_58875
		), .Z(n_355467718));
	notech_ao4 i_75852323(.A(n_443768021), .B(n_58411), .C(n_443668020), .D(n_60537
		), .Z(n_355367717));
	notech_ao4 i_76052321(.A(n_379264323), .B(n_31496), .C(n_119226519), .D(n_33284
		), .Z(n_355267716));
	notech_nand3 i_63452447(.A(n_354767711), .B(n_354667710), .C(n_354567709
		), .Z(n_354967713));
	notech_ao4 i_63152450(.A(n_101026337), .B(n_118526512), .C(n_443368017),
		 .D(n_58920), .Z(n_354767711));
	notech_ao4 i_63052451(.A(n_443268016), .B(\nbus_11283[25] ), .C(n_443168015
		), .D(nbus_11271[25]), .Z(n_354667710));
	notech_ao4 i_63252449(.A(n_305744491), .B(n_31501), .C(n_118426511), .D(n_33172
		), .Z(n_354567709));
	notech_and3 i_51453073(.A(n_350328602), .B(n_354267706), .C(n_354167705)
		, .Z(n_354467708));
	notech_ao4 i_55652524(.A(n_30693), .B(n_58875), .C(n_30695), .D(n_58411)
		, .Z(n_354267706));
	notech_ao4 i_55752523(.A(n_30697), .B(n_33284), .C(n_59464), .D(n_30689)
		, .Z(n_354167705));
	notech_nand2 i_52552555(.A(n_353767701), .B(n_353667700), .Z(n_353867702
		));
	notech_ao4 i_52352557(.A(n_117626503), .B(n_33171), .C(n_106826395), .D(n_117726504
		), .Z(n_353767701));
	notech_ao4 i_52252558(.A(n_442568009), .B(\nbus_11290[24] ), .C(n_442668010
		), .D(\nbus_11283[24] ), .Z(n_353667700));
	notech_nao3 i_52452556(.A(n_443068014), .B(n_3434), .C(n_3440), .Z(n_353567699
		));
	notech_nand3 i_51753071(.A(n_350128600), .B(n_353167695), .C(n_353067694
		), .Z(n_353367697));
	notech_ao4 i_48952586(.A(n_30693), .B(n_58920), .C(n_30695), .D(n_58438)
		, .Z(n_353167695));
	notech_ao4 i_49052585(.A(n_30697), .B(n_33172), .C(n_101026337), .D(n_30689
		), .Z(n_353067694));
	notech_nand3 i_2521783(.A(n_352867692), .B(n_3590), .C(n_351667680), .Z(n_352967693
		));
	notech_nao3 i_160651484(.A(n_63796), .B(opc_10[24]), .C(n_337961007), .Z
		(n_352867692));
	notech_nand2 i_160451486(.A(sav_esp[24]), .B(n_61871), .Z(n_352767691)
		);
	notech_or2 i_160551485(.A(n_126226589), .B(n_364628688), .Z(n_351667680)
		);
	notech_or4 i_2521335(.A(n_351467678), .B(n_357867740), .C(n_357367735), 
		.D(n_350267667), .Z(n_351567679));
	notech_ao3 i_112451961(.A(n_63796), .B(opc_10[24]), .C(n_337461002), .Z(n_351467678
		));
	notech_nor2 i_112351962(.A(n_122226549), .B(n_364628688), .Z(n_350267667
		));
	notech_or4 i_2621336(.A(n_349867665), .B(n_356867730), .C(n_356167725), 
		.D(n_348667654), .Z(n_350167666));
	notech_ao3 i_110151984(.A(n_63796), .B(opc_10[25]), .C(n_337461002), .Z(n_349867665
		));
	notech_nor2 i_110051985(.A(n_122226549), .B(n_363350926), .Z(n_348667654
		));
	notech_nand3 i_2320981(.A(n_355767721), .B(n_347567645), .C(n_348267652)
		, .Z(n_348567653));
	notech_nao3 i_75752324(.A(opc_10[22]), .B(n_63758), .C(n_444068024), .Z(n_348267652
		));
	notech_or4 i_75652325(.A(n_340461032), .B(n_339561023), .C(n_57256), .D(n_3464
		), .Z(n_347567645));
	notech_or4 i_2620856(.A(n_353367697), .B(n_354967713), .C(n_347267643), 
		.D(n_3449), .Z(n_347367644));
	notech_ao3 i_62952452(.A(n_63796), .B(opc_10[25]), .C(n_443568019), .Z(n_347267643
		));
	notech_nor2 i_62852453(.A(n_363350926), .B(n_443468018), .Z(n_3449));
	notech_or4 i_2520759(.A(n_353867702), .B(n_353567699), .C(n_3441), .D(n_3433
		), .Z(n_3442));
	notech_ao3 i_52052560(.A(n_63796), .B(opc_10[24]), .C(n_442768011), .Z(n_3441
		));
	notech_ao3 i_51852562(.A(n_57397), .B(opd[24]), .C(n_57170), .Z(n_3440)
		);
	notech_or2 i_50852567(.A(n_442868012), .B(nbus_11271[24]), .Z(n_3434));
	notech_nor2 i_51952561(.A(n_364628688), .B(n_442968013), .Z(n_3433));
	notech_ao4 i_186354134(.A(n_114845640), .B(n_57064), .C(n_3410), .D(n_217373541
		), .Z(n_3423));
	notech_and4 i_186854129(.A(n_3365), .B(n_3421), .C(n_3366), .D(n_3364), 
		.Z(n_3422));
	notech_ao4 i_186554132(.A(n_3343), .B(n_350078503), .C(n_3342), .D(n_3341
		), .Z(n_3421));
	notech_ao4 i_187054127(.A(n_29232), .B(n_3347), .C(n_30743), .D(n_3346),
		 .Z(n_3419));
	notech_ao4 i_187254125(.A(n_3345), .B(n_156594048), .C(n_30786), .D(n_30269
		), .Z(n_3417));
	notech_and2 i_187354124(.A(n_3400), .B(n_3399), .Z(n_3416));
	notech_ao4 i_5855868(.A(n_57637), .B(n_2810), .C(n_32211), .D(n_30798), 
		.Z(n_3410));
	notech_or4 i_188054117(.A(instrc[124]), .B(n_32646), .C(n_30552), .D(n_33153
		), .Z(n_3409));
	notech_nao3 i_188754110(.A(n_32514), .B(n_30377), .C(n_349971384), .Z(n_3404
		));
	notech_nand3 i_7171893(.A(instrc[125]), .B(n_33175), .C(instrc[127]), .Z
		(n_3402));
	notech_nand2 i_101054974(.A(n_321860846), .B(n_57064), .Z(n_3401));
	notech_nand2 i_30162(.A(instrc[99]), .B(n_33178), .Z(n_29236));
	notech_or4 i_101254972(.A(n_436667950), .B(instrc[102]), .C(n_33142), .D
		(n_33161), .Z(n_3400));
	notech_or4 i_101154973(.A(instrc[98]), .B(n_30449), .C(n_33139), .D(n_33159
		), .Z(n_3399));
	notech_or4 i_101954967(.A(n_30552), .B(n_30839), .C(n_33153), .D(instrc[
		124]), .Z(n_3394));
	notech_nao3 i_100354981(.A(instrc[117]), .B(n_290663806), .C(n_3340), .Z
		(n_3366));
	notech_or4 i_100254982(.A(n_339061018), .B(n_76712523), .C(instrc[124]),
		 .D(n_3402), .Z(n_3365));
	notech_or4 i_100154983(.A(n_349671381), .B(n_33242), .C(n_30383), .D(n_3404
		), .Z(n_3364));
	notech_or2 i_100854976(.A(n_57472), .B(n_56704), .Z(n_3357));
	notech_or2 i_98754996(.A(n_337060998), .B(n_337160999), .Z(n_3356));
	notech_or4 i_98654997(.A(n_338661014), .B(n_2382), .C(n_184660383), .D(n_337160999
		), .Z(n_3355));
	notech_nand3 i_2971935(.A(instrc[105]), .B(instrc[107]), .C(n_30829), .Z
		(n_3347));
	notech_nand3 i_5871906(.A(instrc[89]), .B(instrc[91]), .C(n_322260850), 
		.Z(n_3346));
	notech_nao3 i_4971915(.A(instrc[93]), .B(instrc[95]), .C(n_321960847), .Z
		(n_3345));
	notech_and4 i_9455832(.A(n_3394), .B(n_3419), .C(n_3417), .D(n_3416), .Z
		(n_3343));
	notech_and4 i_9355833(.A(n_322760855), .B(n_322860856), .C(n_3410), .D(n_3401
		), .Z(n_3342));
	notech_ao4 i_2955897(.A(n_286263764), .B(n_57472), .C(n_386964400), .D(n_3409
		), .Z(n_3341));
	notech_ao4 i_9255834(.A(n_322560853), .B(n_32211), .C(n_339261020), .D(n_61933
		), .Z(n_3340));
	notech_and4 i_5055876(.A(n_57544), .B(n_184360381), .C(n_336860996), .D(n_328060908
		), .Z(n_3339));
	notech_and4 i_86759838(.A(n_3336), .B(n_3332), .C(n_311167488), .D(n_310067477
		), .Z(n_3338));
	notech_ao4 i_86359842(.A(n_25094), .B(nbus_11271[11]), .C(n_3751), .D(n_23611
		), .Z(n_3336));
	notech_ao4 i_86559840(.A(n_3753), .B(n_23614), .C(n_3752), .D(n_23613), 
		.Z(n_3332));
	notech_and4 i_87359832(.A(n_3329), .B(n_3327), .C(n_3325), .D(n_311467491
		), .Z(n_3331));
	notech_ao4 i_86859837(.A(n_386264393), .B(n_31484), .C(n_23747), .D(n_33258
		), .Z(n_3329));
	notech_ao4 i_87059835(.A(n_431067894), .B(n_23750), .C(\nbus_11290[11] )
		, .D(n_386164392), .Z(n_3327));
	notech_ao4 i_87159834(.A(n_386064391), .B(nbus_11273[11]), .C(n_56035), 
		.D(n_32540), .Z(n_3325));
	notech_and4 i_87859827(.A(n_3321), .B(n_3319), .C(n_312467498), .D(n_310167478
		), .Z(n_3323));
	notech_ao4 i_87459831(.A(n_25094), .B(nbus_11271[12]), .C(n_368767787), 
		.D(n_23611), .Z(n_3321));
	notech_ao4 i_87659829(.A(n_3689), .B(n_23614), .C(n_3688), .D(n_23613), 
		.Z(n_3319));
	notech_and4 i_88459821(.A(n_3316), .B(n_331467636), .C(n_3313), .D(n_3128
		), .Z(n_3318));
	notech_ao4 i_87959826(.A(n_23747), .B(n_33250), .C(n_3907), .D(n_23750),
		 .Z(n_3316));
	notech_ao4 i_88159824(.A(n_386164392), .B(\nbus_11290[12] ), .C(n_386064391
		), .D(nbus_11273[12]), .Z(n_331467636));
	notech_ao4 i_88259823(.A(n_56035), .B(n_32541), .C(n_58702), .D(n_309867475
		), .Z(n_3313));
	notech_and4 i_91159794(.A(n_330867634), .B(n_330667633), .C(n_313867507)
		, .D(n_310267479), .Z(n_331167635));
	notech_ao4 i_90759798(.A(n_25094), .B(nbus_11271[15]), .C(n_3691), .D(n_23611
		), .Z(n_330867634));
	notech_ao4 i_90959796(.A(n_3693), .B(n_23614), .C(n_3692), .D(n_23613), 
		.Z(n_330667633));
	notech_and4 i_91759788(.A(n_3302), .B(n_330067631), .C(n_329967630), .D(n_314167510
		), .Z(n_3305));
	notech_ao4 i_91259793(.A(n_23747), .B(n_33248), .C(n_3910), .D(n_23750),
		 .Z(n_3302));
	notech_ao4 i_91459791(.A(n_386164392), .B(\nbus_11290[15] ), .C(n_386064391
		), .D(nbus_11273[15]), .Z(n_330067631));
	notech_ao4 i_91559790(.A(n_56035), .B(n_32545), .C(n_58702), .D(n_309967476
		), .Z(n_329967630));
	notech_and4 i_92359782(.A(n_329667627), .B(n_329467625), .C(n_329367624)
		, .D(n_314867517), .Z(n_329867629));
	notech_ao4 i_91859787(.A(n_61106), .B(n_30772), .C(n_381264343), .D(n_31488
		), .Z(n_329667627));
	notech_ao4 i_92059785(.A(n_3690), .B(n_381564346), .C(n_3910), .D(n_381364344
		), .Z(n_329467625));
	notech_ao4 i_92159784(.A(n_381464345), .B(n_33248), .C(n_381664347), .D(\nbus_11290[15] 
		), .Z(n_329367624));
	notech_and4 i_92959776(.A(n_329067621), .B(n_328867619), .C(n_328767618)
		, .D(n_315667524), .Z(n_329267623));
	notech_ao4 i_92459781(.A(n_3693), .B(n_24542), .C(n_3692), .D(n_24541), 
		.Z(n_329067621));
	notech_ao4 i_92659779(.A(n_3691), .B(n_24539), .C(n_24528), .D(n_33241),
		 .Z(n_328867619));
	notech_ao4 i_92759778(.A(n_24527), .B(n_33240), .C(n_3610), .D(n_24716),
		 .Z(n_328767618));
	notech_and4 i_100559701(.A(n_328467615), .B(n_3282), .C(n_328167613), .D
		(n_326860896), .Z(n_328667617));
	notech_ao4 i_100059706(.A(n_25094), .B(\nbus_11290[2] ), .C(n_58051), .D
		(n_31474), .Z(n_328467615));
	notech_ao4 i_100259704(.A(n_325960887), .B(n_188084307), .C(n_326160889)
		, .D(n_57383), .Z(n_3282));
	notech_ao4 i_100359703(.A(n_326360891), .B(n_57260), .C(n_382664357), .D
		(n_100842449), .Z(n_328167613));
	notech_and4 i_101259694(.A(n_327867611), .B(n_327767610), .C(n_327367608
		), .D(n_3272), .Z(n_3280));
	notech_ao4 i_100659700(.A(n_382864359), .B(n_33167), .C(n_326260890), .D
		(n_383064361), .Z(n_327867611));
	notech_ao4 i_100759699(.A(n_56035), .B(n_32554), .C(n_30590), .D(n_326060888
		), .Z(n_327767610));
	notech_ao4 i_100959697(.A(n_326660894), .B(n_179284222), .C(n_179384223)
		, .D(n_326760895), .Z(n_327367608));
	notech_ao4 i_101059696(.A(n_326460892), .B(n_179484224), .C(n_326560893)
		, .D(n_179584225), .Z(n_3272));
	notech_and3 i_110059615(.A(n_5774), .B(n_317567542), .C(n_310067477), .Z
		(n_327067606));
	notech_ao4 i_110159614(.A(n_441868002), .B(n_3752), .C(n_3753), .D(n_4533
		), .Z(n_326767604));
	notech_and4 i_111159606(.A(n_3264), .B(n_3262), .C(n_3261), .D(n_318467547
		), .Z(n_3266));
	notech_ao4 i_110459611(.A(n_440667990), .B(n_3750), .C(n_441668000), .D(\nbus_11290[11] 
		), .Z(n_3264));
	notech_ao4 i_110759609(.A(n_56036), .B(n_32563), .C(n_385464385), .D(n_3751
		), .Z(n_3262));
	notech_ao4 i_110859608(.A(n_385664387), .B(n_33258), .C(n_385864389), .D
		(n_431067894), .Z(n_3261));
	notech_and4 i_111659601(.A(n_3258), .B(n_3256), .C(n_310167478), .D(n_319367556
		), .Z(n_326067602));
	notech_ao4 i_111259605(.A(n_31485), .B(n_441968003), .C(n_3688), .D(n_441868002
		), .Z(n_3258));
	notech_ao4 i_111459603(.A(n_441768001), .B(nbus_11273[12]), .C(n_440667990
		), .D(n_368667786), .Z(n_3256));
	notech_and4 i_112159596(.A(n_3253), .B(n_325167598), .C(n_319667559), .D
		(n_319967562), .Z(n_3255));
	notech_ao4 i_111759600(.A(n_56036), .B(n_32564), .C(n_30590), .D(n_309867475
		), .Z(n_3253));
	notech_ao4 i_111959598(.A(n_385664387), .B(n_33250), .C(n_385864389), .D
		(n_3907), .Z(n_325167598));
	notech_ao3 i_114959572(.A(n_320067563), .B(n_310267479), .C(n_335060978)
		, .Z(n_324967596));
	notech_ao4 i_115059571(.A(n_3693), .B(n_4533), .C(n_441768001), .D(nbus_11273
		[15]), .Z(n_324667593));
	notech_and4 i_115859563(.A(n_324367590), .B(n_324167588), .C(n_324067587
		), .D(n_320767568), .Z(n_324567592));
	notech_ao4 i_115359568(.A(n_441668000), .B(\nbus_11290[15] ), .C(n_56036
		), .D(n_32567), .Z(n_324367590));
	notech_ao4 i_115559566(.A(n_30590), .B(n_309967476), .C(n_385464385), .D
		(n_3691), .Z(n_324167588));
	notech_ao4 i_115659565(.A(n_385664387), .B(n_33248), .C(n_385864389), .D
		(n_3910), .Z(n_324067587));
	notech_ao4 i_156259197(.A(n_431067894), .B(n_30503), .C(n_30496), .D(\nbus_11290[11] 
		), .Z(n_3239));
	notech_ao4 i_156359196(.A(n_30499), .B(nbus_11273[11]), .C(n_30501), .D(n_33258
		), .Z(n_323767585));
	notech_ao4 i_156559194(.A(n_3907), .B(n_30503), .C(n_30496), .D(\nbus_11290[12] 
		), .Z(n_3236));
	notech_ao4 i_156759193(.A(n_30499), .B(nbus_11273[12]), .C(n_30501), .D(n_33250
		), .Z(n_3234));
	notech_ao4 i_157559185(.A(n_3910), .B(n_30503), .C(n_30496), .D(\nbus_11290[15] 
		), .Z(n_323367583));
	notech_ao4 i_157659184(.A(n_30499), .B(nbus_11273[15]), .C(n_30501), .D(n_33248
		), .Z(n_323167581));
	notech_or2 i_126160754(.A(n_440667990), .B(n_25121), .Z(n_4533));
	notech_nand2 i_76059945(.A(n_61623), .B(read_data[15]), .Z(n_3228));
	notech_nand2 i_74559960(.A(n_61623), .B(read_data[12]), .Z(n_322367576)
		);
	notech_nand2 i_74059965(.A(n_61632), .B(read_data[11]), .Z(n_3216));
	notech_or4 i_42160252(.A(n_63718), .B(n_440667990), .C(n_63758), .D(nbus_11273
		[15]), .Z(n_320767568));
	notech_nao3 i_42460249(.A(n_63766), .B(opc[15]), .C(n_441868002), .Z(n_320367565
		));
	notech_nand2 i_42660248(.A(n_30354), .B(opd[15]), .Z(n_320067563));
	notech_or4 i_37660289(.A(n_384964380), .B(n_30553), .C(n_61933), .D(n_31623
		), .Z(n_319967562));
	notech_or2 i_37960286(.A(n_441668000), .B(\nbus_11290[12] ), .Z(n_319667559
		));
	notech_or4 i_38360283(.A(n_63718), .B(n_4533), .C(n_61933), .D(nbus_11273
		[12]), .Z(n_319367556));
	notech_or2 i_36960296(.A(n_441768001), .B(nbus_11273[11]), .Z(n_318467547
		));
	notech_nand2 i_37260293(.A(n_30354), .B(opd[11]), .Z(n_318167544));
	notech_or2 i_37360292(.A(n_30590), .B(n_433367917), .Z(n_317567542));
	notech_or2 i_18460458(.A(n_381764348), .B(nbus_11273[15]), .Z(n_315667524
		));
	notech_or4 i_19160451(.A(n_61871), .B(n_61675), .C(n_19680), .D(n_31523)
		, .Z(n_314867517));
	notech_or2 i_17260470(.A(n_386264393), .B(n_31488), .Z(n_314167510));
	notech_or4 i_17560467(.A(n_63718), .B(n_386364394), .C(n_63762), .D(nbus_11273
		[15]), .Z(n_313867507));
	notech_or2 i_13860504(.A(n_386264393), .B(n_31485), .Z(n_3128));
	notech_or4 i_14160501(.A(n_63718), .B(n_386364394), .C(n_63758), .D(nbus_11273
		[12]), .Z(n_312467498));
	notech_or2 i_12660516(.A(n_58702), .B(n_433367917), .Z(n_311467491));
	notech_or4 i_12960513(.A(n_63718), .B(n_386364394), .C(n_63754), .D(nbus_11273
		[11]), .Z(n_311167488));
	notech_nand2 i_79259913(.A(n_115442595), .B(n_32219), .Z(n_310667483));
	notech_nand2 i_77559930(.A(n_244036119), .B(n_25121), .Z(n_310567482));
	notech_nao3 i_77459931(.A(n_58597), .B(n_30495), .C(n_384764378), .Z(n_310467481
		));
	notech_nao3 i_77159934(.A(n_244036119), .B(n_58601), .C(n_384764378), .Z
		(n_310367480));
	notech_and3 i_48860679(.A(n_323167581), .B(n_323367583), .C(n_3228), .Z(n_310267479
		));
	notech_and3 i_48560682(.A(n_3234), .B(n_3236), .C(n_322367576), .Z(n_310167478
		));
	notech_and3 i_48160685(.A(n_323767585), .B(n_3239), .C(n_3216), .Z(n_310067477
		));
	notech_or2 i_48060686(.A(n_3610), .B(n_30719), .Z(n_309967476));
	notech_or2 i_46960690(.A(n_3609), .B(n_30719), .Z(n_309867475));
	notech_and4 i_106262336(.A(n_28158), .B(n_58055), .C(n_309467471), .D(n_309367470
		), .Z(n_309767474));
	notech_ao4 i_105562342(.A(n_24528), .B(n_33239), .C(n_24527), .D(n_33238
		), .Z(n_309467471));
	notech_and3 i_106162337(.A(n_309067467), .B(n_309267469), .C(n_293467311
		), .Z(n_309367470));
	notech_ao4 i_105762340(.A(n_60449), .B(n_31510), .C(n_24717), .D(n_336160989
		), .Z(n_309267469));
	notech_ao4 i_105962339(.A(n_381164342), .B(n_31474), .C(n_326160889), .D
		(n_380764338), .Z(n_309067467));
	notech_ao4 i_106362335(.A(n_381064341), .B(n_33167), .C(n_100842449), .D
		(n_380964340), .Z(n_308767464));
	notech_ao4 i_106462334(.A(n_325960887), .B(n_24430), .C(n_326360891), .D
		(n_24424), .Z(n_308667463));
	notech_and3 i_107262329(.A(n_294367320), .B(n_308267459), .C(n_308467461
		), .Z(n_308567462));
	notech_ao4 i_106762332(.A(n_326260890), .B(n_24421), .C(n_326660894), .D
		(n_24431), .Z(n_308467461));
	notech_ao4 i_106862331(.A(n_326460892), .B(n_24429), .C(n_326760895), .D
		(n_24425), .Z(n_308267459));
	notech_and4 i_116662235(.A(n_307967456), .B(n_307767454), .C(n_307667453
		), .D(n_294667323), .Z(n_308167458));
	notech_ao4 i_116162240(.A(n_24528), .B(n_33237), .C(n_24527), .D(n_33236
		), .Z(n_307967456));
	notech_ao4 i_116362238(.A(n_60449), .B(n_31519), .C(n_3753), .D(n_24542)
		, .Z(n_307767454));
	notech_ao4 i_116462237(.A(n_3752), .B(n_24541), .C(n_3751), .D(n_24539),
		 .Z(n_307667453));
	notech_and4 i_117262229(.A(n_307367450), .B(n_307167448), .C(n_307067447
		), .D(n_295367330), .Z(n_307567452));
	notech_ao4 i_116762234(.A(n_431067894), .B(n_381364344), .C(nbus_11273[
		11]), .D(n_381764348), .Z(n_307367450));
	notech_ao4 i_116962232(.A(n_381664347), .B(\nbus_11290[11] ), .C(n_3750)
		, .D(n_381564346), .Z(n_307167448));
	notech_ao4 i_117062231(.A(n_381264343), .B(n_31484), .C(n_61106), .D(n_30768
		), .Z(n_307067447));
	notech_and4 i_117862223(.A(n_58055), .B(n_306767444), .C(n_306567442), .D
		(n_306467441), .Z(n_306967446));
	notech_ao4 i_117362228(.A(n_3689), .B(n_24542), .C(n_381764348), .D(nbus_11273
		[12]), .Z(n_306767444));
	notech_ao4 i_117562226(.A(n_381664347), .B(\nbus_11290[12] ), .C(n_368667786
		), .D(n_381564346), .Z(n_306567442));
	notech_ao4 i_117662225(.A(n_3688), .B(n_24541), .C(n_368767787), .D(n_24539
		), .Z(n_306467441));
	notech_and4 i_118562216(.A(n_306167438), .B(n_306067437), .C(n_305867435
		), .D(n_305767434), .Z(n_306367440));
	notech_ao4 i_117962222(.A(n_381464345), .B(n_33250), .C(n_3907), .D(n_381364344
		), .Z(n_306167438));
	notech_ao4 i_118062221(.A(n_3609), .B(n_24716), .C(n_24528), .D(n_33235)
		, .Z(n_306067437));
	notech_ao4 i_118262219(.A(n_24527), .B(n_33234), .C(n_381264343), .D(n_31485
		), .Z(n_305867435));
	notech_ao4 i_118362218(.A(n_60449), .B(n_31520), .C(n_61106), .D(n_30769
		), .Z(n_305767434));
	notech_and4 i_123462172(.A(n_305467431), .B(n_305267429), .C(n_305167428
		), .D(n_326860896), .Z(n_305667433));
	notech_ao4 i_122762177(.A(n_326360891), .B(n_151069548), .C(n_383264363)
		, .D(n_61632), .Z(n_305467431));
	notech_ao4 i_122962175(.A(n_326260890), .B(n_150969547), .C(n_57027), .D
		(n_33167), .Z(n_305267429));
	notech_ao4 i_123062174(.A(n_100842449), .B(n_57036), .C(n_57438), .D(n_326160889
		), .Z(n_305167428));
	notech_and4 i_124062166(.A(n_304867425), .B(n_304667423), .C(n_304567422
		), .D(n_297967356), .Z(n_305067427));
	notech_ao4 i_123562171(.A(n_30473), .B(n_326060888), .C(n_325960887), .D
		(n_143769475), .Z(n_304867425));
	notech_ao4 i_123762169(.A(n_326660894), .B(n_143469472), .C(n_326460892)
		, .D(n_143569473), .Z(n_304667423));
	notech_ao4 i_123862168(.A(n_326560893), .B(n_143669474), .C(n_326760895)
		, .D(n_143369471), .Z(n_304567422));
	notech_or4 i_129262119(.A(n_298467361), .B(n_298767364), .C(n_30500), .D
		(n_30508), .Z(n_304467421));
	notech_ao4 i_129062121(.A(n_3751), .B(n_333978345), .C(n_323978248), .D(n_33258
		), .Z(n_304167418));
	notech_nand2 i_129462117(.A(n_303867415), .B(n_299067367), .Z(n_303967416
		));
	notech_ao4 i_129362118(.A(n_57243), .B(nbus_11273[11]), .C(n_57244), .D(\nbus_11290[11] 
		), .Z(n_303867415));
	notech_ao4 i_129562116(.A(n_30473), .B(n_433367917), .C(n_31484), .D(n_58030
		), .Z(n_303667413));
	notech_and4 i_162761788(.A(n_30274), .B(n_303367410), .C(n_303167408), .D
		(n_299867375), .Z(n_303567412));
	notech_ao4 i_162361792(.A(n_1532), .B(n_30891), .C(n_29993), .D(n_30916)
		, .Z(n_303367410));
	notech_ao4 i_162561790(.A(n_29994), .B(n_30914), .C(n_30191), .D(n_33103
		), .Z(n_303167408));
	notech_and4 i_163261783(.A(n_302867405), .B(n_302667403), .C(n_300167378
		), .D(n_300467381), .Z(n_303067407));
	notech_ao4 i_162861787(.A(n_291167288), .B(\nbus_11290[1] ), .C(n_3606),
		 .D(nbus_11273[1]), .Z(n_302867405));
	notech_ao4 i_163061785(.A(n_30896), .B(n_30576), .C(n_291067287), .D(n_30201
		), .Z(n_302667403));
	notech_and4 i_165461761(.A(n_300567382), .B(n_30274), .C(n_302267399), .D
		(n_300867385), .Z(n_302567402));
	notech_ao4 i_165261763(.A(n_323960867), .B(n_33103), .C(n_305344487), .D
		(n_31473), .Z(n_302267399));
	notech_ao4 i_165561760(.A(n_292067297), .B(\nbus_11290[1] ), .C(n_3607),
		 .D(nbus_11273[1]), .Z(n_302067397));
	notech_ao4 i_165661759(.A(n_291967296), .B(n_194866375), .C(n_291867295)
		, .D(n_336860996), .Z(n_301867395));
	notech_mux2 i_165961756(.S(n_323660864), .A(n_30896), .B(n_30914), .Z(n_301767394
		));
	notech_or2 i_31146(.A(n_28551), .B(n_30441), .Z(n_28252));
	notech_or2 i_31147(.A(n_439367977), .B(n_30441), .Z(n_28251));
	notech_ao4 i_31240(.A(n_331360941), .B(\nbus_11290[2] ), .C(n_28240), .D
		(nbus_11273[2]), .Z(n_28158));
	notech_or2 i_88762504(.A(n_57170), .B(n_30280), .Z(n_301367390));
	notech_or2 i_89262499(.A(n_323860866), .B(n_334360971), .Z(n_300867385)
		);
	notech_nao3 i_89362498(.A(n_323660864), .B(n_30484), .C(n_30916), .Z(n_300567382
		));
	notech_or2 i_85062539(.A(n_57122), .B(n_30280), .Z(n_300467381));
	notech_or2 i_85362536(.A(n_30196), .B(n_334360971), .Z(n_300167378));
	notech_or2 i_85662533(.A(n_305244486), .B(n_31473), .Z(n_299867375));
	notech_nor2 i_53362849(.A(n_3750), .B(n_57393), .Z(n_299367370));
	notech_or4 i_53662846(.A(n_58555), .B(n_256563512), .C(n_324078249), .D(n_431067894
		), .Z(n_299067367));
	notech_ao3 i_53962843(.A(n_63766), .B(opc[11]), .C(n_333778343), .Z(n_298767364
		));
	notech_ao3 i_54062842(.A(opa[11]), .B(n_30351), .C(n_60194), .Z(n_298467361
		));
	notech_or2 i_47462903(.A(n_5783), .B(n_31474), .Z(n_297967356));
	notech_or2 i_39562974(.A(n_381464345), .B(n_33258), .Z(n_295367330));
	notech_or2 i_40262967(.A(n_430767891), .B(n_24716), .Z(n_294667323));
	notech_or4 i_27763086(.A(n_61056), .B(n_24430), .C(\nbus_11290[2] ), .D(n_30664
		), .Z(n_294367320));
	notech_nand2 i_28763077(.A(sav_ecx[2]), .B(n_61871), .Z(n_293467311));
	notech_ao4 i_9663261(.A(n_323660864), .B(n_30919), .C(n_60177), .D(nbus_11273
		[1]), .Z(n_292467301));
	notech_ao4 i_9763260(.A(n_323660864), .B(n_30920), .C(n_60177), .D(\nbus_11290[1] 
		), .Z(n_292267299));
	notech_nao3 i_92869345(.A(n_3608), .B(n_32266), .C(n_184660383), .Z(n_292067297
		));
	notech_and2 i_13763222(.A(n_30891), .B(n_301767394), .Z(n_291967296));
	notech_mux2 i_13663223(.S(n_32266), .A(n_292467301), .B(n_292267299), .Z
		(n_291867295));
	notech_ao4 i_9863259(.A(n_30212), .B(n_30919), .C(n_60177), .D(nbus_11273
		[1]), .Z(n_291567292));
	notech_ao4 i_9963258(.A(n_30212), .B(n_30920), .C(n_60177), .D(\nbus_11290[1] 
		), .Z(n_291367290));
	notech_nao3 i_91869346(.A(n_30077), .B(n_32261), .C(n_1481), .Z(n_291167288
		));
	notech_mux2 i_13863221(.S(n_32261), .A(n_291567292), .B(n_291367290), .Z
		(n_291067287));
	notech_nand2 i_105863360(.A(n_330960937), .B(n_28552), .Z(n_290767284)
		);
	notech_nand2 i_104065128(.A(n_290367280), .B(n_238766787), .Z(n_290467281
		));
	notech_ao4 i_103965129(.A(n_3688), .B(n_333778343), .C(n_3907), .D(n_323778246
		), .Z(n_290367280));
	notech_or4 i_104665122(.A(n_239366793), .B(n_239066790), .C(n_30517), .D
		(n_30518), .Z(n_290267279));
	notech_ao4 i_104265126(.A(n_57244), .B(\nbus_11290[12] ), .C(n_57243), .D
		(nbus_11273[12]), .Z(n_290067277));
	notech_ao4 i_104465124(.A(n_30473), .B(n_309867475), .C(n_58030), .D(n_31485
		), .Z(n_289867275));
	notech_nand2 i_105665112(.A(n_289467271), .B(n_239766797), .Z(n_289567272
		));
	notech_ao4 i_105565113(.A(n_3692), .B(n_333778343), .C(n_3910), .D(n_323778246
		), .Z(n_289467271));
	notech_or4 i_106265106(.A(n_240366803), .B(n_240066800), .C(n_30525), .D
		(n_30527), .Z(n_289367270));
	notech_ao4 i_105865110(.A(n_57244), .B(\nbus_11290[15] ), .C(n_57243), .D
		(nbus_11273[15]), .Z(n_289167268));
	notech_ao4 i_106065108(.A(n_57068), .B(n_309967476), .C(n_58030), .D(n_31488
		), .Z(n_288967266));
	notech_ao4 i_107865091(.A(n_28240), .B(nbus_11273[2]), .C(n_26585), .D(n_30971
		), .Z(n_288667263));
	notech_ao4 i_107965090(.A(n_126126588), .B(n_32061), .C(n_125926586), .D
		(n_33233), .Z(n_288567262));
	notech_ao3 i_108465085(.A(n_288167258), .B(n_288367260), .C(n_241166811)
		, .Z(n_288467261));
	notech_ao4 i_108165088(.A(n_336160989), .B(n_26603), .C(n_26600), .D(n_31510
		), .Z(n_288367260));
	notech_ao4 i_108265087(.A(n_326560893), .B(n_26277), .C(n_326760895), .D
		(n_26276), .Z(n_288167258));
	notech_and4 i_109865075(.A(n_241666815), .B(n_287667253), .C(n_287867255
		), .D(n_287567252), .Z(n_288067257));
	notech_ao4 i_108665083(.A(n_326660894), .B(n_26275), .C(n_26271), .D(n_326260890
		), .Z(n_287867255));
	notech_ao4 i_108765082(.A(n_100842449), .B(n_332460952), .C(n_332260950)
		, .D(n_33167), .Z(n_287667253));
	notech_and3 i_109765076(.A(n_287267249), .B(n_287467251), .C(n_242166819
		), .Z(n_287567252));
	notech_ao4 i_109465079(.A(n_325960887), .B(n_26278), .C(n_326160889), .D
		(n_332160949), .Z(n_287467251));
	notech_ao4 i_109565078(.A(n_331160939), .B(\nbus_11290[2] ), .C(n_61106)
		, .D(n_30778), .Z(n_287267249));
	notech_and4 i_118764992(.A(n_286967246), .B(n_286767244), .C(n_286667243
		), .D(n_242466821), .Z(n_287167248));
	notech_ao4 i_118264997(.A(n_126126588), .B(n_32070), .C(n_125926586), .D
		(n_33232), .Z(n_286967246));
	notech_ao4 i_118464995(.A(n_430767891), .B(n_331560943), .C(n_26600), .D
		(n_31519), .Z(n_286767244));
	notech_ao4 i_118564994(.A(n_3753), .B(n_26397), .C(n_3751), .D(n_26396),
		 .Z(n_286667243));
	notech_and4 i_119464985(.A(n_286367240), .B(n_286267239), .C(n_286067237
		), .D(n_285967236), .Z(n_286567242));
	notech_ao4 i_118864991(.A(n_3752), .B(n_26394), .C(n_431067894), .D(n_378864319
		), .Z(n_286367240));
	notech_ao4 i_118964990(.A(n_378964320), .B(n_33258), .C(n_378664317), .D
		(\nbus_11290[11] ), .Z(n_286267239));
	notech_ao4 i_119164988(.A(n_378764318), .B(nbus_11273[11]), .C(n_3750), 
		.D(n_378564316), .Z(n_286067237));
	notech_ao4 i_119264987(.A(n_378464315), .B(n_31484), .C(n_61106), .D(n_30790
		), .Z(n_285967236));
	notech_and4 i_120064979(.A(n_285667233), .B(n_285467231), .C(n_285367230
		), .D(n_244166836), .Z(n_285867235));
	notech_ao4 i_119564984(.A(n_126126588), .B(n_32071), .C(n_125926586), .D
		(n_33231), .Z(n_285667233));
	notech_ao4 i_119764982(.A(n_3609), .B(n_331560943), .C(n_26600), .D(n_31520
		), .Z(n_285467231));
	notech_ao4 i_119864981(.A(n_3689), .B(n_26397), .C(n_368767787), .D(n_26396
		), .Z(n_285367230));
	notech_and4 i_120964972(.A(n_285067227), .B(n_284967226), .C(n_284767224
		), .D(n_284667223), .Z(n_285267229));
	notech_ao4 i_120164978(.A(n_3688), .B(n_26394), .C(n_3907), .D(n_378864319
		), .Z(n_285067227));
	notech_ao4 i_120464977(.A(n_378964320), .B(n_33250), .C(n_378664317), .D
		(\nbus_11290[12] ), .Z(n_284967226));
	notech_ao4 i_120664975(.A(n_378764318), .B(nbus_11273[12]), .C(n_368667786
		), .D(n_378564316), .Z(n_284767224));
	notech_ao4 i_120764974(.A(n_378464315), .B(n_31485), .C(n_61106), .D(n_30791
		), .Z(n_284667223));
	notech_and4 i_123064953(.A(n_284367220), .B(n_284167218), .C(n_284067217
		), .D(n_245766851), .Z(n_284567222));
	notech_ao4 i_122564958(.A(n_126126588), .B(n_32074), .C(n_125926586), .D
		(n_33230), .Z(n_284367220));
	notech_ao4 i_122764956(.A(n_3610), .B(n_331560943), .C(n_26600), .D(n_31523
		), .Z(n_284167218));
	notech_ao4 i_122864955(.A(n_3693), .B(n_26397), .C(n_3691), .D(n_26396),
		 .Z(n_284067217));
	notech_and4 i_123964946(.A(n_283767214), .B(n_283667213), .C(n_283467211
		), .D(n_283367210), .Z(n_283967216));
	notech_ao4 i_123164952(.A(n_3692), .B(n_26394), .C(n_3910), .D(n_378864319
		), .Z(n_283767214));
	notech_ao4 i_123264951(.A(n_378964320), .B(n_33248), .C(n_378664317), .D
		(\nbus_11290[15] ), .Z(n_283667213));
	notech_ao4 i_123464949(.A(n_378764318), .B(nbus_11273[15]), .C(n_3690), 
		.D(n_378564316), .Z(n_283467211));
	notech_ao4 i_123764948(.A(n_378464315), .B(n_31488), .C(n_61106), .D(n_30794
		), .Z(n_283367210));
	notech_and4 i_137864812(.A(n_283067207), .B(n_282867205), .C(n_282767204
		), .D(n_247266865), .Z(n_283267209));
	notech_ao4 i_137364817(.A(n_57012), .B(n_31519), .C(n_3753), .D(n_334278348
		), .Z(n_283067207));
	notech_ao4 i_137564815(.A(n_3751), .B(n_334178347), .C(n_3752), .D(n_334078346
		), .Z(n_282867205));
	notech_ao4 i_137664814(.A(n_431067894), .B(n_57275), .C(n_57274), .D(n_33258
		), .Z(n_282767204));
	notech_and4 i_138464806(.A(n_282467201), .B(n_282267199), .C(n_282167198
		), .D(n_247966872), .Z(n_282667203));
	notech_ao4 i_137964811(.A(n_57128), .B(nbus_11273[11]), .C(n_3750), .D(n_57394
		), .Z(n_282467201));
	notech_ao4 i_138164809(.A(n_58025), .B(n_31484), .C(n_61104), .D(n_30818
		), .Z(n_282267199));
	notech_ao4 i_138264808(.A(n_55913), .B(n_33229), .C(n_55793), .D(n_33228
		), .Z(n_282167198));
	notech_and4 i_139064800(.A(n_281867195), .B(n_281667193), .C(n_281567192
		), .D(n_248666879), .Z(n_282067197));
	notech_ao4 i_138564805(.A(n_57012), .B(n_31520), .C(n_3689), .D(n_334278348
		), .Z(n_281867195));
	notech_ao4 i_138764803(.A(n_368767787), .B(n_334178347), .C(n_3688), .D(n_334078346
		), .Z(n_281667193));
	notech_ao4 i_138864802(.A(n_3907), .B(n_57275), .C(n_57274), .D(n_33250)
		, .Z(n_281567192));
	notech_and4 i_139664794(.A(n_281267189), .B(n_281067187), .C(n_280967186
		), .D(n_249366886), .Z(n_281467191));
	notech_ao4 i_139164799(.A(n_57128), .B(nbus_11273[12]), .C(n_368667786),
		 .D(n_57394), .Z(n_281267189));
	notech_ao4 i_139364797(.A(n_58025), .B(n_31485), .C(n_61103), .D(n_30819
		), .Z(n_281067187));
	notech_ao4 i_139464796(.A(n_55913), .B(n_33227), .C(n_55793), .D(n_33226
		), .Z(n_280967186));
	notech_and4 i_141464776(.A(n_280667183), .B(n_280467181), .C(n_280367180
		), .D(n_250066893), .Z(n_280867185));
	notech_ao4 i_140964781(.A(n_57012), .B(n_31523), .C(n_3693), .D(n_334278348
		), .Z(n_280667183));
	notech_ao4 i_141164779(.A(n_3691), .B(n_334178347), .C(n_3692), .D(n_334078346
		), .Z(n_280467181));
	notech_ao4 i_141264778(.A(n_3910), .B(n_57275), .C(n_57274), .D(n_33248)
		, .Z(n_280367180));
	notech_and4 i_142064770(.A(n_280067177), .B(n_279867175), .C(n_279767174
		), .D(n_250766900), .Z(n_280267179));
	notech_ao4 i_141564775(.A(n_57128), .B(nbus_11273[15]), .C(n_3690), .D(n_57394
		), .Z(n_280067177));
	notech_ao4 i_141764773(.A(n_58025), .B(n_31488), .C(n_61103), .D(n_30821
		), .Z(n_279867175));
	notech_ao4 i_141864772(.A(n_55913), .B(n_33225), .C(n_330560933), .D(n_33224
		), .Z(n_279767174));
	notech_ao4 i_144164749(.A(n_245877510), .B(n_31520), .C(n_200777063), .D
		(n_3689), .Z(n_279567172));
	notech_ao4 i_144264748(.A(n_3688), .B(n_200677062), .C(n_3907), .D(n_57317
		), .Z(n_279367170));
	notech_and4 i_144964741(.A(n_279067167), .B(n_278867165), .C(n_251966912
		), .D(n_252266915), .Z(n_279267169));
	notech_ao4 i_144564745(.A(n_57133), .B(\nbus_11290[12] ), .C(n_57110), .D
		(nbus_11273[12]), .Z(n_279067167));
	notech_ao4 i_144764743(.A(n_57147), .B(n_309867475), .C(n_58053), .D(n_31485
		), .Z(n_278867165));
	notech_ao4 i_146864722(.A(n_178876848), .B(n_31523), .C(n_200777063), .D
		(n_3693), .Z(n_278667163));
	notech_ao4 i_146964721(.A(n_200677062), .B(n_3692), .C(n_3910), .D(n_57317
		), .Z(n_278467161));
	notech_and4 i_147664714(.A(n_278167158), .B(n_277967156), .C(n_253066923
		), .D(n_253366926), .Z(n_278367160));
	notech_ao4 i_147264718(.A(n_57133), .B(\nbus_11290[15] ), .C(n_57110), .D
		(nbus_11273[15]), .Z(n_278167158));
	notech_ao4 i_147464716(.A(n_57147), .B(n_309967476), .C(n_58053), .D(n_31488
		), .Z(n_277967156));
	notech_and4 i_149964691(.A(n_28158), .B(n_277567152), .C(n_118376249), .D
		(n_253466927), .Z(n_277767154));
	notech_ao4 i_149864692(.A(n_333260960), .B(n_33223), .C(n_333360961), .D
		(n_33222), .Z(n_277567152));
	notech_ao4 i_150064690(.A(n_326260890), .B(n_28252), .C(n_326360891), .D
		(n_28251), .Z(n_277367150));
	notech_ao4 i_150164689(.A(n_439667980), .B(n_100842449), .C(n_439567979)
		, .D(n_33167), .Z(n_277267149));
	notech_and4 i_151064680(.A(n_276967146), .B(n_276867145), .C(n_276667143
		), .D(n_276567142), .Z(n_277167148));
	notech_ao4 i_150464686(.A(n_326160889), .B(n_439367977), .C(n_439467978)
		, .D(n_31474), .Z(n_276967146));
	notech_ao4 i_150564685(.A(n_61103), .B(n_30834), .C(n_325960887), .D(n_28260
		), .Z(n_276867145));
	notech_ao4 i_150764683(.A(n_326560893), .B(n_28255), .C(n_326760895), .D
		(n_28258), .Z(n_276667143));
	notech_ao4 i_150864682(.A(n_326460892), .B(n_28259), .C(n_326660894), .D
		(n_28256), .Z(n_276567142));
	notech_and4 i_159864594(.A(n_276267139), .B(n_276067137), .C(n_275967136
		), .D(n_255166944), .Z(n_276467141));
	notech_ao4 i_159364599(.A(n_333260960), .B(n_33221), .C(n_333360961), .D
		(n_33220), .Z(n_276267139));
	notech_ao4 i_159564597(.A(n_3753), .B(n_28368), .C(n_57006), .D(n_31519)
		, .Z(n_276067137));
	notech_ao4 i_159664596(.A(n_3751), .B(n_28365), .C(n_3752), .D(n_28367),
		 .Z(n_275967136));
	notech_and4 i_160464588(.A(n_275667133), .B(n_275467131), .C(n_275367130
		), .D(n_255766950), .Z(n_275867135));
	notech_ao4 i_159964593(.A(n_444568029), .B(n_33258), .C(n_444468028), .D
		(\nbus_11290[11] ), .Z(n_275667133));
	notech_ao4 i_160164591(.A(n_444368027), .B(nbus_11273[11]), .C(n_444768031
		), .D(n_3750), .Z(n_275467131));
	notech_ao4 i_160264590(.A(n_444868032), .B(n_31484), .C(n_61104), .D(n_30846
		), .Z(n_275367130));
	notech_and4 i_161064582(.A(n_275067127), .B(n_274867125), .C(n_274767124
		), .D(n_256466957), .Z(n_275267129));
	notech_ao4 i_160564587(.A(n_333260960), .B(n_33219), .C(n_333360961), .D
		(n_33218), .Z(n_275067127));
	notech_ao4 i_160764585(.A(n_28368), .B(n_3689), .C(n_57001), .D(n_31520)
		, .Z(n_274867125));
	notech_ao4 i_160864584(.A(n_28365), .B(n_368767787), .C(n_28367), .D(n_3688
		), .Z(n_274767124));
	notech_and4 i_161664576(.A(n_2744), .B(n_274267120), .C(n_274167119), .D
		(n_257066963), .Z(n_274667123));
	notech_ao4 i_161164581(.A(n_444568029), .B(n_33250), .C(n_444468028), .D
		(\nbus_11290[12] ), .Z(n_2744));
	notech_ao4 i_161364579(.A(n_444368027), .B(nbus_11273[12]), .C(n_444768031
		), .D(n_368667786), .Z(n_274267120));
	notech_ao4 i_161464578(.A(n_444868032), .B(n_31485), .C(n_61104), .D(n_30847
		), .Z(n_274167119));
	notech_and4 i_164464548(.A(n_273867116), .B(n_273667114), .C(n_273567113
		), .D(n_257766970), .Z(n_274067118));
	notech_ao4 i_163964553(.A(n_333260960), .B(n_33217), .C(n_333360961), .D
		(n_33216), .Z(n_273867116));
	notech_ao4 i_164164551(.A(n_28368), .B(n_3693), .C(n_57001), .D(n_31523)
		, .Z(n_273667114));
	notech_ao4 i_164264550(.A(n_28365), .B(n_3691), .C(n_28367), .D(n_3692),
		 .Z(n_273567113));
	notech_and4 i_165064542(.A(n_273267110), .B(n_272967108), .C(n_272867107
		), .D(n_258366976), .Z(n_273467112));
	notech_ao4 i_164564547(.A(n_444568029), .B(n_33248), .C(n_444468028), .D
		(\nbus_11290[15] ), .Z(n_273267110));
	notech_ao4 i_164764545(.A(n_444368027), .B(nbus_11273[15]), .C(n_444768031
		), .D(n_3690), .Z(n_272967108));
	notech_ao4 i_164864544(.A(n_444868032), .B(n_31488), .C(n_61103), .D(n_30850
		), .Z(n_272867107));
	notech_and4 i_172864464(.A(n_272567104), .B(n_272367102), .C(n_310067477
		), .D(n_259266985), .Z(n_272767106));
	notech_ao4 i_172464468(.A(n_279977810), .B(nbus_11271[11]), .C(n_3753), 
		.D(n_334478350), .Z(n_272567104));
	notech_ao4 i_172664466(.A(n_3752), .B(n_334378349), .C(n_431067894), .D(n_323378242
		), .Z(n_272367102));
	notech_and4 i_173364459(.A(n_271767099), .B(n_271567097), .C(n_259566988
		), .D(n_259866991), .Z(n_272167101));
	notech_ao4 i_172964463(.A(n_57238), .B(n_58974), .C(n_57237), .D(n_58312
		), .Z(n_271767099));
	notech_ao4 i_173164461(.A(n_57609), .B(n_433367917), .C(n_31484), .D(n_58029
		), .Z(n_271567097));
	notech_and4 i_173864454(.A(n_271267094), .B(n_271067092), .C(n_310167478
		), .D(n_260366996), .Z(n_271467096));
	notech_ao4 i_173464458(.A(n_279977810), .B(nbus_11271[12]), .C(n_3689), 
		.D(n_334478350), .Z(n_271267094));
	notech_ao4 i_173664456(.A(n_3688), .B(n_334378349), .C(n_3907), .D(n_323378242
		), .Z(n_271067092));
	notech_and4 i_174364449(.A(n_270667089), .B(n_2704), .C(n_260666999), .D
		(n_261067002), .Z(n_270867091));
	notech_ao4 i_173964453(.A(n_57238), .B(n_59050), .C(n_57237), .D(n_58321
		), .Z(n_270667089));
	notech_ao4 i_174164451(.A(n_57604), .B(n_309867475), .C(n_58029), .D(n_31485
		), .Z(n_2704));
	notech_and4 i_176664426(.A(n_270067085), .B(n_269867083), .C(n_310267479
		), .D(n_261567007), .Z(n_270267087));
	notech_ao4 i_176264430(.A(n_279977810), .B(nbus_11271[15]), .C(n_3693), 
		.D(n_334478350), .Z(n_270067085));
	notech_ao4 i_176464428(.A(n_3692), .B(n_334378349), .C(n_3910), .D(n_323378242
		), .Z(n_269867083));
	notech_and4 i_177164421(.A(n_269567080), .B(n_269367078), .C(n_261867010
		), .D(n_262167013), .Z(n_269767082));
	notech_ao4 i_176764425(.A(n_57238), .B(n_59068), .C(n_57237), .D(nbus_11273
		[15]), .Z(n_269567080));
	notech_ao4 i_176964423(.A(n_57604), .B(n_309967476), .C(n_58029), .D(n_31488
		), .Z(n_269367078));
	notech_nand2 i_181964373(.A(n_268967074), .B(n_262667017), .Z(n_269067075
		));
	notech_ao4 i_181864374(.A(n_3752), .B(n_29418), .C(n_57611), .D(n_431067894
		), .Z(n_268967074));
	notech_or4 i_182564367(.A(n_263267023), .B(n_262967020), .C(n_30561), .D
		(n_30562), .Z(n_268867073));
	notech_ao4 i_182164371(.A(n_444968033), .B(n_58974), .C(n_445068034), .D
		(n_58312), .Z(n_268667071));
	notech_ao4 i_182364369(.A(n_57064), .B(n_433367917), .C(n_445268036), .D
		(n_31484), .Z(n_268467069));
	notech_nand2 i_182964364(.A(n_268067065), .B(n_263667027), .Z(n_268167066
		));
	notech_ao4 i_182864365(.A(n_29418), .B(n_3688), .C(n_57611), .D(n_3907),
		 .Z(n_268067065));
	notech_or4 i_183564358(.A(n_264267033), .B(n_263967030), .C(n_30563), .D
		(n_30564), .Z(n_267967064));
	notech_ao4 i_183164362(.A(n_444968033), .B(n_59050), .C(n_445068034), .D
		(n_58321), .Z(n_267767062));
	notech_ao4 i_183364360(.A(n_57064), .B(n_309867475), .C(n_445268036), .D
		(n_31485), .Z(n_267567060));
	notech_nand2 i_185464339(.A(n_267167056), .B(n_264667037), .Z(n_267267057
		));
	notech_ao4 i_185364340(.A(n_29418), .B(n_3692), .C(n_57611), .D(n_3910),
		 .Z(n_267167056));
	notech_or4 i_186064333(.A(n_265267043), .B(n_264967040), .C(n_30565), .D
		(n_30566), .Z(n_266867055));
	notech_ao4 i_185664337(.A(n_444968033), .B(n_59068), .C(n_445068034), .D
		(n_58348), .Z(n_266667053));
	notech_ao4 i_185864335(.A(n_57064), .B(n_309967476), .C(n_445268036), .D
		(n_31488), .Z(n_266067051));
	notech_ao4 i_189164302(.A(n_31532), .B(n_61675), .C(n_30695), .D(\nbus_11283[24] 
		), .Z(n_265967050));
	notech_ao4 i_189264301(.A(n_30697), .B(n_33171), .C(n_30689), .D(n_106826395
		), .Z(n_265767048));
	notech_nor2 i_100165167(.A(n_30693), .B(n_58893), .Z(n_265667047));
	notech_nao3 i_1566141(.A(n_30441), .B(n_57417), .C(n_439367977), .Z(n_28259
		));
	notech_or4 i_1066146(.A(n_2383), .B(n_439367977), .C(n_32159), .D(n_32161
		), .Z(n_28258));
	notech_or2 i_1666140(.A(n_439367977), .B(n_32544), .Z(n_28256));
	notech_or4 i_966147(.A(n_2383), .B(n_28260), .C(n_32159), .D(n_32161), .Z
		(n_28255));
	notech_nor2 i_98165187(.A(n_445168035), .B(n_3690), .Z(n_265267043));
	notech_ao3 i_98465184(.A(n_30282), .B(\opa_12[15] ), .C(n_386964400), .Z
		(n_264967040));
	notech_or4 i_98765181(.A(n_30269), .B(n_29560), .C(n_61933), .D(n_31626)
		, .Z(n_264667037));
	notech_ao3 i_98865180(.A(opa[15]), .B(n_29417), .C(n_60194), .Z(n_264367034
		));
	notech_nor2 i_95365215(.A(n_445168035), .B(n_368667786), .Z(n_264267033)
		);
	notech_ao3 i_95665212(.A(n_30282), .B(\opa_12[12] ), .C(n_386964400), .Z
		(n_263967030));
	notech_or4 i_95965209(.A(n_30269), .B(n_29560), .C(n_61933), .D(n_31623)
		, .Z(n_263667027));
	notech_ao3 i_96065208(.A(opa[12]), .B(n_29417), .C(n_60194), .Z(n_263367024
		));
	notech_nor2 i_94365225(.A(n_445168035), .B(n_3750), .Z(n_263267023));
	notech_ao3 i_94665222(.A(n_30282), .B(\opa_12[11] ), .C(n_386964400), .Z
		(n_262967020));
	notech_or4 i_94965219(.A(n_61933), .B(n_31622), .C(n_30269), .D(n_29560)
		, .Z(n_262667017));
	notech_ao4 i_130273235(.A(n_293792280), .B(n_31290), .C(n_57435), .D(n_31026
		), .Z(n_208580591));
	notech_ao4 i_130173236(.A(n_292192264), .B(n_4428), .C(n_292292265), .D(n_31323
		), .Z(n_208680592));
	notech_or4 i_41871562(.A(n_28534), .B(n_25713), .C(n_61871), .D(n_61630)
		, .Z(n_208780593));
	notech_and4 i_50238(.A(n_341381880), .B(n_342481891), .C(n_330281779), .D
		(n_208780593), .Z(n_208880594));
	notech_nao3 i_43071550(.A(n_32506), .B(n_4338), .C(n_4085), .Z(n_209180597
		));
	notech_or4 i_43171549(.A(n_340981876), .B(n_57336), .C(n_415382405), .D(n_27823
		), .Z(n_209280598));
	notech_nand3 i_43571545(.A(n_579), .B(n_32485), .C(n_19698), .Z(n_209380599
		));
	notech_ao4 i_55158(.A(n_333681811), .B(n_345881925), .C(n_239446886), .D
		(n_33496), .Z(n_209580601));
	notech_nand2 i_58371397(.A(n_4088), .B(n_209780603), .Z(n_209680602));
	notech_or2 i_58471396(.A(n_57001), .B(n_239346885), .Z(n_209780603));
	notech_nand2 i_2269241(.A(n_321860846), .B(n_57122), .Z(n_211080616));
	notech_nand3 i_2469239(.A(n_321860846), .B(n_57122), .C(n_63754), .Z(n_211480617
		));
	notech_nao3 i_2369240(.A(n_323060858), .B(n_211480617), .C(n_322960857),
		 .Z(n_211680619));
	notech_nand2 i_2569238(.A(n_219380694), .B(n_219280693), .Z(n_211780620)
		);
	notech_and4 i_2669237(.A(n_322760855), .B(n_322860856), .C(n_218880689),
		 .D(n_211080616), .Z(n_211880621));
	notech_or2 i_3669227(.A(n_212080623), .B(n_30266), .Z(n_211980622));
	notech_ao4 i_2769236(.A(n_323160859), .B(instrc[124]), .C(n_304344477), 
		.D(n_219180692), .Z(n_212080623));
	notech_or4 i_3769226(.A(instrc[121]), .B(n_111445606), .C(n_2577), .D(n_32161
		), .Z(n_212380626));
	notech_nao3 i_3269231(.A(n_63796), .B(n_30212), .C(n_218880689), .Z(n_212480627
		));
	notech_nand3 i_3369230(.A(instrc[119]), .B(n_275560604), .C(n_211680619)
		, .Z(n_212580628));
	notech_nand2 i_3469229(.A(n_30869), .B(n_211780620), .Z(n_212680629));
	notech_or4 i_3569228(.A(instrc[121]), .B(n_1481), .C(n_211880621), .D(n_32305
		), .Z(n_212780630));
	notech_and4 i_53765(.A(n_219980700), .B(n_212780630), .C(n_212680629), .D
		(n_211980622), .Z(n_212880631));
	notech_and2 i_15869107(.A(n_32203), .B(imm[31]), .Z(n_212980632));
	notech_nand2 i_44468842(.A(n_213280635), .B(opa[14]), .Z(n_213180634));
	notech_ao4 i_43568851(.A(n_304244476), .B(n_33214), .C(n_30077), .D(n_30483
		), .Z(n_213280635));
	notech_nao3 i_43768849(.A(n_30212), .B(n_30428), .C(n_377264303), .Z(n_213380636
		));
	notech_and4 i_1520845(.A(n_220780708), .B(n_220680707), .C(n_220580706),
		 .D(n_213180634), .Z(n_214080643));
	notech_or2 i_65068641(.A(n_29758), .B(n_379364324), .Z(n_214180644));
	notech_nand2 i_65868633(.A(n_214380646), .B(opa[14]), .Z(n_214280645));
	notech_nand2 i_64968642(.A(n_214180644), .B(n_376964300), .Z(n_214380646
		));
	notech_nao3 i_65168640(.A(n_63786), .B(opc_10[14]), .C(n_442182452), .Z(n_214480647
		));
	notech_and4 i_1520973(.A(n_221480715), .B(n_221380714), .C(n_221280713),
		 .D(n_214280645), .Z(n_215180654));
	notech_ao3 i_74768544(.A(opa[9]), .B(n_442082451), .C(n_60194), .Z(n_215380655
		));
	notech_or2 i_75668535(.A(n_62142062), .B(n_31482), .Z(n_216380664));
	notech_nand3 i_1020968(.A(n_221880719), .B(n_221780718), .C(n_222580726)
		, .Z(n_216480665));
	notech_and2 i_84368452(.A(n_3770), .B(n_445968043), .Z(n_216580666));
	notech_and2 i_84468451(.A(n_446068044), .B(n_214180644), .Z(n_216680667)
		);
	notech_or4 i_84668449(.A(n_379164322), .B(n_327760905), .C(n_33173), .D(n_30733
		), .Z(n_216780668));
	notech_nao3 i_85168444(.A(n_63786), .B(opc[0]), .C(n_376764298), .Z(n_217280673
		));
	notech_and4 i_120959(.A(n_222980730), .B(n_222880729), .C(n_223280733), 
		.D(n_222780728), .Z(n_217580676));
	notech_ao3 i_178967577(.A(n_60605), .B(\nbus_11290[31] ), .C(n_56428), .Z
		(n_217680677));
	notech_ao4 i_178867578(.A(n_4424), .B(n_384582276), .C(n_4347), .D(n_212980632
		), .Z(n_218580686));
	notech_ao3 i_179067576(.A(opb[31]), .B(nbus_11271[31]), .C(n_56428), .Z(n_218680687
		));
	notech_or4 i_3212926(.A(n_218580686), .B(n_218680687), .C(n_217680677), 
		.D(n_30347), .Z(n_218780688));
	notech_ao4 i_144969285(.A(n_57638), .B(n_2810), .C(n_30798), .D(n_125342694
		), .Z(n_218880689));
	notech_nao3 i_2969234(.A(n_63818), .B(n_33162), .C(n_211880621), .Z(n_219180692
		));
	notech_ao4 i_1569248(.A(n_30554), .B(n_30248), .C(n_30751), .D(n_4464), 
		.Z(n_219280693));
	notech_ao4 i_1869245(.A(n_30815), .B(n_375464285), .C(n_30822), .D(n_375364284
		), .Z(n_219380694));
	notech_ao4 i_3969224(.A(n_57122), .B(n_114845640), .C(n_30835), .D(n_375564286
		), .Z(n_219680697));
	notech_and4 i_4269221(.A(n_212380626), .B(n_219680697), .C(n_212480627),
		 .D(n_212580628), .Z(n_219980700));
	notech_or4 i_169258(.A(n_32589), .B(n_28534), .C(n_60157), .D(n_61632), 
		.Z(n_220280703));
	notech_ao4 i_44868840(.A(n_304644480), .B(n_97342414), .C(n_377164302), 
		.D(n_30075), .Z(n_220480705));
	notech_and3 i_45168837(.A(n_220480705), .B(n_377364304), .C(n_213380636)
		, .Z(n_220580706));
	notech_ao4 i_44968839(.A(n_4924), .B(\nbus_11290[14] ), .C(n_304744481),
		 .D(n_33215), .Z(n_220680707));
	notech_ao4 i_45068838(.A(n_4922), .B(n_31487), .C(n_377064301), .D(n_57122
		), .Z(n_220780708));
	notech_ao4 i_66068631(.A(n_445968043), .B(n_97342414), .C(n_377164302), 
		.D(n_4418), .Z(n_221180712));
	notech_and3 i_66368628(.A(n_221180712), .B(n_377364304), .C(n_214480647)
		, .Z(n_221280713));
	notech_ao4 i_66168630(.A(n_62742068), .B(\nbus_11290[14] ), .C(n_446068044
		), .D(n_33215), .Z(n_221380714));
	notech_ao4 i_66268629(.A(n_62142062), .B(n_31487), .C(n_377064301), .D(n_57141
		), .Z(n_221480715));
	notech_ao4 i_76068531(.A(n_62642067), .B(nbus_11273[9]), .C(n_62742068),
		 .D(\nbus_11290[9] ), .Z(n_221780718));
	notech_ao4 i_76168530(.A(n_326960897), .B(n_57141), .C(n_327060898), .D(n_62442065
		), .Z(n_221880719));
	notech_nor2 i_75768534(.A(n_215380655), .B(n_30917), .Z(n_222080721));
	notech_ao4 i_75868533(.A(n_327160899), .B(n_4418), .C(n_327260900), .D(n_442182452
		), .Z(n_222280723));
	notech_ao4 i_75968532(.A(n_446068044), .B(n_33168), .C(n_445968043), .D(n_99942440
		), .Z(n_222380724));
	notech_and4 i_76568526(.A(n_222380724), .B(n_222280723), .C(n_216380664)
		, .D(n_222080721), .Z(n_222580726));
	notech_and3 i_85768438(.A(n_327860906), .B(n_216780668), .C(n_217280673)
		, .Z(n_222780728));
	notech_ao4 i_85568440(.A(n_376964300), .B(n_33169), .C(n_376864299), .D(n_101142452
		), .Z(n_222880729));
	notech_ao4 i_85668439(.A(n_54741988), .B(n_31472), .C(n_57141), .D(n_327560903
		), .Z(n_222980730));
	notech_ao4 i_86068435(.A(nbus_11273[0]), .B(n_216680667), .C(\nbus_11290[0] 
		), .D(n_216580666), .Z(n_223280733));
	notech_ao4 i_179167575(.A(n_4348), .B(n_31539), .C(n_112042561), .D(n_32345
		), .Z(n_223380734));
	notech_ao4 i_179267574(.A(n_4350), .B(n_33463), .C(n_4349), .D(n_33462),
		 .Z(n_223480735));
	notech_ao4 i_179367573(.A(n_4351), .B(n_32912), .C(n_24142), .D(n_33464)
		, .Z(n_223680737));
	notech_ao4 i_179467572(.A(n_4353), .B(nbus_11271[31]), .C(n_4352), .D(\nbus_11283[31] 
		), .Z(n_223780738));
	notech_and4 i_179767569(.A(n_223780738), .B(n_223680737), .C(n_223480735
		), .D(n_223380734), .Z(n_223980740));
	notech_or2 i_21165946(.A(n_26585), .B(n_30985), .Z(n_224480745));
	notech_or2 i_30165860(.A(n_26585), .B(n_31028), .Z(n_225980760));
	notech_or2 i_29765863(.A(n_337761005), .B(nbus_11271[30]), .Z(n_226280763
		));
	notech_or2 i_29365866(.A(n_126926596), .B(n_33194), .Z(n_226580766));
	notech_or2 i_68465484(.A(n_336660994), .B(n_331760945), .Z(n_227280773)
		);
	notech_or2 i_67765491(.A(n_99942440), .B(n_444668030), .Z(n_227980780)
		);
	notech_or4 i_78465384(.A(n_63718), .B(n_57666), .C(n_63754), .D(nbus_11273
		[2]), .Z(n_229280793));
	notech_or4 i_81065358(.A(n_63718), .B(n_57666), .C(n_63780), .D(nbus_11273
		[7]), .Z(n_230580806));
	notech_or4 i_82565343(.A(n_61933), .B(n_31620), .C(n_30319), .D(n_323578244
		), .Z(n_231480815));
	notech_nao3 i_82265346(.A(n_30300), .B(\opa_12[9] ), .C(n_376064291), .Z
		(n_231780818));
	notech_or4 i_81965349(.A(n_63718), .B(n_57387), .C(n_63754), .D(nbus_11273
		[9]), .Z(n_232080821));
	notech_or2 i_89865270(.A(n_386464395), .B(n_31474), .Z(n_232980830));
	notech_or2 i_92465244(.A(n_386464395), .B(n_31480), .Z(n_234280843));
	notech_ao3 i_94065228(.A(opa[9]), .B(n_29417), .C(n_60194), .Z(n_234780848
		));
	notech_or4 i_93965229(.A(n_61938), .B(n_31620), .C(n_30269), .D(n_29560)
		, .Z(n_235080851));
	notech_ao3 i_93665232(.A(n_30282), .B(\opa_12[9] ), .C(n_386964400), .Z(n_235380854
		));
	notech_nor2 i_93365235(.A(n_327060898), .B(n_445168035), .Z(n_235680857)
		);
	notech_nao3 i_32411(.A(n_33153), .B(n_33162), .C(n_323160859), .Z(n_26987
		));
	notech_or4 i_32420(.A(n_30449), .B(instrc[99]), .C(n_30618), .D(n_30343)
		, .Z(n_26978));
	notech_ao4 i_181464378(.A(n_326960897), .B(n_57064), .C(n_445268036), .D
		(n_31482), .Z(n_235880859));
	notech_ao4 i_181264380(.A(n_444968033), .B(\nbus_11290[9] ), .C(n_445068034
		), .D(nbus_11273[9]), .Z(n_236080861));
	notech_or4 i_181664376(.A(n_235680857), .B(n_235380854), .C(n_30349), .D
		(n_30348), .Z(n_236280863));
	notech_ao4 i_180964383(.A(n_29418), .B(n_327160899), .C(n_99942440), .D(n_57611
		), .Z(n_236380864));
	notech_nand2 i_181064382(.A(n_236380864), .B(n_235080851), .Z(n_236480865
		));
	notech_ao4 i_180564387(.A(n_324260870), .B(n_29337), .C(n_324360871), .D
		(n_29340), .Z(n_236780868));
	notech_ao4 i_180464388(.A(n_324760875), .B(n_29341), .C(n_324460872), .D
		(n_29338), .Z(n_236880869));
	notech_ao4 i_180264390(.A(n_323760865), .B(n_57064), .C(n_29533), .D(\nbus_11290[7] 
		), .Z(n_237080871));
	notech_and4 i_180764385(.A(n_237080871), .B(n_236880869), .C(n_236780868
		), .D(n_234280843), .Z(n_237280873));
	notech_ao4 i_179964393(.A(n_324160869), .B(n_29342), .C(n_324060868), .D
		(n_378364314), .Z(n_237380874));
	notech_ao4 i_179864394(.A(n_100242443), .B(n_29540), .C(n_29550), .D(n_33165
		), .Z(n_237480875));
	notech_ao4 i_179664396(.A(n_324660874), .B(n_29334), .C(n_324560873), .D
		(n_29333), .Z(n_237680877));
	notech_and4 i_180164391(.A(n_324860876), .B(n_237680877), .C(n_237480875
		), .D(n_237380874), .Z(n_237880879));
	notech_ao4 i_178164411(.A(n_326660894), .B(n_29337), .C(n_29340), .D(n_326560893
		), .Z(n_237980880));
	notech_ao4 i_178064412(.A(n_326460892), .B(n_29341), .C(n_326760895), .D
		(n_29338), .Z(n_238080881));
	notech_ao4 i_177864414(.A(n_326060888), .B(n_57064), .C(n_29533), .D(\nbus_11290[2] 
		), .Z(n_238280883));
	notech_and4 i_178364409(.A(n_238280883), .B(n_238080881), .C(n_237980880
		), .D(n_232980830), .Z(n_238480885));
	notech_ao4 i_177564417(.A(n_325960887), .B(n_29342), .C(n_326160889), .D
		(n_378364314), .Z(n_238580886));
	notech_ao4 i_177464418(.A(n_100842449), .B(n_29540), .C(n_29550), .D(n_33167
		), .Z(n_238680887));
	notech_ao4 i_177264420(.A(n_326260890), .B(n_29334), .C(n_326360891), .D
		(n_29333), .Z(n_238880889));
	notech_and4 i_177764415(.A(n_238880889), .B(n_238680887), .C(n_238580886
		), .D(n_326860896), .Z(n_239080891));
	notech_ao4 i_171164481(.A(n_326960897), .B(n_57604), .C(n_58029), .D(n_31482
		), .Z(n_239180892));
	notech_ao4 i_170964483(.A(n_57238), .B(\nbus_11290[9] ), .C(n_57237), .D
		(nbus_11273[9]), .Z(n_239380894));
	notech_and4 i_171364479(.A(n_239380894), .B(n_239180892), .C(n_231780818
		), .D(n_232080821), .Z(n_239580896));
	notech_ao4 i_170664486(.A(n_327160899), .B(n_334378349), .C(n_99942440),
		 .D(n_323378242), .Z(n_239680897));
	notech_ao4 i_170464488(.A(n_279977810), .B(nbus_11271[9]), .C(n_327360901
		), .D(n_334478350), .Z(n_239880899));
	notech_and4 i_170864484(.A(n_239880899), .B(n_239680897), .C(n_231480815
		), .D(n_327460902), .Z(n_240080901));
	notech_ao4 i_170164491(.A(n_324460872), .B(n_140176467), .C(n_324360871)
		, .D(n_139876464), .Z(n_240180902));
	notech_ao4 i_170064492(.A(n_324260870), .B(n_140076466), .C(n_324760875)
		, .D(n_139976465), .Z(n_240280903));
	notech_ao4 i_169864494(.A(n_323760865), .B(n_57604), .C(n_58044), .D(n_31480
		), .Z(n_240480905));
	notech_and4 i_170364489(.A(n_230580806), .B(n_240480905), .C(n_240280903
		), .D(n_240180902), .Z(n_240680907));
	notech_ao4 i_169564497(.A(n_192676984), .B(n_33165), .C(n_324160869), .D
		(n_169676762), .Z(n_240780908));
	notech_ao4 i_169464498(.A(n_324560873), .B(n_200477060), .C(n_100242443)
		, .D(n_323278241), .Z(n_240880909));
	notech_ao4 i_169264500(.A(n_279977810), .B(nbus_11271[7]), .C(n_324660874
		), .D(n_200377059), .Z(n_241080911));
	notech_and4 i_169764495(.A(n_324860876), .B(n_241080911), .C(n_240880909
		), .D(n_240780908), .Z(n_241280913));
	notech_ao4 i_167764515(.A(n_326760895), .B(n_140176467), .C(n_326560893)
		, .D(n_139876464), .Z(n_241380914));
	notech_ao4 i_167664516(.A(n_326660894), .B(n_140076466), .C(n_326460892)
		, .D(n_139976465), .Z(n_241480915));
	notech_ao4 i_167464518(.A(n_326060888), .B(n_57604), .C(n_58044), .D(n_31474
		), .Z(n_241680917));
	notech_and4 i_167964513(.A(n_241680917), .B(n_241480915), .C(n_241380914
		), .D(n_229280793), .Z(n_241880919));
	notech_ao4 i_167164521(.A(n_192676984), .B(n_33167), .C(n_325960887), .D
		(n_169676762), .Z(n_241980920));
	notech_ao4 i_167064522(.A(n_200477060), .B(n_326360891), .C(n_100842449)
		, .D(n_323278241), .Z(n_242080921));
	notech_ao4 i_166864524(.A(n_279977810), .B(nbus_11271[2]), .C(n_326260890
		), .D(n_200377059), .Z(n_242380923));
	notech_and4 i_167364519(.A(n_242380923), .B(n_242080921), .C(n_241980920
		), .D(n_326860896), .Z(n_242680925));
	notech_ao4 i_157864614(.A(n_444868032), .B(n_31482), .C(n_61103), .D(n_30844
		), .Z(n_242780926));
	notech_ao4 i_157764615(.A(n_444368027), .B(nbus_11273[9]), .C(n_327060898
		), .D(n_444768031), .Z(n_242980927));
	notech_ao4 i_157564617(.A(n_444568029), .B(n_33168), .C(n_444468028), .D
		(\nbus_11290[9] ), .Z(n_243280929));
	notech_and4 i_158064612(.A(n_243280929), .B(n_242980927), .C(n_242780926
		), .D(n_227980780), .Z(n_243680931));
	notech_ao4 i_157264620(.A(n_327260900), .B(n_28365), .C(n_327160899), .D
		(n_28367), .Z(n_243880932));
	notech_ao4 i_157164621(.A(n_57001), .B(n_31517), .C(n_327360901), .D(n_28368
		), .Z(n_243980933));
	notech_ao4 i_156964623(.A(n_333260960), .B(n_33466), .C(n_333360961), .D
		(n_33465), .Z(n_244380935));
	notech_and4 i_157464618(.A(n_244380935), .B(n_243980933), .C(n_243880932
		), .D(n_227280773), .Z(n_244680937));
	notech_ao4 i_124864937(.A(n_26600), .B(n_31538), .C(n_61103), .D(n_30808
		), .Z(n_244780938));
	notech_ao4 i_124764938(.A(n_337861006), .B(n_31506), .C(n_126226589), .D
		(n_5750), .Z(n_244880939));
	notech_ao4 i_124564940(.A(n_126726594), .B(\nbus_11283[30] ), .C(n_126826595
		), .D(\nbus_11290[30] ), .Z(n_245080941));
	notech_and4 i_125164935(.A(n_245080941), .B(n_244880939), .C(n_244780938
		), .D(n_226580766), .Z(n_245280943));
	notech_ao4 i_124264943(.A(n_337961007), .B(n_318771158), .C(n_127026597)
		, .D(n_5758), .Z(n_245380944));
	notech_ao4 i_124064945(.A(n_126126588), .B(n_32089), .C(n_125926586), .D
		(n_33467), .Z(n_245580946));
	notech_and4 i_124464941(.A(n_245580946), .B(n_245380944), .C(n_225980760
		), .D(n_226280763), .Z(n_245780948));
	notech_ao4 i_116665013(.A(n_31482), .B(n_378464315), .C(n_61103), .D(n_30787
		), .Z(n_245880949));
	notech_ao4 i_116565014(.A(n_378764318), .B(nbus_11273[9]), .C(n_327060898
		), .D(n_378564316), .Z(n_245980950));
	notech_ao4 i_116365016(.A(n_378964320), .B(n_33168), .C(n_378664317), .D
		(\nbus_11290[9] ), .Z(n_246180952));
	notech_ao4 i_116265017(.A(n_327160899), .B(n_26394), .C(n_99942440), .D(n_378864319
		), .Z(n_246280953));
	notech_and4 i_116865011(.A(n_246280953), .B(n_246180952), .C(n_245980950
		), .D(n_245880949), .Z(n_246480955));
	notech_ao4 i_115965020(.A(n_327360901), .B(n_26397), .C(n_327260900), .D
		(n_26396), .Z(n_246580956));
	notech_ao4 i_115865021(.A(n_336660994), .B(n_331560943), .C(n_26600), .D
		(n_31517), .Z(n_246680957));
	notech_ao4 i_115665023(.A(n_126126588), .B(n_32068), .C(n_125926586), .D
		(n_33468), .Z(n_246880959));
	notech_and4 i_116165018(.A(n_246880959), .B(n_246680957), .C(n_246580956
		), .D(n_224480745), .Z(n_247180961));
	notech_and2 i_49363350(.A(n_264881138), .B(n_264781137), .Z(n_30339));
	notech_mux2 i_13963220(.S(n_32259), .A(n_247680966), .B(n_247480964), .Z
		(n_247280962));
	notech_ao4 i_10163256(.A(n_29891), .B(n_30920), .C(n_60177), .D(\nbus_11290[1] 
		), .Z(n_247480964));
	notech_ao4 i_10063257(.A(n_30919), .B(n_29891), .C(n_60177), .D(nbus_11273
		[1]), .Z(n_247680966));
	notech_nao3 i_93562457(.A(n_57679), .B(n_32323), .C(n_32321), .Z(n_247980969
		));
	notech_or2 i_23063129(.A(n_25094), .B(nbus_11271[9]), .Z(n_250880998));
	notech_or2 i_22563134(.A(n_23747), .B(n_33168), .Z(n_251581005));
	notech_or2 i_37262995(.A(n_336660994), .B(n_24716), .Z(n_252281012));
	notech_or2 i_36563002(.A(n_381464345), .B(n_33168), .Z(n_252981019));
	notech_or4 i_48962888(.A(n_63718), .B(n_57438), .C(n_63794), .D(nbus_11273
		[5]), .Z(n_253881028));
	notech_or2 i_48662891(.A(n_334860976), .B(n_57036), .Z(n_254181031));
	notech_nao3 i_51762864(.A(n_63790), .B(opc[7]), .C(n_151069548), .Z(n_255081040
		));
	notech_or4 i_51462867(.A(n_63718), .B(n_57438), .C(n_63762), .D(nbus_11273
		[7]), .Z(n_255381043));
	notech_ao3 i_53062852(.A(opa[9]), .B(n_30351), .C(n_60189), .Z(n_255881048
		));
	notech_nao3 i_52962853(.A(n_63768), .B(opc[9]), .C(n_333778343), .Z(n_256181051
		));
	notech_nor2 i_52662856(.A(n_99942440), .B(n_323778246), .Z(n_256481054)
		);
	notech_nor2 i_52362859(.A(n_327060898), .B(n_57393), .Z(n_256781057));
	notech_or2 i_73462649(.A(n_31122), .B(n_140076466), .Z(n_257681066));
	notech_or4 i_77062613(.A(n_63718), .B(n_378364314), .C(n_63756), .D(nbus_11273
		[5]), .Z(n_258981079));
	notech_or4 i_79362590(.A(n_232463321), .B(n_32259), .C(n_29758), .D(nbus_11273
		[1]), .Z(n_259881088));
	notech_or4 i_79062593(.A(n_232463321), .B(n_29758), .C(n_57494), .D(\nbus_11290[1] 
		), .Z(n_260181091));
	notech_or4 i_78762596(.A(n_29891), .B(n_94542386), .C(n_60189), .D(nbus_11273
		[1]), .Z(n_260481094));
	notech_or4 i_83762552(.A(n_61056), .B(n_57494), .C(n_376564296), .D(\nbus_11290[5] 
		), .Z(n_260981099));
	notech_or4 i_83462555(.A(n_63718), .B(n_94542386), .C(n_63758), .D(nbus_11273
		[5]), .Z(n_261281102));
	notech_nao3 i_87362517(.A(n_63790), .B(opc[5]), .C(n_29994), .Z(n_262181111
		));
	notech_or2 i_87062520(.A(n_31122), .B(n_30001), .Z(n_262481114));
	notech_nao3 i_90962482(.A(n_63774), .B(opc[5]), .C(n_30391), .Z(n_263381123
		));
	notech_or4 i_90662485(.A(n_60177), .B(n_303944473), .C(nbus_11273[5]), .D
		(n_32266), .Z(n_263681126));
	notech_nao3 i_5163306(.A(n_32323), .B(n_32310), .C(n_334960977), .Z(n_30338
		));
	notech_or2 i_93262460(.A(n_30379), .B(n_334860976), .Z(n_264581135));
	notech_ao4 i_170661709(.A(n_30373), .B(\nbus_11290[5] ), .C(n_61675), .D
		(n_31513), .Z(n_264681136));
	notech_and2 i_170761708(.A(n_264681136), .B(n_264581135), .Z(n_264781137
		));
	notech_ao4 i_170561710(.A(n_30378), .B(nbus_11273[5]), .C(n_30376), .D(n_33135
		), .Z(n_264881138));
	notech_ao4 i_166861747(.A(n_334860976), .B(n_323860866), .C(n_57170), .D
		(n_30338), .Z(n_264981139));
	notech_ao4 i_166761748(.A(n_31478), .B(n_305344487), .C(n_323960867), .D
		(n_33135), .Z(n_265081140));
	notech_ao4 i_166561750(.A(n_31099), .B(n_30578), .C(n_31098), .D(n_303944473
		), .Z(n_265281142));
	notech_and4 i_167061745(.A(n_265281142), .B(n_265081140), .C(n_264981139
		), .D(n_263681126), .Z(n_265481144));
	notech_ao4 i_166261753(.A(n_31123), .B(n_30390), .C(n_31125), .D(n_30387
		), .Z(n_265581145));
	notech_ao4 i_166061755(.A(n_31126), .B(n_30394), .C(n_31119), .D(n_30393
		), .Z(n_265781147));
	notech_and4 i_166461751(.A(n_30339), .B(n_265781147), .C(n_265581145), .D
		(n_263381123), .Z(n_265981149));
	notech_ao4 i_164161774(.A(n_57122), .B(n_30338), .C(n_31099), .D(n_30576
		), .Z(n_266081150));
	notech_ao4 i_164061775(.A(n_30191), .B(n_33135), .C(n_334860976), .D(n_30196
		), .Z(n_266181151));
	notech_ao4 i_163861777(.A(n_31098), .B(n_1532), .C(n_31478), .D(n_305244486
		), .Z(n_266381153));
	notech_and4 i_164361772(.A(n_266381153), .B(n_266181151), .C(n_266081150
		), .D(n_262481114), .Z(n_266581155));
	notech_ao4 i_163561780(.A(n_31123), .B(n_30002), .C(n_31125), .D(n_29998
		), .Z(n_266681156));
	notech_ao4 i_163361782(.A(n_31126), .B(n_29997), .C(n_31119), .D(n_29993
		), .Z(n_266881158));
	notech_and4 i_163761778(.A(n_30339), .B(n_266881158), .C(n_266681156), .D
		(n_262181111), .Z(n_267081160));
	notech_ao4 i_161361802(.A(n_31099), .B(n_376564296), .C(n_31118), .D(n_376764298
		), .Z(n_267181161));
	notech_ao4 i_161261803(.A(n_57141), .B(n_30338), .C(n_31119), .D(n_376664297
		), .Z(n_267281162));
	notech_ao4 i_161061805(.A(n_376964300), .B(n_33135), .C(n_334860976), .D
		(n_376864299), .Z(n_267481164));
	notech_and4 i_161561800(.A(n_267481164), .B(n_267281162), .C(n_267181161
		), .D(n_261281102), .Z(n_267681166));
	notech_ao4 i_160761808(.A(n_31122), .B(n_29680), .C(n_54741988), .D(n_31478
		), .Z(n_267781167));
	notech_ao4 i_160561810(.A(n_31126), .B(n_29681), .C(n_31123), .D(n_29678
		), .Z(n_267981169));
	notech_and4 i_160961806(.A(n_30339), .B(n_267981169), .C(n_267781167), .D
		(n_260981099), .Z(n_268181171));
	notech_ao4 i_154861867(.A(n_376764298), .B(n_30914), .C(n_247280962), .D
		(n_29888), .Z(n_268281172));
	notech_ao4 i_154661869(.A(n_57141), .B(n_30280), .C(n_376664297), .D(n_30916
		), .Z(n_268481174));
	notech_and4 i_155061865(.A(n_260181091), .B(n_268481174), .C(n_268281172
		), .D(n_260481094), .Z(n_268681176));
	notech_ao4 i_154361872(.A(n_376964300), .B(n_33103), .C(n_376864299), .D
		(n_334360971), .Z(n_268781177));
	notech_ao4 i_154161874(.A(n_54741988), .B(n_31473), .C(n_94542386), .D(n_30891
		), .Z(n_268981179));
	notech_and4 i_154561870(.A(n_30274), .B(n_268981179), .C(n_268781177), .D
		(n_259881088), .Z(n_269181181));
	notech_ao4 i_152961884(.A(n_57064), .B(n_30338), .C(n_31099), .D(n_29342
		), .Z(n_269281182));
	notech_ao4 i_152861885(.A(n_334860976), .B(n_29540), .C(n_29533), .D(\nbus_11290[5] 
		), .Z(n_269381183));
	notech_ao4 i_152661887(.A(n_386464395), .B(n_31478), .C(n_29550), .D(n_33135
		), .Z(n_269581185));
	notech_and4 i_153161882(.A(n_269581185), .B(n_269381183), .C(n_269281182
		), .D(n_258981079), .Z(n_269781187));
	notech_ao4 i_152361890(.A(n_31125), .B(n_29340), .C(n_31122), .D(n_29337
		), .Z(n_269881188));
	notech_ao4 i_152261891(.A(n_31118), .B(n_29333), .C(n_31123), .D(n_29338
		), .Z(n_269981189));
	notech_ao4 i_152061893(.A(n_31126), .B(n_29341), .C(n_31119), .D(n_29334
		), .Z(n_270181191));
	notech_and4 i_152561888(.A(n_30339), .B(n_270181191), .C(n_269981189), .D
		(n_269881188), .Z(n_270381193));
	notech_ao4 i_150061913(.A(n_57604), .B(n_30338), .C(n_31099), .D(n_169676762
		), .Z(n_270481194));
	notech_ao4 i_149961914(.A(n_33135), .B(n_192676984), .C(n_334860976), .D
		(n_323278241), .Z(n_270581195));
	notech_ao4 i_149761916(.A(n_31098), .B(n_57666), .C(n_58044), .D(n_31478
		), .Z(n_270781197));
	notech_and4 i_150261911(.A(n_270781197), .B(n_270581195), .C(n_270481194
		), .D(n_257681066), .Z(n_270981199));
	notech_ao4 i_149461919(.A(n_31123), .B(n_140176467), .C(n_31125), .D(n_139876464
		), .Z(n_271081200));
	notech_ao4 i_149361920(.A(n_31119), .B(n_200377059), .C(n_31118), .D(n_200477060
		), .Z(n_271181201));
	notech_ao4 i_149161922(.A(n_279977810), .B(nbus_11271[5]), .C(n_31126), 
		.D(n_139976465), .Z(n_271381203));
	notech_and4 i_149661917(.A(n_30339), .B(n_271381203), .C(n_271181201), .D
		(n_271081200), .Z(n_271581205));
	notech_ao4 i_128662125(.A(n_326960897), .B(n_57068), .C(n_58030), .D(n_31482
		), .Z(n_271781206));
	notech_ao4 i_128462127(.A(n_57243), .B(nbus_11273[9]), .C(n_57244), .D(\nbus_11290[9] 
		), .Z(n_271981208));
	notech_or4 i_128862123(.A(n_256781057), .B(n_256481054), .C(n_30353), .D
		(n_30352), .Z(n_272181210));
	notech_ao4 i_128162130(.A(n_327260900), .B(n_333978345), .C(n_323978248)
		, .D(n_33168), .Z(n_272281211));
	notech_nand2 i_128262129(.A(n_272281211), .B(n_256181051), .Z(n_272781212
		));
	notech_ao4 i_127662134(.A(n_324360871), .B(n_143669474), .C(n_324460872)
		, .D(n_143369471), .Z(n_273081215));
	notech_ao4 i_127562135(.A(n_324260870), .B(n_143469472), .C(n_324760875)
		, .D(n_143569473), .Z(n_273181216));
	notech_ao4 i_127362137(.A(n_5783), .B(n_31480), .C(n_324160869), .D(n_143769475
		), .Z(n_273981218));
	notech_and4 i_127862132(.A(n_255381043), .B(n_273981218), .C(n_273181216
		), .D(n_273081215), .Z(n_274181220));
	notech_ao4 i_127062140(.A(n_100242443), .B(n_57036), .C(n_57027), .D(n_33165
		), .Z(n_274281221));
	notech_ao4 i_126862142(.A(n_323760865), .B(n_57068), .C(n_150969547), .D
		(n_324660874), .Z(n_274481223));
	notech_and4 i_127262138(.A(n_324860876), .B(n_274481223), .C(n_274281221
		), .D(n_255081040), .Z(n_274781225));
	notech_ao4 i_125162157(.A(n_31125), .B(n_143669474), .C(n_31123), .D(n_143369471
		), .Z(n_274881226));
	notech_ao4 i_125062158(.A(n_31122), .B(n_143469472), .C(n_31126), .D(n_143569473
		), .Z(n_274981227));
	notech_ao4 i_124862160(.A(n_31099), .B(n_143769475), .C(n_57068), .D(n_30338
		), .Z(n_275181229));
	notech_and4 i_125362155(.A(n_275181229), .B(n_274981227), .C(n_274881226
		), .D(n_254181031), .Z(n_275381231));
	notech_ao4 i_124562163(.A(n_5783), .B(n_31478), .C(n_57027), .D(n_33135)
		, .Z(n_275481232));
	notech_ao4 i_124362165(.A(n_31119), .B(n_150969547), .C(n_31118), .D(n_151069548
		), .Z(n_275681234));
	notech_and4 i_124762161(.A(n_30339), .B(n_275681234), .C(n_275481232), .D
		(n_253881028), .Z(n_275881236));
	notech_ao4 i_114562256(.A(n_31482), .B(n_381264343), .C(n_61103), .D(n_30766
		), .Z(n_275981237));
	notech_ao4 i_114462257(.A(n_381664347), .B(\nbus_11290[9] ), .C(n_327060898
		), .D(n_381564346), .Z(n_276081238));
	notech_ao4 i_114262259(.A(n_99942440), .B(n_381364344), .C(n_381764348),
		 .D(nbus_11273[9]), .Z(n_276281240));
	notech_and4 i_114762254(.A(n_276281240), .B(n_276081238), .C(n_275981237
		), .D(n_252981019), .Z(n_276481242));
	notech_ao4 i_113962262(.A(n_327160899), .B(n_24541), .C(n_327260900), .D
		(n_24539), .Z(n_276581243));
	notech_ao4 i_113862263(.A(n_60453), .B(n_31517), .C(n_327360901), .D(n_24542
		), .Z(n_276681244));
	notech_ao4 i_113662265(.A(n_24528), .B(n_33470), .C(n_24527), .D(n_33469
		), .Z(n_276881246));
	notech_and4 i_114162260(.A(n_276881246), .B(n_276681244), .C(n_276581243
		), .D(n_252281012), .Z(n_277081248));
	notech_ao4 i_101662380(.A(n_326960897), .B(n_58702), .C(n_31482), .D(n_386264393
		), .Z(n_277181249));
	notech_ao4 i_101562381(.A(n_386164392), .B(\nbus_11290[9] ), .C(n_327060898
		), .D(n_386364394), .Z(n_277281250));
	notech_ao4 i_101362383(.A(n_99942440), .B(n_23750), .C(nbus_11273[9]), .D
		(n_386064391), .Z(n_277481252));
	notech_and4 i_101862378(.A(n_277481252), .B(n_277281250), .C(n_277181249
		), .D(n_251581005), .Z(n_277681254));
	notech_ao4 i_101062386(.A(n_327160899), .B(n_23613), .C(n_327260900), .D
		(n_23611), .Z(n_277781255));
	notech_ao4 i_100962387(.A(n_56036), .B(n_32538), .C(n_327360901), .D(n_23614
		), .Z(n_277881256));
	notech_ao3 i_100762388(.A(n_327460902), .B(n_250880998), .C(n_335060978)
		, .Z(n_278181259));
	notech_ao4 i_100362392(.A(n_334560973), .B(n_324060868), .C(n_334460972)
		, .D(n_31480), .Z(n_278381261));
	notech_ao4 i_100262393(.A(n_391164442), .B(n_100242443), .C(n_391264443)
		, .D(n_33165), .Z(n_278481262));
	notech_ao4 i_100062395(.A(n_23510), .B(n_324560873), .C(n_23519), .D(n_324160869
		), .Z(n_278681264));
	notech_ao4 i_99962396(.A(n_23517), .B(n_324760875), .C(n_23511), .D(n_324660874
		), .Z(n_278781265));
	notech_and4 i_100562390(.A(n_278781265), .B(n_278681264), .C(n_278481262
		), .D(n_278381261), .Z(n_278981267));
	notech_ao4 i_99562399(.A(n_23514), .B(n_324260870), .C(n_23518), .D(n_324360871
		), .Z(n_279081268));
	notech_ao4 i_99462400(.A(n_58702), .B(n_323760865), .C(n_23515), .D(n_324460872
		), .Z(n_279181269));
	notech_ao4 i_99262402(.A(n_25094), .B(nbus_11271[7]), .C(n_56036), .D(n_32535
		), .Z(n_279381271));
	notech_and4 i_99862397(.A(n_324860876), .B(n_279381271), .C(n_279181269)
		, .D(n_279081268), .Z(n_279581273));
	notech_ao4 i_97662418(.A(n_391164442), .B(n_334860976), .C(n_58702), .D(n_30338
		), .Z(n_279681274));
	notech_ao4 i_97562419(.A(n_334460972), .B(n_56983), .C(n_391264443), .D(n_33135
		), .Z(n_279781275));
	notech_ao4 i_97262421(.A(n_23519), .B(n_31099), .C(n_334560973), .D(n_31098
		), .Z(n_279981277));
	notech_ao4 i_97162422(.A(n_31125), .B(n_23518), .C(n_31122), .D(n_23514)
		, .Z(n_280081278));
	notech_and4 i_97862416(.A(n_280081278), .B(n_279981277), .C(n_279781275)
		, .D(n_279681274), .Z(n_280281280));
	notech_ao4 i_96762425(.A(n_23510), .B(n_31118), .C(n_23515), .D(n_31123)
		, .Z(n_280381281));
	notech_ao4 i_96662426(.A(n_23517), .B(n_31126), .C(n_23511), .D(n_31119)
		, .Z(n_280481282));
	notech_ao4 i_96462428(.A(n_56036), .B(n_32533), .C(n_25094), .D(nbus_11271
		[5]), .Z(n_280681284));
	notech_and4 i_97062423(.A(n_30339), .B(n_280681284), .C(n_280481282), .D
		(n_280381281), .Z(n_280881286));
	notech_or2 i_171860649(.A(n_334560973), .B(n_32249), .Z(n_23514));
	notech_or4 i_171960648(.A(n_32275), .B(n_334560973), .C(instrc[122]), .D
		(instrc[120]), .Z(n_23515));
	notech_nao3 i_174160643(.A(n_23763), .B(n_58566), .C(n_334560973), .Z(n_23517
		));
	notech_or4 i_174460642(.A(n_32275), .B(n_23519), .C(instrc[122]), .D(instrc
		[120]), .Z(n_23518));
	notech_or4 i_35160314(.A(n_336660994), .B(n_30719), .C(n_340461032), .D(n_2830
		), .Z(n_286581343));
	notech_nand2 i_35060315(.A(opd[9]), .B(n_30354), .Z(n_286881346));
	notech_or2 i_34760318(.A(n_441768001), .B(nbus_11273[9]), .Z(n_287181349
		));
	notech_nao3 i_58060123(.A(n_63790), .B(opc[5]), .C(n_200977065), .Z(n_287881356
		));
	notech_nor2 i_58360120(.A(n_324760875), .B(n_178576845), .Z(n_290781385)
		);
	notech_ao4 i_142759320(.A(n_324260870), .B(n_178676846), .C(n_178776847)
		, .D(n_324460872), .Z(n_290881386));
	notech_ao4 i_142659321(.A(n_324160869), .B(n_178376843), .C(n_324360871)
		, .D(n_178476844), .Z(n_291081388));
	notech_ao3 i_142959318(.A(n_290881386), .B(n_291081388), .C(n_290781385)
		, .Z(n_291181389));
	notech_ao4 i_142459323(.A(nbus_11273[7]), .B(n_30401), .C(n_323760865), 
		.D(n_57147), .Z(n_291281390));
	notech_ao4 i_142359324(.A(n_56783), .B(n_31515), .C(n_197877035), .D(\nbus_11290[7] 
		), .Z(n_291381391));
	notech_ao4 i_142059327(.A(n_204977105), .B(n_33165), .C(n_100242443), .D
		(n_57289), .Z(n_291681394));
	notech_ao4 i_141859328(.A(n_324060868), .B(n_57432), .C(n_58019), .D(n_31480
		), .Z(n_291781395));
	notech_ao4 i_141659330(.A(n_324660874), .B(n_200877064), .C(n_57426), .D
		(n_4448), .Z(n_291981397));
	notech_ao4 i_141559331(.A(n_56896), .B(n_30943), .C(n_324560873), .D(n_200977065
		), .Z(n_292081398));
	notech_and4 i_142259325(.A(n_292081398), .B(n_291981397), .C(n_291781395
		), .D(n_291681394), .Z(n_292281400));
	notech_ao4 i_141259334(.A(n_31123), .B(n_178776847), .C(n_31513), .D(n_178876848
		), .Z(n_292381401));
	notech_ao4 i_141159335(.A(n_31126), .B(n_178576845), .C(n_31122), .D(n_178676846
		), .Z(n_292481402));
	notech_ao4 i_140959337(.A(n_31099), .B(n_178376843), .C(n_31125), .D(n_178476844
		), .Z(n_292681404));
	notech_ao4 i_140859338(.A(nbus_11273[5]), .B(n_30322), .C(n_57010), .D(n_33135
		), .Z(n_292781405));
	notech_and4 i_141459332(.A(n_292781405), .B(n_292681404), .C(n_292481402
		), .D(n_292381401), .Z(n_292981407));
	notech_ao4 i_140559341(.A(n_58019), .B(n_56983), .C(\nbus_11290[5] ), .D
		(n_197877035), .Z(n_293081408));
	notech_ao4 i_140459342(.A(n_57432), .B(n_31098), .C(n_57147), .D(n_30338
		), .Z(n_293181409));
	notech_ao4 i_140259344(.A(n_31119), .B(n_200877064), .C(n_334860976), .D
		(n_57289), .Z(n_293381411));
	notech_and4 i_140759339(.A(n_293381411), .B(n_293181409), .C(n_293081408
		), .D(n_287881356), .Z(n_293581413));
	notech_ao4 i_108159630(.A(n_385664387), .B(n_33168), .C(n_99942440), .D(n_385864389
		), .Z(n_293681414));
	notech_ao4 i_107959631(.A(n_56036), .B(n_32561), .C(n_327260900), .D(n_385464385
		), .Z(n_293781415));
	notech_ao4 i_107659633(.A(n_327060898), .B(n_440667990), .C(n_441668000)
		, .D(\nbus_11290[9] ), .Z(n_293981417));
	notech_and4 i_108359628(.A(n_293981417), .B(n_293781415), .C(n_293681414
		), .D(n_287181349), .Z(n_294181419));
	notech_ao4 i_107359636(.A(n_327160899), .B(n_441868002), .C(n_327360901)
		, .D(n_4533), .Z(n_294281420));
	notech_ao3 i_107259637(.A(n_286581343), .B(n_55802), .C(n_30917), .Z(n_294581423
		));
	notech_ao4 i_106859641(.A(n_179484224), .B(n_324760875), .C(n_179584225)
		, .D(n_324360871), .Z(n_294781425));
	notech_ao4 i_106659642(.A(n_179284222), .B(n_324260870), .C(n_179384223)
		, .D(n_324460872), .Z(n_294881426));
	notech_ao4 i_106459644(.A(n_56036), .B(n_32559), .C(n_323760865), .D(n_30590
		), .Z(n_295081428));
	notech_ao4 i_106359645(.A(n_382864359), .B(n_33165), .C(n_383064361), .D
		(n_324660874), .Z(n_295181429));
	notech_and4 i_107059639(.A(n_295181429), .B(n_295081428), .C(n_294881426
		), .D(n_294781425), .Z(n_295381431));
	notech_ao4 i_106059648(.A(n_57260), .B(n_324560873), .C(n_382664357), .D
		(n_100242443), .Z(n_295481432));
	notech_ao4 i_105959649(.A(n_188084307), .B(n_324160869), .C(n_57383), .D
		(n_324060868), .Z(n_295581433));
	notech_ao4 i_105759651(.A(n_25094), .B(\nbus_11290[7] ), .C(n_58051), .D
		(n_31480), .Z(n_295781435));
	notech_and4 i_106259646(.A(n_324860876), .B(n_295781435), .C(n_295581433
		), .D(n_295481432), .Z(n_295981437));
	notech_ao4 i_103859668(.A(n_31126), .B(n_179484224), .C(n_31125), .D(n_179584225
		), .Z(n_296081438));
	notech_ao4 i_103759669(.A(n_179284222), .B(n_31122), .C(n_31123), .D(n_179384223
		), .Z(n_296181439));
	notech_ao4 i_103559671(.A(n_383064361), .B(n_31119), .C(n_56036), .D(n_32557
		), .Z(n_296381441));
	notech_ao4 i_103459672(.A(n_382664357), .B(n_334860976), .C(n_382864359)
		, .D(n_33135), .Z(n_296481442));
	notech_and4 i_104059666(.A(n_296481442), .B(n_296381441), .C(n_296181439
		), .D(n_296081438), .Z(n_296681444));
	notech_ao4 i_103159675(.A(n_57383), .B(n_31098), .C(n_57260), .D(n_31118
		), .Z(n_296781445));
	notech_ao4 i_103059676(.A(n_58051), .B(n_56983), .C(n_188084307), .D(n_31099
		), .Z(n_296881446));
	notech_ao4 i_102859678(.A(n_25094), .B(\nbus_11290[5] ), .C(n_30590), .D
		(n_30338), .Z(n_297081448));
	notech_and4 i_102959677(.A(n_264881138), .B(n_55802), .C(n_297081448), .D
		(n_264781137), .Z(n_297281450));
	notech_ao4 i_84859857(.A(n_23517), .B(n_31075), .C(n_23518), .D(n_31074)
		, .Z(n_297481452));
	notech_ao4 i_84759858(.A(n_23514), .B(n_31071), .C(n_23515), .D(n_31072)
		, .Z(n_297581453));
	notech_ao4 i_84559860(.A(n_58702), .B(n_187176929), .C(n_31048), .D(n_23519
		), .Z(n_297781455));
	notech_ao4 i_84459861(.A(n_391264443), .B(n_33104), .C(n_56036), .D(n_32532
		), .Z(n_297881456));
	notech_and4 i_85059855(.A(n_297881456), .B(n_297781455), .C(n_297581453)
		, .D(n_297481452), .Z(n_298081458));
	notech_ao4 i_84159864(.A(n_334460972), .B(n_31477), .C(n_391164442), .D(n_334660974
		), .Z(n_298181459));
	notech_ao4 i_84059865(.A(n_23510), .B(n_31067), .C(n_334560973), .D(n_31047
		), .Z(n_298281460));
	notech_ao4 i_83859867(.A(n_25094), .B(nbus_11271[4]), .C(n_23511), .D(n_31068
		), .Z(n_298481462));
	notech_ao3 i_83959866(.A(n_298481462), .B(n_187576933), .C(n_335060978),
		 .Z(n_298681464));
	notech_ao4 i_83459871(.A(n_326460892), .B(n_23517), .C(n_23518), .D(n_326560893
		), .Z(n_298881466));
	notech_ao4 i_83359872(.A(n_23514), .B(n_326660894), .C(n_23515), .D(n_326760895
		), .Z(n_298981467));
	notech_ao4 i_83159874(.A(n_326060888), .B(n_58702), .C(n_23519), .D(n_325960887
		), .Z(n_299181469));
	notech_ao4 i_83059875(.A(n_391264443), .B(n_33167), .C(n_56036), .D(n_32530
		), .Z(n_299281470));
	notech_and4 i_83659869(.A(n_299281470), .B(n_299181469), .C(n_298981467)
		, .D(n_298881466), .Z(n_299481472));
	notech_ao4 i_82759878(.A(n_25094), .B(nbus_11271[2]), .C(n_391164442), .D
		(n_100842449), .Z(n_299581473));
	notech_ao4 i_82659879(.A(n_334560973), .B(n_326160889), .C(n_334460972),
		 .D(n_31474), .Z(n_299681474));
	notech_ao4 i_82459881(.A(n_23511), .B(n_326260890), .C(n_23510), .D(n_326360891
		), .Z(n_299881476));
	notech_ao3 i_82559880(.A(n_299881476), .B(n_326860896), .C(n_335060978),
		 .Z(n_300081478));
	notech_nand2 i_16655782(.A(tsc[29]), .B(n_30615), .Z(n_300481482));
	notech_or2 i_16555783(.A(n_131426641), .B(nbus_11271[29]), .Z(n_300781485
		));
	notech_nao3 i_16055788(.A(n_57397), .B(opd[29]), .C(n_58702), .Z(n_301281490
		));
	notech_or2 i_24555703(.A(n_25110), .B(nbus_11271[29]), .Z(n_301681494)
		);
	notech_nand3 i_24055708(.A(n_57397), .B(n_32219), .C(opd[29]), .Z(n_302181499
		));
	notech_or2 i_29855657(.A(n_26585), .B(n_31020), .Z(n_302481502));
	notech_or2 i_29555660(.A(n_337761005), .B(nbus_11271[26]), .Z(n_302781505
		));
	notech_or2 i_29255663(.A(n_127026597), .B(n_5720), .Z(n_303081508));
	notech_or2 i_31155644(.A(n_26585), .B(n_31022), .Z(n_303781515));
	notech_or2 i_30855647(.A(n_337761005), .B(nbus_11271[27]), .Z(n_304081518
		));
	notech_or2 i_30555650(.A(n_127026597), .B(n_5711), .Z(n_304381521));
	notech_or2 i_32455631(.A(n_26585), .B(n_31024), .Z(n_305081528));
	notech_or2 i_32155634(.A(n_337761005), .B(nbus_11271[28]), .Z(n_305381531
		));
	notech_or2 i_31855637(.A(n_4427), .B(n_127026597), .Z(n_305681534));
	notech_or2 i_33755618(.A(n_26585), .B(n_31026), .Z(n_306381541));
	notech_or2 i_33455621(.A(n_337761005), .B(nbus_11271[29]), .Z(n_306681544
		));
	notech_or2 i_33155624(.A(n_4428), .B(n_127026597), .Z(n_306981547));
	notech_nand3 i_58755379(.A(n_164196010), .B(n_171160315), .C(n_1765), .Z
		(n_307681554));
	notech_or2 i_58455382(.A(n_122726554), .B(\nbus_11283[29] ), .Z(n_307981557
		));
	notech_or2 i_58155385(.A(n_122826555), .B(n_33197), .Z(n_308281560));
	notech_nand2 i_57855388(.A(sav_edi[29]), .B(n_61871), .Z(n_308581563));
	notech_or2 i_61955347(.A(n_28867), .B(nbus_11271[29]), .Z(n_308681564)
		);
	notech_nao3 i_61455352(.A(n_57397), .B(opd[29]), .C(n_57195), .Z(n_309381571
		));
	notech_nand3 i_70255264(.A(n_57397), .B(n_32211), .C(opd[29]), .Z(n_310181579
		));
	notech_or2 i_73955227(.A(n_443668020), .B(nbus_11271[29]), .Z(n_310281580
		));
	notech_nand3 i_73455232(.A(n_57395), .B(n_32224), .C(opd[29]), .Z(n_310981587
		));
	notech_or2 i_77155195(.A(n_443168015), .B(nbus_11271[29]), .Z(n_311081588
		));
	notech_nand3 i_76655200(.A(n_57395), .B(n_125342694), .C(opd[29]), .Z(n_311781595
		));
	notech_nand3 i_84355129(.A(n_57395), .B(n_32220), .C(opd[29]), .Z(n_311981596
		));
	notech_nao3 i_83855134(.A(n_63790), .B(opc_10[29]), .C(n_442768011), .Z(n_312681603
		));
	notech_nand2 i_2055922(.A(n_63790), .B(opc_10[29]), .Z(n_94229643));
	notech_ao4 i_181854179(.A(n_31672), .B(n_57230), .C(n_57103), .D(n_31601
		), .Z(n_315981636));
	notech_ao4 i_181754180(.A(n_59100), .B(n_31928), .C(n_31437), .D(n_57218
		), .Z(n_316081637));
	notech_ao4 i_181554182(.A(n_31896), .B(n_57091), .C(n_58702), .D(n_31993
		), .Z(n_316281639));
	notech_ao4 i_181454183(.A(n_31704), .B(n_57064), .C(n_57068), .D(n_31832
		), .Z(n_316381640));
	notech_and4 i_182054177(.A(n_316381640), .B(n_316281639), .C(n_316081637
		), .D(n_315981636), .Z(n_316581642));
	notech_ao4 i_181154186(.A(n_57195), .B(n_31736), .C(n_30679), .D(n_31961
		), .Z(n_316681643));
	notech_ao4 i_181054187(.A(n_31864), .B(n_57170), .C(n_32025), .D(n_30590
		), .Z(n_316781644));
	notech_and2 i_181254185(.A(n_316781644), .B(n_316681643), .Z(n_316881645
		));
	notech_ao4 i_180854189(.A(n_31768), .B(n_57141), .C(n_57147), .D(n_33489
		), .Z(n_316981646));
	notech_ao4 i_180754190(.A(n_57122), .B(n_31800), .C(n_33488), .D(n_57604
		), .Z(n_317081647));
	notech_nand2 i_1955923(.A(n_63790), .B(opc_10[28]), .Z(n_7636));
	notech_ao4 i_179454203(.A(n_57218), .B(n_31436), .C(n_57230), .D(n_31671
		), .Z(n_317381650));
	notech_ao4 i_179354204(.A(n_58702), .B(n_31992), .C(n_59100), .D(n_31927
		), .Z(n_317481651));
	notech_ao4 i_179154206(.A(n_57091), .B(n_31895), .C(n_57097), .D(n_31600
		), .Z(n_317681653));
	notech_ao4 i_179054207(.A(n_57064), .B(n_31703), .C(n_57068), .D(n_31831
		), .Z(n_317781654));
	notech_and4 i_179654201(.A(n_317781654), .B(n_317681653), .C(n_317481651
		), .D(n_317381650), .Z(n_317981656));
	notech_ao4 i_178754210(.A(n_57195), .B(n_31735), .C(n_30679), .D(n_31960
		), .Z(n_318081657));
	notech_ao4 i_178654211(.A(n_57170), .B(n_31863), .C(n_30590), .D(n_32024
		), .Z(n_318181658));
	notech_and2 i_178854209(.A(n_318181658), .B(n_318081657), .Z(n_318281659
		));
	notech_ao4 i_178454213(.A(n_57141), .B(n_31767), .C(n_57147), .D(n_33487
		), .Z(n_318381660));
	notech_ao4 i_178354214(.A(n_57122), .B(n_31799), .C(n_57604), .D(n_33486
		), .Z(n_318481661));
	notech_ao4 i_171854278(.A(n_442868012), .B(n_60620), .C(n_442968013), .D
		(n_4387), .Z(n_318781664));
	notech_ao4 i_171754279(.A(n_442568009), .B(\nbus_11290[29] ), .C(n_442668010
		), .D(\nbus_11283[29] ), .Z(n_318981666));
	notech_and3 i_172054276(.A(n_318781664), .B(n_318981666), .C(n_312681603
		), .Z(n_319081667));
	notech_ao4 i_171554281(.A(n_117626503), .B(n_33197), .C(n_4428), .D(n_117726504
		), .Z(n_319181668));
	notech_ao4 i_162054372(.A(n_4387), .B(n_443468018), .C(n_443568019), .D(n_94229643
		), .Z(n_319481671));
	notech_ao4 i_161954373(.A(n_4428), .B(n_118526512), .C(n_118426511), .D(n_33197
		), .Z(n_319681673));
	notech_and3 i_162254370(.A(n_319481671), .B(n_319681673), .C(n_311781595
		), .Z(n_319781674));
	notech_ao4 i_161754375(.A(n_443268016), .B(\nbus_11283[29] ), .C(n_443368017
		), .D(\nbus_11290[29] ), .Z(n_319881675));
	notech_ao4 i_159254400(.A(n_4387), .B(n_443968023), .C(n_94229643), .D(n_444068024
		), .Z(n_320181678));
	notech_ao4 i_159154401(.A(n_4428), .B(n_119326520), .C(n_119226519), .D(n_33197
		), .Z(n_320381680));
	notech_and3 i_159454398(.A(n_320181678), .B(n_320381680), .C(n_310981587
		), .Z(n_320481681));
	notech_ao4 i_158954403(.A(n_443768021), .B(\nbus_11283[29] ), .C(n_443868022
		), .D(\nbus_11290[29] ), .Z(n_320581682));
	notech_ao4 i_155854434(.A(n_4387), .B(n_303822063), .C(n_94229643), .D(n_299122016
		), .Z(n_320881685));
	notech_ao4 i_155754435(.A(n_4428), .B(n_57320), .C(n_57319), .D(n_33197)
		, .Z(n_321081687));
	notech_and3 i_156054432(.A(n_320881685), .B(n_321081687), .C(n_310181579
		), .Z(n_321181688));
	notech_ao4 i_155554437(.A(n_57363), .B(n_58474), .C(n_57362), .D(n_58947
		), .Z(n_321281689));
	notech_ao4 i_155454438(.A(n_303922064), .B(n_60620), .C(n_31537), .D(n_61675
		), .Z(n_321381690));
	notech_ao4 i_144254548(.A(n_4387), .B(n_28852), .C(n_94229643), .D(n_28869
		), .Z(n_321581692));
	notech_ao4 i_144154549(.A(n_4428), .B(n_388264413), .C(n_388364414), .D(n_33197
		), .Z(n_321781694));
	notech_and3 i_144454546(.A(n_321581692), .B(n_321781694), .C(n_309381571
		), .Z(n_321881695));
	notech_ao4 i_143954551(.A(n_28874), .B(n_58474), .C(n_28863), .D(n_58947
		), .Z(n_321981696));
	notech_ao4 i_141454576(.A(n_4387), .B(n_122226549), .C(n_94229643), .D(n_337461002
		), .Z(n_322281699));
	notech_ao4 i_141254578(.A(n_57001), .B(n_31537), .C(n_331060938), .D(n_31505
		), .Z(n_322481701));
	notech_and4 i_141654574(.A(n_322481701), .B(n_322281699), .C(n_308281560
		), .D(n_308581563), .Z(n_322681703));
	notech_ao4 i_140954581(.A(n_122626553), .B(n_58947), .C(n_4428), .D(n_122926556
		), .Z(n_322781704));
	notech_ao4 i_140754583(.A(n_333360961), .B(n_33471), .C(n_337361001), .D
		(n_60620), .Z(n_322981706));
	notech_and4 i_141154579(.A(n_322981706), .B(n_322781704), .C(n_307681554
		), .D(n_307981557), .Z(n_323181708));
	notech_ao4 i_120454786(.A(n_4387), .B(n_126226589), .C(n_337961007), .D(n_94229643
		), .Z(n_323281709));
	notech_ao4 i_120354787(.A(n_337861006), .B(n_31505), .C(n_61103), .D(n_30807
		), .Z(n_323381710));
	notech_ao4 i_120154789(.A(n_126926596), .B(n_33197), .C(n_55946), .D(n_31537
		), .Z(n_323581712));
	notech_and4 i_120654784(.A(n_323581712), .B(n_323381710), .C(n_323281709
		), .D(n_306981547), .Z(n_323781714));
	notech_ao4 i_119854792(.A(n_126726594), .B(n_58474), .C(n_126826595), .D
		(n_58947), .Z(n_323881715));
	notech_ao4 i_119654794(.A(n_126126588), .B(n_32088), .C(n_125926586), .D
		(n_33472), .Z(n_324081717));
	notech_and4 i_120054790(.A(n_324081717), .B(n_323881715), .C(n_306381541
		), .D(n_306681544), .Z(n_324281719));
	notech_ao4 i_119354797(.A(n_126226589), .B(n_440082450), .C(n_337961007)
		, .D(n_7636), .Z(n_324381720));
	notech_ao4 i_119254798(.A(n_337861006), .B(n_31504), .C(n_61104), .D(n_30806
		), .Z(n_324481721));
	notech_ao4 i_119054800(.A(n_126926596), .B(n_33196), .C(n_55946), .D(n_31536
		), .Z(n_324681723));
	notech_and4 i_119554795(.A(n_324681723), .B(n_324481721), .C(n_324381720
		), .D(n_305681534), .Z(n_324881725));
	notech_ao4 i_118754803(.A(n_126726594), .B(\nbus_11283[28] ), .C(n_126826595
		), .D(\nbus_11290[28] ), .Z(n_324981726));
	notech_ao4 i_118554805(.A(n_55975), .B(n_32087), .C(n_55966), .D(n_33473
		), .Z(n_325181728));
	notech_and4 i_118954801(.A(n_325181728), .B(n_305381531), .C(n_324981726
		), .D(n_305081528), .Z(n_325381730));
	notech_ao4 i_118254808(.A(n_126226589), .B(n_284131522), .C(n_337961007)
		, .D(n_172669762), .Z(n_325481731));
	notech_ao4 i_118154809(.A(n_337861006), .B(n_31503), .C(n_61104), .D(n_30805
		), .Z(n_325581732));
	notech_ao4 i_117954811(.A(n_126926596), .B(n_33195), .C(n_55946), .D(n_31535
		), .Z(n_325781734));
	notech_and4 i_118454806(.A(n_325781734), .B(n_325581732), .C(n_325481731
		), .D(n_304381521), .Z(n_325981736));
	notech_ao4 i_117654814(.A(n_126726594), .B(\nbus_11283[27] ), .C(n_126826595
		), .D(\nbus_11290[27] ), .Z(n_326081737));
	notech_ao4 i_117454816(.A(n_55975), .B(n_32086), .C(n_55966), .D(n_33474
		), .Z(n_326281739));
	notech_and4 i_117854812(.A(n_326281739), .B(n_304081518), .C(n_326081737
		), .D(n_303781515), .Z(n_326481741));
	notech_ao4 i_117154819(.A(n_126226589), .B(n_284231523), .C(n_175169787)
		, .D(n_337961007), .Z(n_326581742));
	notech_ao4 i_117054820(.A(n_337861006), .B(n_31502), .C(n_61104), .D(n_30802
		), .Z(n_326681743));
	notech_ao4 i_116854822(.A(n_126926596), .B(n_33198), .C(n_55946), .D(n_31534
		), .Z(n_326881745));
	notech_and4 i_117354817(.A(n_326881745), .B(n_326681743), .C(n_326581742
		), .D(n_303081508), .Z(n_327081747));
	notech_ao4 i_116554825(.A(n_126726594), .B(\nbus_11283[26] ), .C(n_126826595
		), .D(\nbus_11290[26] ), .Z(n_327181748));
	notech_ao4 i_116354827(.A(n_55975), .B(n_32085), .C(n_55966), .D(n_33475
		), .Z(n_327381750));
	notech_and4 i_116754823(.A(n_327381750), .B(n_302781505), .C(n_327181748
		), .D(n_302481502), .Z(n_327581752));
	notech_ao4 i_112754861(.A(n_4387), .B(n_25090), .C(n_94229643), .D(n_365428694
		), .Z(n_327681753));
	notech_ao4 i_112654862(.A(n_4428), .B(n_365328693), .C(n_365228692), .D(n_33197
		), .Z(n_327881755));
	notech_and3 i_112954859(.A(n_327681753), .B(n_327881755), .C(n_302181499
		), .Z(n_327981756));
	notech_ao4 i_112354865(.A(n_365628696), .B(n_58474), .C(n_365528695), .D
		(n_58947), .Z(n_328081757));
	notech_ao4 i_112254866(.A(n_56036), .B(n_32580), .C(n_31537), .D(n_61675
		), .Z(n_328281759));
	notech_ao4 i_105554933(.A(n_4387), .B(n_388064411), .C(n_94229643), .D(n_388164412
		), .Z(n_328481761));
	notech_ao4 i_105454934(.A(n_4428), .B(n_131626643), .C(n_131526642), .D(n_33197
		), .Z(n_328681763));
	notech_ao4 i_105154937(.A(n_387864409), .B(n_58474), .C(n_387964410), .D
		(n_58947), .Z(n_328881765));
	notech_and4 i_105354935(.A(n_222077272), .B(n_328881765), .C(n_300481482
		), .D(n_300781485), .Z(n_329181768));
	notech_ao4 i_35392(.A(n_19698), .B(n_343481901), .C(n_340981876), .D(n_4106
		), .Z(n_329281769));
	notech_or4 i_253065(.A(n_32396), .B(n_28008), .C(\opcode[1] ), .D(n_61940
		), .Z(n_329381770));
	notech_nao3 i_153066(.A(n_30524), .B(n_32548), .C(n_19672), .Z(n_329681773
		));
	notech_nand2 i_33265(.A(n_19603), .B(n_19612), .Z(n_26133));
	notech_nor2 i_2853043(.A(n_343481901), .B(n_19698), .Z(n_329781774));
	notech_and4 i_3853036(.A(n_32590), .B(n_1817), .C(n_2033), .D(n_59515), 
		.Z(n_330081777));
	notech_ao4 i_52131(.A(n_330081777), .B(n_61846), .C(n_340781874), .D(n_3456
		), .Z(n_330181778));
	notech_or4 i_196953086(.A(n_32396), .B(n_28534), .C(n_61846), .D(n_60157
		), .Z(n_330281779));
	notech_or4 i_7253002(.A(n_61892), .B(n_316760795), .C(n_61725), .D(n_61871
		), .Z(n_330381780));
	notech_or4 i_7353001(.A(n_61675), .B(n_415382405), .C(n_340981876), .D(n_61873
		), .Z(n_330481781));
	notech_or4 i_7552999(.A(n_4106), .B(n_340981876), .C(n_61873), .D(n_61675
		), .Z(n_330581782));
	notech_nao3 i_8052994(.A(n_63718), .B(n_61940), .C(n_330881785), .Z(n_330781784
		));
	notech_ao4 i_1853052(.A(n_25681), .B(n_32383), .C(n_32573), .D(n_31160),
		 .Z(n_330881785));
	notech_or4 i_7952995(.A(n_32576), .B(n_28534), .C(\opcode[1] ), .D(n_61940
		), .Z(n_331181788));
	notech_and4 i_4653028(.A(n_331181788), .B(n_341481881), .C(n_341581882),
		 .D(n_330781784), .Z(n_331281789));
	notech_and3 i_4553029(.A(n_25485), .B(n_4025), .C(n_25680), .Z(n_331381790
		));
	notech_or4 i_8652988(.A(n_30304), .B(n_61892), .C(n_57001), .D(n_33242),
		 .Z(n_331481791));
	notech_or4 i_9052985(.A(n_57001), .B(n_30538), .C(n_56755), .D(n_38705),
		 .Z(n_331581792));
	notech_or4 i_8952986(.A(n_61846), .B(n_61940), .C(n_61958), .D(n_331381790
		), .Z(n_331681793));
	notech_or4 i_8852987(.A(n_61725), .B(n_61892), .C(n_331281789), .D(n_61871
		), .Z(n_331781794));
	notech_or2 i_9752978(.A(n_330281779), .B(n_27843), .Z(n_331881795));
	notech_and3 i_50239(.A(n_341381880), .B(n_342481891), .C(n_331881795), .Z
		(n_331981796));
	notech_nand2 i_10152974(.A(n_1806), .B(n_31160), .Z(n_332081797));
	notech_and4 i_11352962(.A(readio_ack), .B(n_4338), .C(n_19663), .D(n_32508
		), .Z(n_332181798));
	notech_and4 i_4453030(.A(n_343181898), .B(n_342981896), .C(n_342881895),
		 .D(n_363850921), .Z(n_332281799));
	notech_and4 i_4353031(.A(n_58597), .B(n_30664), .C(n_58566), .D(n_58555)
		, .Z(n_332381800));
	notech_nor2 i_4253032(.A(n_332181798), .B(n_329781774), .Z(n_332481801)
		);
	notech_or4 i_11752958(.A(n_340561033), .B(n_28534), .C(n_61846), .D(n_332381800
		), .Z(n_332581802));
	notech_nao3 i_11852957(.A(n_61104), .B(n_61632), .C(n_332481801), .Z(n_332681803
		));
	notech_or4 i_11652959(.A(n_61725), .B(n_61892), .C(n_332281799), .D(n_61871
		), .Z(n_332781804));
	notech_or4 i_12552950(.A(n_61892), .B(n_333081807), .C(n_61725), .D(n_61871
		), .Z(n_332981806));
	notech_and4 i_3953035(.A(n_1800), .B(n_1804), .C(n_1803), .D(n_1799), .Z
		(n_333081807));
	notech_and4 i_52438(.A(n_344281909), .B(n_341381880), .C(n_344381910), .D
		(n_332981806), .Z(n_333181808));
	notech_and3 i_18552890(.A(n_4351), .B(n_24142), .C(n_344881915), .Z(n_333381809
		));
	notech_and3 i_19052885(.A(n_2112), .B(n_416182412), .C(n_2111), .Z(n_333581810
		));
	notech_and4 i_19352882(.A(n_344981916), .B(n_4085), .C(n_333781812), .D(n_329681773
		), .Z(n_333681811));
	notech_or2 i_4053034(.A(n_2039), .B(n_411482388), .Z(n_333781812));
	notech_nand2 i_19152884(.A(n_344981916), .B(n_30868), .Z(n_333881813));
	notech_nao3 i_19252883(.A(n_329681773), .B(n_344981916), .C(n_32506), .Z
		(n_333981814));
	notech_or4 i_82452261(.A(n_340461032), .B(n_32217), .C(n_57256), .D(n_364628688
		), .Z(n_334081815));
	notech_nao3 i_82352262(.A(n_57395), .B(opd[24]), .C(n_57057), .Z(n_334981821
		));
	notech_nao3 i_82552260(.A(n_63774), .B(opc_10[24]), .C(n_299122016), .Z(n_335181822
		));
	notech_nand3 i_2521015(.A(n_346481931), .B(n_335181822), .C(n_334081815)
		, .Z(n_335281823));
	notech_or4 i_182851264(.A(n_340461032), .B(n_2830), .C(n_57251), .D(n_363350926
		), .Z(n_335381824));
	notech_or2 i_182751265(.A(n_25110), .B(nbus_11271[25]), .Z(n_335981827)
		);
	notech_or2 i_182251270(.A(n_365628696), .B(n_58438), .Z(n_336181828));
	notech_or2 i_182551267(.A(n_365228692), .B(n_33172), .Z(n_336481831));
	notech_nao3 i_182651266(.A(n_63790), .B(opc_10[25]), .C(n_365428694), .Z
		(n_336581832));
	notech_nand3 i_2621912(.A(n_336581832), .B(n_347281939), .C(n_335381824)
		, .Z(n_336681833));
	notech_or4 i_184751246(.A(n_340461032), .B(n_2830), .C(n_57251), .D(n_364628688
		), .Z(n_336781834));
	notech_or2 i_184651247(.A(n_25110), .B(nbus_11271[24]), .Z(n_337081837)
		);
	notech_or2 i_184151252(.A(n_365628696), .B(n_58429), .Z(n_337181838));
	notech_or2 i_184451249(.A(n_365228692), .B(n_33171), .Z(n_337481841));
	notech_nao3 i_184551248(.A(n_63790), .B(opc_10[24]), .C(n_365428694), .Z
		(n_337581842));
	notech_nand3 i_2521911(.A(n_348281948), .B(n_337581842), .C(n_336781834)
		, .Z(n_337681843));
	notech_or4 i_188451209(.A(n_340461032), .B(n_2830), .C(n_57251), .D(n_3464
		), .Z(n_337781844));
	notech_nand2 i_187651217(.A(tsc[54]), .B(n_30615), .Z(n_337881845));
	notech_or2 i_188351210(.A(n_25110), .B(n_60537), .Z(n_338081847));
	notech_or2 i_187851215(.A(n_365628696), .B(n_58411), .Z(n_338181848));
	notech_or2 i_188151212(.A(n_365228692), .B(n_33284), .Z(n_338481851));
	notech_nao3 i_188251211(.A(opc_10[22]), .B(n_63756), .C(n_365428694), .Z
		(n_338581852));
	notech_nand3 i_2321909(.A(n_349181957), .B(n_338581852), .C(n_337781844)
		, .Z(n_338681853));
	notech_or4 i_4153033(.A(n_49651676), .B(n_32397), .C(n_32383), .D(n_31407
		), .Z(n_338981856));
	notech_or4 i_216150933(.A(n_4106), .B(n_61871), .C(n_61675), .D(n_19680)
		, .Z(n_339081857));
	notech_or2 i_216050934(.A(vliw_pc[0]), .B(n_353728636), .Z(n_339181858)
		);
	notech_nand3 i_126958(.A(n_32186), .B(n_339181858), .C(n_339081857), .Z(n_339281859
		));
	notech_or4 i_6053014(.A(instrc[4]), .B(instrc[3]), .C(instrc[7]), .D(instrc
		[5]), .Z(n_339781864));
	notech_or4 i_6353011(.A(instrc[2]), .B(instrc[1]), .C(n_33321), .D(n_339781864
		), .Z(n_339881865));
	notech_or4 i_6153013(.A(fsmf[3]), .B(fsmf[0]), .C(fsmf[1]), .D(instrc[6]
		), .Z(n_340181868));
	notech_or4 i_6253012(.A(fsmf[4]), .B(fsmf[2]), .C(n_32548), .D(n_32091),
		 .Z(n_340481871));
	notech_or4 i_24577(.A(n_340481871), .B(n_340181868), .C(n_339881865), .D
		(n_30356), .Z(n_340781874));
	notech_nao3 i_79753069(.A(n_30383), .B(n_4338), .C(n_348471370), .Z(n_340981876
		));
	notech_and3 i_2553046(.A(n_330481781), .B(n_330381780), .C(n_330581782),
		 .Z(n_341381880));
	notech_ao4 i_8252992(.A(n_25676), .B(n_332760955), .C(n_383182262), .D(n_28008
		), .Z(n_341481881));
	notech_and2 i_8152993(.A(n_4090), .B(n_4089), .Z(n_341581882));
	notech_and3 i_9452981(.A(n_50148), .B(n_331581792), .C(n_331481791), .Z(n_342281889
		));
	notech_and3 i_9652979(.A(n_331681793), .B(n_342281889), .C(n_331781794),
		 .Z(n_342481891));
	notech_and4 i_10852967(.A(n_1808), .B(n_1805), .C(n_1809), .D(n_23326), 
		.Z(n_342881895));
	notech_and4 i_10652969(.A(n_1824), .B(n_1834), .C(n_4109), .D(n_23350), 
		.Z(n_342981896));
	notech_and4 i_10752968(.A(n_1807), .B(n_1844), .C(n_1820), .D(n_316860796
		), .Z(n_343181898));
	notech_nand3 i_2353047(.A(n_315760785), .B(n_32485), .C(n_316260790), .Z
		(n_343481901));
	notech_and4 i_12152954(.A(n_332581802), .B(n_364350916), .C(n_332681803)
		, .D(n_332781804), .Z(n_344281909));
	notech_ao4 i_12352952(.A(n_61846), .B(n_365128691), .C(n_1849), .D(n_28082
		), .Z(n_344381910));
	notech_and4 i_18952886(.A(n_1840), .B(n_4353), .C(n_4352), .D(n_4350), .Z
		(n_344881915));
	notech_ao4 i_653062(.A(n_61846), .B(n_333581810), .C(n_61859), .D(n_333381809
		), .Z(n_344981916));
	notech_or4 i_2753044(.A(n_19629), .B(n_59560), .C(n_19620), .D(n_349671381
		), .Z(n_345681923));
	notech_nand3 i_19552880(.A(n_62441), .B(n_333881813), .C(n_333981814), .Z
		(n_345881925));
	notech_ao4 i_82652259(.A(n_303922064), .B(nbus_11271[24]), .C(n_31532), 
		.D(n_61679), .Z(n_345981926));
	notech_ao4 i_82752258(.A(n_57362), .B(n_58893), .C(n_57363), .D(n_58429)
		, .Z(n_346181928));
	notech_ao4 i_82852257(.A(n_57319), .B(n_33171), .C(n_106826395), .D(n_57320
		), .Z(n_346281929));
	notech_and4 i_83152254(.A(n_346281929), .B(n_346181928), .C(n_345981926)
		, .D(n_334981821), .Z(n_346481931));
	notech_ao4 i_183351259(.A(n_101026337), .B(n_365328693), .C(n_365528695)
		, .D(n_58920), .Z(n_346681933));
	notech_ao4 i_182951263(.A(n_382264353), .B(n_31501), .C(n_56035), .D(n_32577
		), .Z(n_346781934));
	notech_and3 i_183151261(.A(n_350128600), .B(n_346781934), .C(n_335981827
		), .Z(n_346981936));
	notech_and4 i_183551257(.A(n_346681933), .B(n_336181828), .C(n_346981936
		), .D(n_336481831), .Z(n_347281939));
	notech_ao4 i_185351240(.A(n_365328693), .B(n_106826395), .C(n_365528695)
		, .D(n_58893), .Z(n_347481941));
	notech_ao4 i_184951244(.A(n_31500), .B(n_382264353), .C(n_56030), .D(n_32572
		), .Z(n_347681943));
	notech_and4 i_185151242(.A(n_55802), .B(n_347681943), .C(n_337081837), .D
		(n_437167955), .Z(n_347881945));
	notech_and4 i_185551238(.A(n_347881945), .B(n_347481941), .C(n_337181838
		), .D(n_337481841), .Z(n_348281948));
	notech_ao4 i_189051203(.A(n_59464), .B(n_365328693), .C(n_365528695), .D
		(n_58875), .Z(n_348481950));
	notech_ao4 i_188651207(.A(n_382264353), .B(n_31496), .C(n_31530), .D(n_61680
		), .Z(n_348681952));
	notech_and4 i_188851205(.A(n_55802), .B(n_348681952), .C(n_337881845), .D
		(n_338081847), .Z(n_348881954));
	notech_and4 i_189251201(.A(n_348881954), .B(n_348481950), .C(n_338181848
		), .D(n_338481851), .Z(n_349181957));
	notech_nand3 i_50349245(.A(n_61104), .B(n_61632), .C(read_data[3]), .Z(n_349581961
		));
	notech_or2 i_27649458(.A(n_55955), .B(n_30999), .Z(n_351881984));
	notech_nao3 i_27349461(.A(n_19612), .B(read_data[16]), .C(n_35412112), .Z
		(n_352181987));
	notech_or2 i_27049464(.A(n_126726594), .B(\nbus_11283[16] ), .Z(n_352481990
		));
	notech_or2 i_28949445(.A(n_55955), .B(n_31002), .Z(n_353181997));
	notech_nao3 i_28649448(.A(n_19612), .B(read_data[17]), .C(n_35412112), .Z
		(n_353482000));
	notech_or2 i_28349451(.A(n_126726594), .B(\nbus_11283[17] ), .Z(n_353782003
		));
	notech_or2 i_30249432(.A(n_55955), .B(n_31004), .Z(n_354482010));
	notech_nao3 i_29949435(.A(n_19612), .B(read_data[18]), .C(n_35412112), .Z
		(n_354782013));
	notech_or2 i_29649438(.A(n_126726594), .B(\nbus_11283[18] ), .Z(n_355082016
		));
	notech_or2 i_31549419(.A(n_55955), .B(n_31006), .Z(n_356282023));
	notech_nao3 i_31249422(.A(n_19612), .B(read_data[19]), .C(n_35412112), .Z
		(n_356882026));
	notech_or2 i_30949425(.A(n_126726594), .B(\nbus_11283[19] ), .Z(n_357182029
		));
	notech_nand3 i_50249246(.A(n_55904), .B(n_171160315), .C(n_1713), .Z(n_358182034
		));
	notech_ao3 i_79448958(.A(n_61680), .B(\opa_12[3] ), .C(n_2805), .Z(n_360082053
		));
	notech_ao4 i_196747826(.A(n_242970425), .B(n_31074), .C(n_242870424), .D
		(n_31072), .Z(n_365182102));
	notech_ao4 i_196647827(.A(n_243270428), .B(n_31075), .C(n_243170427), .D
		(n_31071), .Z(n_365282103));
	notech_ao4 i_196447829(.A(n_262170616), .B(n_31048), .C(n_57441), .D(n_31047
		), .Z(n_365582105));
	notech_ao4 i_196347830(.A(n_249970494), .B(n_31068), .C(n_249870493), .D
		(n_31067), .Z(n_365682106));
	notech_and4 i_196947824(.A(n_365682106), .B(n_365582105), .C(n_365282103
		), .D(n_365182102), .Z(n_365882108));
	notech_ao4 i_196047833(.A(n_321271180), .B(n_334760975), .C(n_30326), .D
		(n_30410), .Z(n_365982109));
	notech_ao4 i_195947834(.A(n_57034), .B(n_33476), .C(n_61104), .D(n_30866
		), .Z(n_366082110));
	notech_ao4 i_195747836(.A(n_58042), .B(n_31477), .C(n_56992), .D(n_31512
		), .Z(n_366282112));
	notech_ao4 i_195647837(.A(n_309771080), .B(n_33104), .C(n_309671079), .D
		(n_334660974), .Z(n_366382113));
	notech_and4 i_196247831(.A(n_366382113), .B(n_366282112), .C(n_366082110
		), .D(n_365982109), .Z(n_366582115));
	notech_ao4 i_193947854(.A(n_75522858), .B(n_242970425), .C(n_75622859), 
		.D(n_242870424), .Z(n_366682116));
	notech_ao4 i_193847855(.A(n_75222855), .B(n_243270428), .C(n_75322856), 
		.D(n_243170427), .Z(n_366782117));
	notech_ao4 i_193647857(.A(n_74822851), .B(n_262170616), .C(n_74922852), 
		.D(n_249870493), .Z(n_366982119));
	notech_ao4 i_193547858(.A(n_74522848), .B(n_249970494), .C(n_74622849), 
		.D(n_57441), .Z(n_367082120));
	notech_and4 i_194147852(.A(n_367082120), .B(n_366982119), .C(n_366782117
		), .D(n_366682116), .Z(n_367282122));
	notech_ao4 i_193247861(.A(n_30409), .B(n_30326), .C(n_338161009), .D(n_321271180
		), .Z(n_367382123));
	notech_ao4 i_193147862(.A(n_57034), .B(n_33477), .C(n_61104), .D(n_30863
		), .Z(n_367482124));
	notech_ao4 i_192947864(.A(n_58042), .B(n_31476), .C(n_56992), .D(n_31511
		), .Z(n_367682126));
	notech_ao4 i_192847865(.A(n_309771080), .B(n_33118), .C(n_338361011), .D
		(n_309671079), .Z(n_367782127));
	notech_and4 i_193447859(.A(n_367782127), .B(n_367682126), .C(n_367482124
		), .D(n_367382123), .Z(n_367982129));
	notech_ao4 i_192547868(.A(n_242970425), .B(n_326560893), .C(n_242870424)
		, .D(n_326760895), .Z(n_368082130));
	notech_ao4 i_192447869(.A(n_243270428), .B(n_326460892), .C(n_243170427)
		, .D(n_326660894), .Z(n_368182131));
	notech_ao4 i_192247871(.A(n_249870493), .B(n_326360891), .C(n_30326), .D
		(n_30408), .Z(n_368382133));
	notech_ao4 i_192147872(.A(n_325960887), .B(n_262170616), .C(n_249970494)
		, .D(n_326260890), .Z(n_368482134));
	notech_and4 i_192747866(.A(n_368482134), .B(n_368382133), .C(n_368182131
		), .D(n_368082130), .Z(n_368782136));
	notech_ao4 i_191847875(.A(n_321271180), .B(n_336160989), .C(n_326160889)
		, .D(n_57441), .Z(n_368882137));
	notech_ao4 i_191747876(.A(n_57034), .B(n_33478), .C(n_61104), .D(n_30862
		), .Z(n_368982138));
	notech_ao4 i_191547878(.A(n_58042), .B(n_31474), .C(n_56992), .D(n_31510
		), .Z(n_369182140));
	notech_ao4 i_191447879(.A(n_309771080), .B(n_33167), .C(n_309671079), .D
		(n_100842449), .Z(n_369282141));
	notech_and4 i_192047873(.A(n_369282141), .B(n_369182140), .C(n_368982138
		), .D(n_368882137), .Z(n_369482143));
	notech_nao3 i_47949736(.A(n_32310), .B(n_32323), .C(n_338161009), .Z(n_66222765
		));
	notech_ao4 i_187247921(.A(n_338361011), .B(n_30379), .C(n_61680), .D(n_31511
		), .Z(n_369582144));
	notech_ao4 i_187147922(.A(n_30378), .B(nbus_11273[3]), .C(n_30373), .D(\nbus_11290[3] 
		), .Z(n_369782146));
	notech_ao3 i_49149735(.A(n_369582144), .B(n_369782146), .C(n_360082053),
		 .Z(n_65022753));
	notech_ao4 i_162048173(.A(n_75222855), .B(n_28259), .C(n_28251), .D(n_74922852
		), .Z(n_369882147));
	notech_ao4 i_161948174(.A(n_75622859), .B(n_28258), .C(n_75322856), .D(n_28256
		), .Z(n_369982148));
	notech_ao4 i_161748176(.A(n_28260), .B(n_74822851), .C(n_75522858), .D(n_28255
		), .Z(n_370182150));
	notech_ao4 i_161648177(.A(n_74522848), .B(n_28252), .C(n_439367977), .D(n_74622849
		), .Z(n_370282151));
	notech_and4 i_162248171(.A(n_370282151), .B(n_370182150), .C(n_369982148
		), .D(n_369882147), .Z(n_370482153));
	notech_ao4 i_161348180(.A(n_61104), .B(n_30836), .C(n_338161009), .D(n_331660944
		), .Z(n_370582154));
	notech_ao4 i_161248181(.A(n_338361011), .B(n_439667980), .C(n_439467978)
		, .D(n_31476), .Z(n_370682155));
	notech_ao4 i_161048183(.A(n_55884), .B(n_33479), .C(n_439567979), .D(n_33118
		), .Z(n_370882157));
	notech_and4 i_161148182(.A(n_246070456), .B(n_370882157), .C(n_349581961
		), .D(n_358182034), .Z(n_371082159));
	notech_ao4 i_147248321(.A(n_337961007), .B(n_232870324), .C(n_337761005)
		, .D(nbus_11271[19]), .Z(n_371282161));
	notech_ao4 i_147148322(.A(n_127026597), .B(n_5356), .C(n_126226589), .D(n_319725273
		), .Z(n_371382162));
	notech_ao4 i_146948324(.A(n_126826595), .B(\nbus_11290[19] ), .C(n_126926596
		), .D(n_33202), .Z(n_371582164));
	notech_and4 i_147448319(.A(n_371582164), .B(n_371382162), .C(n_371282161
		), .D(n_357182029), .Z(n_371782166));
	notech_ao4 i_146648327(.A(n_61104), .B(n_30801), .C(n_337861006), .D(n_31492
		), .Z(n_371882167));
	notech_ao4 i_146448329(.A(n_55975), .B(n_32078), .C(n_55966), .D(n_33480
		), .Z(n_372082169));
	notech_and4 i_146848325(.A(n_372082169), .B(n_371882167), .C(n_356282023
		), .D(n_356882026), .Z(n_372282171));
	notech_ao4 i_146148332(.A(n_337961007), .B(n_235370349), .C(n_337761005)
		, .D(nbus_11271[18]), .Z(n_372382172));
	notech_ao4 i_146048333(.A(n_127026597), .B(n_5436), .C(n_126226589), .D(n_319825274
		), .Z(n_372482173));
	notech_ao4 i_145848335(.A(n_126826595), .B(\nbus_11290[18] ), .C(n_126926596
		), .D(n_33201), .Z(n_372682175));
	notech_and4 i_146348330(.A(n_372682175), .B(n_372482173), .C(n_372382172
		), .D(n_355082016), .Z(n_372882177));
	notech_ao4 i_145548338(.A(n_61104), .B(n_30799), .C(n_337861006), .D(n_31491
		), .Z(n_372982178));
	notech_ao4 i_145348340(.A(n_55975), .B(n_32077), .C(n_55966), .D(n_33481
		), .Z(n_373182180));
	notech_and4 i_145748336(.A(n_373182180), .B(n_372982178), .C(n_354482010
		), .D(n_354782013), .Z(n_373382182));
	notech_ao4 i_145048343(.A(n_337961007), .B(n_237870374), .C(n_337761005)
		, .D(nbus_11271[17]), .Z(n_373482183));
	notech_ao4 i_144948344(.A(n_5397), .B(n_127026597), .C(n_126226589), .D(n_319951172
		), .Z(n_373582184));
	notech_ao4 i_144748346(.A(n_126826595), .B(\nbus_11290[17] ), .C(n_126926596
		), .D(n_33200), .Z(n_373782186));
	notech_and4 i_145248341(.A(n_373782186), .B(n_373582184), .C(n_373482183
		), .D(n_353782003), .Z(n_373982188));
	notech_ao4 i_144448349(.A(n_61087), .B(n_30797), .C(n_337861006), .D(n_31490
		), .Z(n_374082189));
	notech_ao4 i_144248351(.A(n_55975), .B(n_32076), .C(n_55966), .D(n_33482
		), .Z(n_374282191));
	notech_and4 i_144648347(.A(n_374282191), .B(n_374082189), .C(n_353181997
		), .D(n_353482000), .Z(n_374482193));
	notech_ao4 i_143948354(.A(n_337961007), .B(n_240370399), .C(n_337761005)
		, .D(nbus_11271[16]), .Z(n_374582194));
	notech_ao4 i_143848355(.A(n_127026597), .B(n_5444), .C(n_126226589), .D(n_320051171
		), .Z(n_374682195));
	notech_ao4 i_143648357(.A(n_126826595), .B(\nbus_11290[16] ), .C(n_126926596
		), .D(n_33199), .Z(n_374882197));
	notech_and4 i_144148352(.A(n_374882197), .B(n_374682195), .C(n_374582194
		), .D(n_352481990), .Z(n_375082199));
	notech_ao4 i_143348360(.A(n_61087), .B(n_30795), .C(n_337861006), .D(n_31489
		), .Z(n_375182200));
	notech_ao4 i_143148362(.A(n_55975), .B(n_32075), .C(n_55966), .D(n_33483
		), .Z(n_375382202));
	notech_and4 i_143548358(.A(n_375382202), .B(n_375182200), .C(n_351881984
		), .D(n_352181987), .Z(n_375582204));
	notech_ao4 i_122348558(.A(n_74922852), .B(n_23510), .C(n_58702), .D(n_66222765
		), .Z(n_375682205));
	notech_ao4 i_122248559(.A(n_75322856), .B(n_23514), .C(n_75222855), .D(n_23517
		), .Z(n_375782206));
	notech_ao4 i_122048561(.A(n_75522858), .B(n_23518), .C(n_75622859), .D(n_23515
		), .Z(n_375982208));
	notech_ao4 i_121948562(.A(n_74622849), .B(n_334560973), .C(n_74822851), 
		.D(n_23519), .Z(n_3760));
	notech_and4 i_122548556(.A(n_3760), .B(n_375982208), .C(n_375782206), .D
		(n_375682205), .Z(n_376282210));
	notech_ao4 i_121648565(.A(n_334460972), .B(n_31476), .C(n_74522848), .D(n_23511
		), .Z(n_3763));
	notech_ao4 i_121548566(.A(n_391264443), .B(n_33118), .C(n_338361011), .D
		(n_391164442), .Z(n_376482211));
	notech_ao4 i_121348568(.A(n_56030), .B(n_32531), .C(n_58664), .D(nbus_11271
		[3]), .Z(n_376682213));
	notech_and4 i_121848563(.A(n_65022753), .B(n_376682213), .C(n_376482211)
		, .D(n_3763), .Z(n_376882214));
	notech_nao3 i_82963398(.A(n_57494), .B(n_30658), .C(n_29758), .Z(n_376982215
		));
	notech_nao3 i_91563392(.A(n_32259), .B(n_30658), .C(n_29758), .Z(n_3770)
		);
	notech_nand2 i_103145425(.A(n_32224), .B(n_115442595), .Z(n_377382218)
		);
	notech_nao3 i_103245424(.A(n_57494), .B(n_30658), .C(n_379164322), .Z(n_377482219
		));
	notech_or2 i_43445985(.A(n_55955), .B(n_31030), .Z(n_377782222));
	notech_or2 i_43145988(.A(n_337761005), .B(nbus_11271[31]), .Z(n_378082225
		));
	notech_or2 i_42845991(.A(n_5243), .B(n_127026597), .Z(n_3783));
	notech_nao3 i_76145678(.A(n_19655), .B(read_data[9]), .C(n_60453), .Z(n_379082232
		));
	notech_nand2 i_75445685(.A(n_300322028), .B(opd[9]), .Z(n_379782238));
	notech_ao4 i_180744706(.A(n_327160899), .B(n_265070645), .C(n_327360901)
		, .D(n_264970644), .Z(n_3802));
	notech_ao4 i_180644707(.A(n_299222017), .B(n_59032), .C(n_327260900), .D
		(n_265370646), .Z(n_380382242));
	notech_ao4 i_180444709(.A(n_327060898), .B(n_299422019), .C(n_265570648)
		, .D(n_58294), .Z(n_3805));
	notech_and4 i_180944704(.A(n_3805), .B(n_380382242), .C(n_3802), .D(n_379782238
		), .Z(n_3807));
	notech_ao4 i_180144712(.A(n_309871081), .B(n_336660994), .C(n_30326), .D
		(n_30412), .Z(n_3808));
	notech_ao4 i_180044713(.A(n_310771089), .B(n_99942440), .C(n_61087), .D(n_30874
		), .Z(n_380982245));
	notech_ao4 i_179844715(.A(n_57034), .B(n_33484), .C(n_310371085), .D(n_33168
		), .Z(n_381182247));
	notech_and4 i_180344710(.A(n_381182247), .B(n_380982245), .C(n_3808), .D
		(n_379082232), .Z(n_3813));
	notech_ao4 i_148645020(.A(n_300822033), .B(n_126226589), .C(n_337961007)
		, .D(n_262470619), .Z(n_3814));
	notech_ao4 i_148545021(.A(n_337861006), .B(n_31507), .C(n_61087), .D(n_30809
		), .Z(n_3815));
	notech_ao4 i_148345023(.A(n_126926596), .B(n_33206), .C(n_55946), .D(n_31539
		), .Z(n_3817));
	notech_and4 i_148845018(.A(n_3817), .B(n_3815), .C(n_3814), .D(n_3783), 
		.Z(n_381982250));
	notech_ao4 i_148045026(.A(n_126726594), .B(\nbus_11283[31] ), .C(n_126826595
		), .D(\nbus_11290[31] ), .Z(n_382082251));
	notech_ao4 i_147845028(.A(n_55975), .B(n_32090), .C(n_55966), .D(n_33485
		), .Z(n_382282253));
	notech_and4 i_148245024(.A(n_382282253), .B(n_378082225), .C(n_382082251
		), .D(n_377782222), .Z(n_382482255));
	notech_ao4 i_161443316(.A(n_32590), .B(n_61630), .C(n_30364), .D(n_30361
		), .Z(n_382582256));
	notech_or4 i_101943285(.A(n_61912), .B(n_61901), .C(n_61892), .D(n_32397
		), .Z(n_25705));
	notech_nand3 i_20743083(.A(n_57472), .B(n_30363), .C(n_57461), .Z(n_382682257
		));
	notech_or4 i_22943061(.A(mask8b[1]), .B(mask8b[0]), .C(n_30370), .D(n_31069
		), .Z(n_382882259));
	notech_or4 i_35342937(.A(n_61725), .B(n_61892), .C(n_4440), .D(\nbus_11290[7] 
		), .Z(n_382982260));
	notech_and2 i_159943351(.A(n_26637), .B(n_339661024), .Z(n_383182262));
	notech_or4 i_56942722(.A(n_301960648), .B(n_61725), .C(n_61680), .D(n_19734
		), .Z(n_383382264));
	notech_nand2 i_57042721(.A(n_31069), .B(n_414582401), .Z(n_383482265));
	notech_or4 i_57242719(.A(instrc[121]), .B(n_2577), .C(instrc[122]), .D(n_32265
		), .Z(n_383582266));
	notech_and2 i_58242711(.A(n_4036), .B(n_1823), .Z(n_384082271));
	notech_and2 i_106942271(.A(instrc[106]), .B(n_32227), .Z(n_384382274));
	notech_and3 i_107142269(.A(n_19672), .B(n_61630), .C(n_30374), .Z(n_384582276
		));
	notech_or4 i_14443145(.A(n_340561033), .B(n_32627), .C(n_61630), .D(nbus_11271
		[11]), .Z(n_384682277));
	notech_nand2 i_14343146(.A(resb_shiftbox[3]), .B(n_30417), .Z(n_384982280
		));
	notech_or4 i_14043149(.A(n_4025), .B(n_60177), .C(n_61630), .D(n_31476),
		 .Z(n_385282283));
	notech_or2 i_13743152(.A(n_61016485), .B(nbus_11271[3]), .Z(n_385582286)
		);
	notech_or2 i_13243157(.A(n_61516490), .B(n_58974), .Z(n_386082290));
	notech_nand2 i_12943160(.A(read_data[27]), .B(n_26116136), .Z(n_386382293
		));
	notech_nand2 i_12643163(.A(n_30416), .B(add_src[3]), .Z(n_3866));
	notech_or4 i_23243058(.A(n_28534), .B(n_60189), .C(n_32576), .D(n_61630)
		, .Z(n_386982298));
	notech_or4 i_33542955(.A(n_28098), .B(n_340561033), .C(n_61630), .D(nbus_11271
		[5]), .Z(n_387082299));
	notech_or2 i_33042960(.A(n_60316478), .B(n_31486), .Z(n_387782304));
	notech_nand2 i_32142969(.A(add_src[13]), .B(n_30416), .Z(n_3886));
	notech_or2 i_54042750(.A(n_60516480), .B(n_58474), .Z(n_3891));
	notech_or4 i_53742753(.A(n_61892), .B(n_3964), .C(n_61725), .D(n_33161),
		 .Z(n_3894));
	notech_or4 i_31466(.A(n_32396), .B(n_28534), .C(n_63700), .D(n_63756), .Z
		(n_27932));
	notech_and2 i_20625(.A(n_61680), .B(opb[7]), .Z(n_21074));
	notech_and2 i_106842272(.A(imm[7]), .B(n_32216), .Z(n_3931));
	notech_ao4 i_176041594(.A(n_57472), .B(n_31703), .C(n_57456), .D(n_31671
		), .Z(n_3934));
	notech_ao4 i_175941595(.A(n_57627), .B(n_33486), .C(n_30363), .D(n_31735
		), .Z(n_3935));
	notech_ao4 i_175741597(.A(n_57506), .B(n_31799), .C(n_57494), .D(n_31767
		), .Z(n_393782333));
	notech_ao4 i_175641598(.A(n_57517), .B(n_31863), .C(n_58550), .D(n_31831
		), .Z(n_3938));
	notech_and4 i_176241592(.A(n_3938), .B(n_393782333), .C(n_3935), .D(n_3934
		), .Z(n_3940));
	notech_ao4 i_175341601(.A(n_57417), .B(n_31927), .C(n_57407), .D(n_31895
		), .Z(n_3941));
	notech_ao4 i_175241602(.A(n_57449), .B(n_31600), .C(n_57435), .D(n_31960
		), .Z(n_3942));
	notech_and2 i_175441600(.A(n_3942), .B(n_3941), .Z(n_3943));
	notech_ao4 i_175041604(.A(n_30664), .B(n_31436), .C(n_57524), .D(n_33487
		), .Z(n_3944));
	notech_ao4 i_174941605(.A(n_58597), .B(n_32024), .C(n_58566), .D(n_31992
		), .Z(n_394582334));
	notech_ao4 i_174641608(.A(n_57467), .B(n_31704), .C(n_57456), .D(n_31672
		), .Z(n_3948));
	notech_ao4 i_174541609(.A(n_57627), .B(n_33488), .C(n_30363), .D(n_31736
		), .Z(n_394982337));
	notech_ao4 i_174341611(.A(n_57506), .B(n_31800), .C(n_57489), .D(n_31768
		), .Z(n_3951));
	notech_ao4 i_174241612(.A(n_57517), .B(n_31864), .C(n_58550), .D(n_31832
		), .Z(n_3952));
	notech_and4 i_174841606(.A(n_3952), .B(n_3951), .C(n_394982337), .D(n_3948
		), .Z(n_3954));
	notech_ao4 i_173941615(.A(n_57412), .B(n_31928), .C(n_57407), .D(n_31896
		), .Z(n_3955));
	notech_ao4 i_173841616(.A(n_57444), .B(n_31601), .C(n_57435), .D(n_31961
		), .Z(n_3956));
	notech_and2 i_174041614(.A(n_3956), .B(n_3955), .Z(n_3957));
	notech_ao4 i_173641618(.A(n_30664), .B(n_31437), .C(n_57524), .D(n_33489
		), .Z(n_395882339));
	notech_ao4 i_173541619(.A(n_58597), .B(n_32025), .C(n_58566), .D(n_31993
		), .Z(n_3959));
	notech_and3 i_199743269(.A(n_19672), .B(n_61630), .C(n_32487), .Z(n_396382340
		));
	notech_or2 i_63143315(.A(n_382582256), .B(n_33157), .Z(n_61816493));
	notech_or4 i_171641638(.A(n_32574), .B(n_25681), .C(n_63758), .D(n_61958
		), .Z(n_3964));
	notech_or4 i_64443311(.A(n_61912), .B(n_61901), .C(n_61892), .D(n_3964),
		 .Z(n_61116486));
	notech_or4 i_67143308(.A(n_61912), .B(n_61901), .C(n_61892), .D(n_384082271
		), .Z(n_61016485));
	notech_nand3 i_64743310(.A(n_27823), .B(n_30364), .C(n_396382340), .Z(n_60916484
		));
	notech_or4 i_62843317(.A(n_60189), .B(n_32574), .C(n_25681), .D(n_61632)
		, .Z(n_60516480));
	notech_or4 i_64343312(.A(n_61892), .B(n_4025), .C(n_60177), .D(n_61725),
		 .Z(n_60316478));
	notech_or2 i_63843313(.A(n_382582256), .B(instrc[107]), .Z(n_60216477)
		);
	notech_ao4 i_643324(.A(n_33164), .B(n_57622), .C(instrc[121]), .D(n_32305
		), .Z(n_396682342));
	notech_or4 i_60543318(.A(n_32396), .B(n_28534), .C(n_60157), .D(n_61632)
		, .Z(n_59316468));
	notech_ao4 i_139643284(.A(n_4432), .B(n_58116456), .C(n_61816493), .D(n_4441
		), .Z(n_58016455));
	notech_ao4 i_168741666(.A(n_61716492), .B(n_32264), .C(n_4438), .D(n_31537
		), .Z(n_396782343));
	notech_ao4 i_168641667(.A(n_323151206), .B(n_58947), .C(n_4436), .D(n_32343
		), .Z(n_396882344));
	notech_ao4 i_168441669(.A(n_60916484), .B(n_32238), .C(n_61016485), .D(n_60620
		), .Z(n_3970));
	notech_and4 i_168941664(.A(n_3894), .B(n_3970), .C(n_396882344), .D(n_396782343
		), .Z(n_397282345));
	notech_ao4 i_168141672(.A(n_4428), .B(n_60216477), .C(n_60316478), .D(n_31505
		), .Z(n_3973));
	notech_ao4 i_167941674(.A(n_4437), .B(n_32189), .C(n_59316468), .D(n_32732
		), .Z(n_3975));
	notech_and4 i_168341670(.A(n_325885670), .B(n_3975), .C(n_3973), .D(n_3891
		), .Z(n_3977));
	notech_or4 i_71343301(.A(n_32576), .B(n_60177), .C(n_28534), .D(n_61632)
		, .Z(n_40616281));
	notech_or2 i_70043306(.A(n_59316468), .B(n_27843), .Z(n_40316278));
	notech_or4 i_70943304(.A(n_25681), .B(n_25705), .C(n_32646), .D(n_63800)
		, .Z(n_40216277));
	notech_or2 i_70143305(.A(n_59316468), .B(n_30521), .Z(n_40116276));
	notech_ao4 i_183743274(.A(n_58541), .B(n_61632), .C(n_27909), .D(n_383182262
		), .Z(n_397882347));
	notech_ao4 i_148441861(.A(n_61716492), .B(n_32262), .C(n_4438), .D(n_31521
		), .Z(n_3979));
	notech_ao4 i_148341862(.A(n_40616281), .B(n_32257), .C(n_443982453), .D(\nbus_11290[13] 
		), .Z(n_398182349));
	notech_and3 i_148641859(.A(n_3979), .B(n_398182349), .C(n_3886), .Z(n_398282350
		));
	notech_ao4 i_148141864(.A(n_40116276), .B(n_32878), .C(n_40216277), .D(n_31505
		), .Z(n_398382351));
	notech_ao4 i_148041865(.A(n_61016485), .B(nbus_11271[13]), .C(n_40316278
		), .D(n_32716), .Z(n_398482352));
	notech_ao4 i_147641869(.A(n_61116486), .B(n_33147), .C(n_60916484), .D(n_32213
		), .Z(n_398782355));
	notech_ao4 i_147541870(.A(n_60516480), .B(nbus_11273[13]), .C(n_60216477
		), .D(n_375064281), .Z(n_398982357));
	notech_ao4 i_147341872(.A(n_56929), .B(n_58947), .C(n_4437), .D(n_32170)
		, .Z(n_3991));
	notech_and4 i_147441871(.A(n_58016455), .B(n_3991), .C(n_382982260), .D(n_387082299
		), .Z(n_3993));
	notech_and4 i_147941866(.A(n_387782304), .B(n_398782355), .C(n_398982357
		), .D(n_3993), .Z(n_3994));
	notech_or4 i_75143296(.A(n_30370), .B(mask8b[0]), .C(n_31069), .D(n_31066
		), .Z(n_26716142));
	notech_and4 i_75043297(.A(mask8b[0]), .B(n_414582401), .C(mask8b[2]), .D
		(n_31066), .Z(n_26316138));
	notech_and4 i_74743298(.A(mask8b[0]), .B(mask8b[1]), .C(mask8b[2]), .D(n_414582401
		), .Z(n_26116136));
	notech_ao4 i_138241959(.A(n_25468), .B(n_61632), .C(n_25705), .D(n_4025)
		, .Z(n_4000));
	notech_nao3 i_98843287(.A(n_382682257), .B(instrc[107]), .C(n_382582256)
		, .Z(n_23916114));
	notech_ao4 i_98343289(.A(n_58116456), .B(n_4432), .C(n_396682342), .D(n_61816493
		), .Z(n_22216097));
	notech_nao3 i_130242039(.A(instrc[121]), .B(n_59558), .C(n_32305), .Z(n_400482361
		));
	notech_ao4 i_129842043(.A(n_23916114), .B(n_32260), .C(n_61816493), .D(n_400482361
		), .Z(n_400582362));
	notech_ao4 i_129642045(.A(n_30605), .B(n_31519), .C(n_26716142), .D(n_31527
		), .Z(n_400782364));
	notech_and4 i_130042041(.A(n_400782364), .B(n_400582362), .C(n_3866), .D
		(n_386382293), .Z(n_400982366));
	notech_ao4 i_129342048(.A(n_40616281), .B(n_32258), .C(n_4434), .D(n_31511
		), .Z(n_401082367));
	notech_ao4 i_129242049(.A(n_40116276), .B(n_32868), .C(n_40216277), .D(n_31492
		), .Z(n_401282369));
	notech_and4 i_130142040(.A(n_401082367), .B(n_401282369), .C(n_400982366
		), .D(n_386082290), .Z(n_4014));
	notech_ao4 i_128842053(.A(n_4433), .B(\nbus_11290[3] ), .C(n_40316278), 
		.D(n_32706), .Z(n_4015));
	notech_ao4 i_128642055(.A(n_61116486), .B(n_32150), .C(n_60916484), .D(n_32201
		), .Z(n_4017));
	notech_and4 i_129042051(.A(n_4017), .B(n_4015), .C(n_385282283), .D(n_385582286
		), .Z(n_4019));
	notech_ao4 i_128342058(.A(n_60516480), .B(nbus_11273[3]), .C(n_60216477)
		, .D(n_338361011), .Z(n_4020));
	notech_and4 i_128542056(.A(n_22216097), .B(n_4020), .C(n_384982280), .D(n_384682277
		), .Z(n_4023));
	notech_or4 i_54540114(.A(n_32184), .B(n_314960777), .C(n_32646), .D(n_61823
		), .Z(n_4025));
	notech_or4 i_63940112(.A(n_32576), .B(n_28098), .C(n_60159), .D(n_61632)
		, .Z(n_25433));
	notech_or2 i_57940091(.A(n_4086), .B(n_19548), .Z(n_24134));
	notech_nand3 i_63340089(.A(sign_div), .B(n_30371), .C(opd[31]), .Z(n_24138
		));
	notech_nand2 i_63540088(.A(n_30371), .B(n_24147), .Z(n_24144));
	notech_or4 i_64540087(.A(n_32576), .B(n_32397), .C(n_28534), .D(n_61632)
		, .Z(n_24141));
	notech_and3 i_64940085(.A(n_405882374), .B(n_4057), .C(n_57878), .Z(n_24127
		));
	notech_nao3 i_70540082(.A(n_28092), .B(n_316260790), .C(n_61892), .Z(n_23989
		));
	notech_and4 i_5340023(.A(n_4453), .B(n_444982454), .C(n_4028), .D(n_30365
		), .Z(n_4026));
	notech_nao3 i_109139016(.A(n_317051260), .B(n_406282377), .C(n_56930), .Z
		(n_4028));
	notech_mux2 i_8439992(.S(n_32321), .A(\nbus_11283[31] ), .B(n_58348), .Z
		(n_4030));
	notech_or2 i_110439003(.A(n_27843), .B(\nbus_11283[31] ), .Z(n_4033));
	notech_or4 i_110639001(.A(n_61917), .B(n_61903), .C(n_61892), .D(n_4036)
		, .Z(n_4035));
	notech_ao4 i_55440132(.A(n_26637), .B(n_32627), .C(n_60189), .D(n_4025),
		 .Z(n_4036));
	notech_nand2 i_110938998(.A(n_56572), .B(n_56661), .Z(n_4039));
	notech_or4 i_94839158(.A(n_30636), .B(n_30343), .C(n_61680), .D(n_31528)
		, .Z(n_4040));
	notech_ao4 i_94939157(.A(n_4442), .B(n_23845), .C(opc[3]), .D(opc[2]), .Z
		(n_4056));
	notech_nand2 i_35562(.A(rep_en1), .B(n_406282377), .Z(n_23836));
	notech_or4 i_35559(.A(n_4086), .B(n_57336), .C(n_19548), .D(n_27823), .Z
		(n_23839));
	notech_or4 i_109339014(.A(n_340561033), .B(n_28008), .C(n_61632), .D(n_4030
		), .Z(n_4057));
	notech_or4 i_109439013(.A(n_26637), .B(n_28098), .C(nbus_11271[15]), .D(n_61632
		), .Z(n_405882374));
	notech_nor2 i_33953(.A(n_59120), .B(n_61632), .Z(n_405982375));
	notech_or4 i_31489(.A(n_61917), .B(n_61903), .C(n_61892), .D(n_28008), .Z
		(n_27909));
	notech_ao3 i_178340065(.A(n_30364), .B(n_30691), .C(n_4086), .Z(n_406282377
		));
	notech_ao4 i_212338026(.A(n_57679), .B(nbus_11273[7]), .C(n_336360991), 
		.D(n_58348), .Z(n_406382378));
	notech_nand2 i_190838232(.A(nbus_11271[4]), .B(opc[3]), .Z(n_406882382)
		);
	notech_or4 i_190738233(.A(n_23847), .B(nbus_11271[0]), .C(nbus_11271[1])
		, .D(nbus_11271[2]), .Z(n_406982383));
	notech_ao4 i_190338237(.A(n_4026), .B(nbus_11271[4]), .C(n_406882382), .D
		(n_406982383), .Z(n_4071));
	notech_ao4 i_190238238(.A(n_24141), .B(nbus_11271[28]), .C(n_23989), .D(n_33392
		), .Z(n_4072));
	notech_ao4 i_190038240(.A(n_24138), .B(n_33490), .C(n_24144), .D(nbus_11270
		[4]), .Z(n_407482384));
	notech_ao4 i_189938241(.A(n_23836), .B(n_33491), .C(n_218373551), .D(n_33493
		), .Z(n_4075));
	notech_and4 i_190538235(.A(n_4075), .B(n_407482384), .C(n_4072), .D(n_4071
		), .Z(n_407782385));
	notech_ao4 i_189638244(.A(n_25433), .B(n_59050), .C(n_23839), .D(n_33492
		), .Z(n_4078));
	notech_ao4 i_189538245(.A(n_4446), .B(\nbus_11290[4] ), .C(n_4447), .D(n_31615
		), .Z(n_4079));
	notech_ao4 i_189338247(.A(n_30712), .B(n_32918), .C(n_4444), .D(n_1839),
		 .Z(n_4081));
	notech_and3 i_189438246(.A(n_24127), .B(n_4081), .C(n_4040), .Z(n_4083)
		);
	notech_or4 i_207637602(.A(n_61917), .B(n_61903), .C(n_317460802), .D(n_33242
		), .Z(n_4085));
	notech_nand3 i_56937535(.A(n_30636), .B(n_32481), .C(n_61632), .Z(n_4086
		));
	notech_and3 i_78737516(.A(n_32353), .B(n_32481), .C(n_30450), .Z(n_29906
		));
	notech_ao4 i_166237476(.A(n_24142), .B(n_61859), .C(n_4458), .D(n_61846)
		, .Z(n_4088));
	notech_and3 i_177237472(.A(n_4036), .B(n_32590), .C(n_415882410), .Z(n_4089
		));
	notech_and4 i_183837469(.A(n_1824), .B(n_1834), .C(n_4109), .D(n_4108), 
		.Z(n_4090));
	notech_or4 i_202737447(.A(instrc[94]), .B(n_32484), .C(instrc[92]), .D(n_61684
		), .Z(n_28572));
	notech_or4 i_202937446(.A(instrc[90]), .B(n_32484), .C(instrc[88]), .D(n_61680
		), .Z(n_28581));
	notech_nand3 i_11637382(.A(n_4146), .B(n_4088), .C(n_4468), .Z(n_4091)
		);
	notech_ao4 i_15937341(.A(n_30628), .B(n_331271269), .C(n_311371095), .D(n_30307
		), .Z(n_409282386));
	notech_nao3 i_16037340(.A(n_414482400), .B(n_4097), .C(n_4143), .Z(n_4093
		));
	notech_and4 i_16137339(.A(n_56794), .B(n_22474), .C(n_22467), .D(n_348071366
		), .Z(n_4094));
	notech_and4 i_16237338(.A(n_4319), .B(n_4460), .C(n_22481), .D(n_4461), 
		.Z(n_4095));
	notech_or2 i_27737265(.A(n_57105), .B(n_33242), .Z(n_4097));
	notech_nand2 i_28737256(.A(n_4099), .B(n_33495), .Z(n_4098));
	notech_nand2 i_19513(.A(n_33495), .B(n_4329), .Z(n_4099));
	notech_and4 i_11737381(.A(n_56930), .B(n_30691), .C(n_415282404), .D(n_56572
		), .Z(n_4102));
	notech_nand2 i_11837380(.A(n_57336), .B(n_30937), .Z(n_4105));
	notech_or2 i_553063(.A(n_340781874), .B(n_30364), .Z(n_4106));
	notech_and3 i_43337127(.A(n_316471137), .B(n_30560), .C(n_3469), .Z(n_4107
		));
	notech_or4 i_47237089(.A(n_32576), .B(n_28098), .C(n_63720), .D(n_63782)
		, .Z(n_4108));
	notech_or4 i_47337088(.A(calc_sz[3]), .B(calc_sz[2]), .C(n_317960807), .D
		(n_58541), .Z(n_4109));
	notech_ao4 i_11037388(.A(n_4292), .B(n_30374), .C(n_2039), .D(n_411482388
		), .Z(n_4110));
	notech_or4 i_50237061(.A(n_61859), .B(n_61632), .C(n_33496), .D(n_4112),
		 .Z(n_4111));
	notech_and3 i_11137387(.A(n_4288), .B(n_4287), .C(n_4291), .Z(n_4112));
	notech_or4 i_3253042(.A(n_26133), .B(n_4106), .C(n_345681923), .D(n_349971384
		), .Z(n_411482388));
	notech_ao3 i_9937399(.A(n_323060858), .B(n_4179), .C(n_322960857), .Z(n_411582389
		));
	notech_and4 i_10037398(.A(n_116645658), .B(n_30798), .C(n_339261020), .D
		(n_4178), .Z(n_411682390));
	notech_ao4 i_10137397(.A(n_59312350), .B(n_4276), .C(n_58566), .D(n_365964190
		), .Z(n_411782391));
	notech_nand3 i_58936994(.A(n_376464295), .B(n_412082394), .C(n_417782425
		), .Z(n_411982393));
	notech_or4 i_11537383(.A(n_32575), .B(n_32383), .C(n_63700), .D(n_61940)
		, .Z(n_412082394));
	notech_nand2 i_59036993(.A(n_391464445), .B(n_391364444), .Z(n_412182395
		));
	notech_and3 i_9437404(.A(n_71912476), .B(n_4193), .C(n_4192), .Z(n_412282396
		));
	notech_ao3 i_9337405(.A(n_4262), .B(n_4459), .C(n_30375), .Z(n_412382397
		));
	notech_and3 i_9637402(.A(n_4364), .B(n_418882429), .C(n_4257), .Z(n_412482398
		));
	notech_and4 i_9837400(.A(n_30679), .B(n_418882429), .C(n_4364), .D(n_4257
		), .Z(n_412582399));
	notech_ao4 i_8537413(.A(n_32697), .B(n_30965), .C(n_247980969), .D(n_32323
		), .Z(n_4126));
	notech_or4 i_63736952(.A(n_72112478), .B(n_4086), .C(n_19637), .D(n_4251
		), .Z(n_4128));
	notech_nor2 i_3637431(.A(n_4236), .B(n_4219), .Z(n_4129));
	notech_ao4 i_9537403(.A(n_4200), .B(n_30336), .C(n_33242), .D(n_4238), .Z
		(n_4130));
	notech_nao3 i_27237269(.A(n_32506), .B(n_30650), .C(n_4085), .Z(n_4134)
		);
	notech_and4 i_26737274(.A(n_61632), .B(n_61087), .C(n_4093), .D(n_4338),
		 .Z(n_4141));
	notech_or4 i_27837264(.A(n_30304), .B(n_61892), .C(n_316260790), .D(read_ack
		), .Z(n_4142));
	notech_ao3 i_27437267(.A(n_30382), .B(n_30381), .C(n_347671363), .Z(n_4143
		));
	notech_nand2 i_27637266(.A(n_33242), .B(n_30680), .Z(n_414482400));
	notech_or4 i_35410(.A(n_317460802), .B(n_61723), .C(n_30343), .D(n_61680
		), .Z(n_23988));
	notech_and2 i_33709(.A(n_19734), .B(n_61628), .Z(n_414582401));
	notech_and2 i_19105(.A(n_4091), .B(n_62441), .Z(\nbus_11289[0] ));
	notech_or2 i_42337136(.A(n_4102), .B(n_4465), .Z(n_4146));
	notech_nao3 i_42737132(.A(n_30691), .B(n_4105), .C(n_4465), .Z(n_4148)
		);
	notech_nand3 i_42937131(.A(n_579), .B(n_19698), .C(n_30869), .Z(n_414982402
		));
	notech_or4 i_43037130(.A(n_348471370), .B(n_4106), .C(n_59560), .D(n_2091
		), .Z(n_4150));
	notech_nand2 i_42437135(.A(rep_en5), .B(n_30372), .Z(n_415282404));
	notech_nao3 i_31485(.A(n_2113), .B(n_30364), .C(n_313471111), .Z(n_415382405
		));
	notech_nao3 i_46837093(.A(pipe_mul[1]), .B(n_28092), .C(pipe_mul[0]), .Z
		(n_415482406));
	notech_or4 i_47137090(.A(n_32576), .B(n_59120), .C(n_61940), .D(n_61958)
		, .Z(n_415782409));
	notech_or4 i_47437087(.A(n_32576), .B(n_32627), .C(n_63700), .D(n_63782)
		, .Z(n_415882410));
	notech_nao3 i_49837063(.A(n_62441), .B(n_30377), .C(n_4110), .Z(n_415982411
		));
	notech_or4 i_50137062(.A(n_348889370), .B(n_19680), .C(n_19672), .D(n_59100
		), .Z(n_4160));
	notech_and2 i_37176(.A(n_4337), .B(n_329381770), .Z(n_416182412));
	notech_or4 i_58037002(.A(instrc[98]), .B(instrc[97]), .C(n_26978), .D(n_30550
		), .Z(n_416982420));
	notech_or4 i_57737005(.A(instrc[113]), .B(instrc[114]), .C(n_2830), .D(n_114845640
		), .Z(n_4172));
	notech_nao3 i_57237010(.A(n_29906), .B(n_33142), .C(n_375264283), .Z(n_417382423
		));
	notech_or4 i_57337009(.A(n_30551), .B(n_371764248), .C(n_29232), .D(instrc
		[107]), .Z(n_4174));
	notech_or4 i_57437008(.A(instrc[122]), .B(n_32275), .C(n_111445606), .D(instrc
		[120]), .Z(n_417582424));
	notech_nand2 i_11437384(.A(n_31160), .B(n_412182395), .Z(n_417782425));
	notech_nand2 i_58436998(.A(n_321860846), .B(n_58702), .Z(n_4178));
	notech_nand3 i_58336999(.A(n_321860846), .B(n_58701), .C(n_63758), .Z(n_4179
		));
	notech_or4 i_63336956(.A(n_61940), .B(n_56003), .C(n_32323), .D(n_30904)
		, .Z(n_418882429));
	notech_nand3 i_63136958(.A(n_57638), .B(n_63758), .C(n_30788), .Z(n_418982430
		));
	notech_nand3 i_63236957(.A(n_30903), .B(n_32273), .C(n_32323), .Z(n_419082431
		));
	notech_and4 i_62336963(.A(n_4126), .B(n_33162), .C(\opcode[0] ), .D(n_30842
		), .Z(n_419182432));
	notech_or4 i_63836951(.A(n_301560644), .B(n_301760646), .C(n_30331), .D(n_4129
		), .Z(n_4192));
	notech_nao3 i_63936950(.A(n_19603), .B(n_19612), .C(n_4130), .Z(n_4193)
		);
	notech_or4 i_64236947(.A(n_4466), .B(n_30839), .C(instrc[127]), .D(instrc
		[124]), .Z(n_4200));
	notech_or2 i_29481(.A(n_323160859), .B(instrc[124]), .Z(n_29917));
	notech_or4 i_136436312(.A(temp_sp[28]), .B(temp_sp[29]), .C(temp_sp[31])
		, .D(temp_sp[30]), .Z(n_420582435));
	notech_or4 i_136136315(.A(temp_sp[25]), .B(temp_sp[27]), .C(temp_sp[26])
		, .D(temp_sp[24]), .Z(n_420882437));
	notech_or4 i_135736319(.A(temp_sp[21]), .B(temp_sp[20]), .C(temp_sp[23])
		, .D(temp_sp[22]), .Z(n_4213));
	notech_or4 i_135436322(.A(temp_sp[17]), .B(temp_sp[16]), .C(temp_sp[19])
		, .D(temp_sp[18]), .Z(n_421682442));
	notech_or4 i_136736310(.A(n_421682442), .B(n_4213), .C(n_420882437), .D(n_420582435
		), .Z(n_4219));
	notech_or4 i_134936327(.A(temp_sp[12]), .B(temp_sp[15]), .C(temp_sp[14])
		, .D(temp_sp[13]), .Z(n_422482445));
	notech_or4 i_134636330(.A(temp_sp[8]), .B(temp_sp[9]), .C(temp_sp[11]), 
		.D(temp_sp[10]), .Z(n_4227));
	notech_or4 i_134236334(.A(temp_sp[5]), .B(temp_sp[4]), .C(temp_sp[7]), .D
		(temp_sp[6]), .Z(n_4231));
	notech_or4 i_133936337(.A(temp_sp[1]), .B(temp_sp[3]), .C(temp_sp[2]), .D
		(temp_sp[0]), .Z(n_4234));
	notech_or4 i_135136325(.A(n_4234), .B(n_4231), .C(n_4227), .D(n_422482445
		), .Z(n_4236));
	notech_nand3 i_133536341(.A(n_347671363), .B(n_30381), .C(n_349671381), 
		.Z(n_4238));
	notech_or4 i_132636350(.A(n_19620), .B(n_2039), .C(n_19629), .D(n_30628)
		, .Z(n_4247));
	notech_or4 i_132536351(.A(n_339061018), .B(n_76712523), .C(instrc[127]),
		 .D(instrc[124]), .Z(n_4248));
	notech_ao4 i_129336376(.A(n_4248), .B(n_4466), .C(n_4247), .D(n_412282396
		), .Z(n_4249));
	notech_nand3 i_130936366(.A(n_32506), .B(n_32485), .C(n_19629), .Z(n_4251
		));
	notech_and2 i_74437519(.A(n_4459), .B(n_4128), .Z(n_4254));
	notech_ao3 i_132036356(.A(n_418982430), .B(n_419082431), .C(n_419182432)
		, .Z(n_4257));
	notech_or2 i_131736359(.A(n_57566), .B(tcmp), .Z(n_4259));
	notech_ao4 i_129736374(.A(n_412582399), .B(n_352678529), .C(n_412482398)
		, .D(n_4259), .Z(n_4262));
	notech_ao4 i_129236377(.A(n_339361021), .B(n_57436), .C(n_412382397), .D
		(n_61859), .Z(n_4263));
	notech_ao4 i_129036379(.A(n_61846), .B(n_30560), .C(n_61087), .D(n_30775
		), .Z(n_4265));
	notech_nao3 i_139137493(.A(n_33175), .B(n_33153), .C(instrc[125]), .Z(n_59312350
		));
	notech_and3 i_123536429(.A(n_417382423), .B(n_417582424), .C(n_4174), .Z
		(n_4272));
	notech_nao3 i_124136425(.A(n_33162), .B(\opcode[0] ), .C(n_390364434), .Z
		(n_4276));
	notech_ao4 i_123236432(.A(n_411782391), .B(n_411682390), .C(n_23763), .D
		(n_411582389), .Z(n_4277));
	notech_ao4 i_122936435(.A(n_28572), .B(n_26662), .C(n_26663), .D(n_28581
		), .Z(n_4280));
	notech_ao4 i_122736437(.A(n_26987), .B(n_79112547), .C(n_370864239), .D(n_23741
		), .Z(n_4284));
	notech_and4 i_123136433(.A(n_4284), .B(n_416982420), .C(n_4280), .D(n_30431
		), .Z(n_4286));
	notech_ao4 i_108736562(.A(n_60194), .B(n_340661034), .C(n_4025), .D(n_60159
		), .Z(n_4287));
	notech_ao4 i_108636563(.A(n_27930), .B(n_27843), .C(n_28098), .D(n_25713
		), .Z(n_4288));
	notech_and4 i_108536564(.A(n_4452), .B(n_4402), .C(n_348171367), .D(n_416182412
		), .Z(n_4291));
	notech_nand2 i_109136558(.A(n_30636), .B(read_ack), .Z(n_4292));
	notech_ao4 i_107136577(.A(n_1861), .B(n_4401), .C(n_340561033), .D(n_28008
		), .Z(n_4296));
	notech_ao4 i_102836614(.A(n_32484), .B(n_309271075), .C(n_4085), .D(n_2081
		), .Z(n_4304));
	notech_nao3 i_77236842(.A(n_32506), .B(n_33242), .C(n_32484), .Z(n_4311)
		);
	notech_or2 i_77036844(.A(n_4086), .B(n_30374), .Z(n_4312));
	notech_ao4 i_75336856(.A(write_ack), .B(n_409282386), .C(n_4312), .D(n_4311
		), .Z(n_4313));
	notech_and4 i_76136849(.A(n_4462), .B(n_58664), .C(n_4142), .D(n_4254), 
		.Z(n_4319));
	notech_ao4 i_75236857(.A(n_4095), .B(n_61859), .C(n_4094), .D(n_61845), 
		.Z(n_4322));
	notech_ao3 i_75536854(.A(n_4313), .B(n_4322), .C(n_4141), .Z(n_4323));
	notech_ao4 i_75036859(.A(n_4470), .B(n_30628), .C(n_577), .D(n_2025), .Z
		(n_4324));
	notech_mux2 i_8192286(.S(n_61680), .A(n_1830), .B(n_57749), .Z(n_4327)
		);
	notech_nand2 i_45492287(.A(n_33242), .B(n_59560), .Z(n_4328));
	notech_nao3 i_1330786(.A(n_31474), .B(n_31476), .C(n_4343), .Z(n_4329)
		);
	notech_or4 i_51692288(.A(n_32575), .B(n_32646), .C(n_63800), .D(n_60159)
		, .Z(n_4330));
	notech_or4 i_55492293(.A(n_32575), .B(n_32391), .C(n_63720), .D(n_63732)
		, .Z(n_4335));
	notech_ao4 i_131892295(.A(n_32397), .B(n_28533), .C(n_315460782), .D(n_60159
		), .Z(n_4337));
	notech_and2 i_162492297(.A(n_32485), .B(n_32481), .Z(n_4338));
	notech_nand3 i_149592299(.A(n_61628), .B(n_61087), .C(n_4338), .Z(n_4340
		));
	notech_or4 i_51292302(.A(opd[0]), .B(opd[1]), .C(opd[4]), .D(opd[5]), .Z
		(n_4343));
	notech_nao3 i_51892303(.A(n_63790), .B(n_63700), .C(n_32575), .Z(n_4344)
		);
	notech_ao4 i_51992304(.A(n_349271377), .B(n_4344), .C(n_60177), .D(n_347471362
		), .Z(n_4345));
	notech_nand2 i_3018012(.A(n_208680592), .B(n_208580591), .Z(write_data_26
		[29]));
	notech_nor2 i_55159(.A(n_333681811), .B(n_345881925), .Z(\nbus_11356[6] 
		));
	notech_and2 i_19222(.A(n_62441), .B(n_209680602), .Z(\nbus_11289[8] ));
	notech_ao4 i_3571929(.A(n_348571371), .B(n_4099), .C(n_2025), .D(n_33494
		), .Z(n_239446886));
	notech_and4 i_3671928(.A(n_329281769), .B(n_209280598), .C(n_209180597),
		 .D(n_209380599), .Z(n_239346885));
	notech_ao3 i_95065218(.A(opa[11]), .B(n_29417), .C(n_60194), .Z(n_262367014
		));
	notech_or4 i_88365285(.A(n_63716), .B(n_57387), .C(n_63732), .D(n_58348)
		, .Z(n_262167013));
	notech_or2 i_19069315(.A(n_212980632), .B(n_4347), .Z(\nbus_11309[31] )
		);
	notech_or4 i_7243322(.A(n_125342694), .B(n_384382274), .C(n_3931), .D(n_4425
		), .Z(n_4347));
	notech_or4 i_57369307(.A(n_61723), .B(n_61890), .C(n_2111), .D(nbus_11271
		[31]), .Z(n_24216));
	notech_or4 i_61769306(.A(n_61890), .B(n_61723), .C(n_2111), .D(\nbus_11290[31] 
		), .Z(n_24298));
	notech_nao3 i_88665282(.A(n_30300), .B(\opa_12[15] ), .C(n_376064291), .Z
		(n_261867010));
	notech_or4 i_88965279(.A(n_61940), .B(n_31626), .C(n_30319), .D(n_323578244
		), .Z(n_261567007));
	notech_nand3 i_37058(.A(n_19672), .B(n_61628), .C(n_19637), .Z(n_4348)
		);
	notech_or4 i_37057(.A(n_32396), .B(n_28008), .C(n_60194), .D(n_61628), .Z
		(n_4349));
	notech_or4 i_62243337(.A(n_59120), .B(n_60189), .C(n_32589), .D(n_61628)
		, .Z(n_4350));
	notech_or4 i_61940146(.A(n_32391), .B(n_32394), .C(n_60159), .D(n_61628)
		, .Z(n_24142));
	notech_or4 i_58643334(.A(n_32396), .B(n_59120), .C(n_60189), .D(n_61628)
		, .Z(n_4351));
	notech_or4 i_62343335(.A(n_61890), .B(n_4025), .C(n_61725), .D(n_60159),
		 .Z(n_4352));
	notech_or4 i_62443336(.A(n_32576), .B(n_60175), .C(n_28098), .D(n_61628)
		, .Z(n_4353));
	notech_ao4 i_82643361(.A(n_19672), .B(n_61679), .C(n_111142552), .D(n_59100
		), .Z(n_112042561));
	notech_nor2 i_57843359(.A(n_4424), .B(n_384582276), .Z(n_111142552));
	notech_and2 i_84446462(.A(n_376864299), .B(n_3770), .Z(n_62742068));
	notech_and2 i_84546463(.A(n_377482219), .B(n_376982215), .Z(n_62642067)
		);
	notech_and2 i_82246461(.A(n_379164322), .B(n_29758), .Z(n_62442065));
	notech_and2 i_44946460(.A(n_379264323), .B(n_377382218), .Z(n_62142062)
		);
	notech_or4 i_1021000(.A(n_30917), .B(n_234780848), .C(n_236480865), .D(n_236280863
		), .Z(n_4354));
	notech_nand2 i_820998(.A(n_237880879), .B(n_237280873), .Z(n_4355));
	notech_nand2 i_320993(.A(n_239080891), .B(n_238480885), .Z(n_4356));
	notech_nand2 i_1021064(.A(n_240080901), .B(n_239580896), .Z(n_4357));
	notech_nand2 i_821062(.A(n_241280913), .B(n_240680907), .Z(n_4358));
	notech_nand2 i_321057(.A(n_242680925), .B(n_241880919), .Z(n_4359));
	notech_nand2 i_1021320(.A(n_244680937), .B(n_243680931), .Z(n_4360));
	notech_nand2 i_3121789(.A(n_245780948), .B(n_245280943), .Z(n_4361));
	notech_nand2 i_1021768(.A(n_247180961), .B(n_246480955), .Z(n_436282448)
		);
	notech_nand3 i_153563376(.A(n_247980969), .B(n_30903), .C(n_32273), .Z(n_4364
		));
	notech_nand2 i_620740(.A(n_265981149), .B(n_265481144), .Z(n_4365));
	notech_nand2 i_620836(.A(n_267081160), .B(n_266581155), .Z(n_4366));
	notech_nand2 i_620964(.A(n_268181171), .B(n_267681166), .Z(n_4367));
	notech_nand2 i_220960(.A(n_269181181), .B(n_268681176), .Z(n_4368));
	notech_nand2 i_620996(.A(n_270381193), .B(n_269781187), .Z(n_4369));
	notech_nand2 i_621060(.A(n_271581205), .B(n_270981199), .Z(n_4370));
	notech_or4 i_1021832(.A(n_30917), .B(n_255881048), .C(n_272781212), .D(n_272181210
		), .Z(n_4371));
	notech_nand2 i_821830(.A(n_274781225), .B(n_274181220), .Z(n_4372));
	notech_nand2 i_621828(.A(n_275881236), .B(n_275381231), .Z(n_437382449)
		);
	notech_nand2 i_1017000(.A(n_277081248), .B(n_276481242), .Z(n_4374));
	notech_and4 i_1017576(.A(n_277881256), .B(n_277781255), .C(n_277681254),
		 .D(n_278181259), .Z(n_4375));
	notech_nand2 i_817574(.A(n_279581273), .B(n_278981267), .Z(n_4376));
	notech_nand2 i_617572(.A(n_280881286), .B(n_280281280), .Z(n_4377));
	notech_and4 i_821350(.A(n_291381391), .B(n_291281390), .C(n_292281400), 
		.D(n_291181389), .Z(n_4378));
	notech_nand2 i_621348(.A(n_293581413), .B(n_292981407), .Z(n_4379));
	notech_and4 i_1021896(.A(n_294281420), .B(n_294181419), .C(n_286881346),
		 .D(n_294581423), .Z(n_4380));
	notech_nand2 i_821894(.A(n_295981437), .B(n_295381431), .Z(n_4381));
	notech_and4 i_621892(.A(n_296881446), .B(n_296781445), .C(n_296681444), 
		.D(n_297281450), .Z(n_4382));
	notech_and4 i_517571(.A(n_298281460), .B(n_298181459), .C(n_298081458), 
		.D(n_298681464), .Z(n_4383));
	notech_and4 i_317569(.A(n_299681474), .B(n_299581473), .C(n_299481472), 
		.D(n_300081478), .Z(n_4384));
	notech_or4 i_85265316(.A(n_63716), .B(n_57387), .C(n_63732), .D(n_58321)
		, .Z(n_261067002));
	notech_ao4 i_52755961(.A(n_57656), .B(n_30904), .C(n_30317), .D(n_4443),
		 .Z(n_4386));
	notech_and4 i_145229811(.A(n_317081647), .B(n_316981646), .C(n_316581642
		), .D(n_316881645), .Z(n_4387));
	notech_and4 i_3020764(.A(n_222077272), .B(n_319181668), .C(n_311981596),
		 .D(n_319081667), .Z(n_4388));
	notech_and4 i_3020860(.A(n_222077272), .B(n_319881675), .C(n_311081588),
		 .D(n_319781674), .Z(n_4389));
	notech_and4 i_3020988(.A(n_222077272), .B(n_320581682), .C(n_310281580),
		 .D(n_320481681), .Z(n_4390));
	notech_nand3 i_3021020(.A(n_321381690), .B(n_321281689), .C(n_321181688)
		, .Z(n_4391));
	notech_and4 i_3021180(.A(n_222077272), .B(n_321981696), .C(n_308681564),
		 .D(n_321881695), .Z(n_4392));
	notech_nand2 i_3021340(.A(n_323181708), .B(n_322681703), .Z(n_4393));
	notech_nand2 i_3021788(.A(n_324281719), .B(n_323781714), .Z(n_4394));
	notech_nand2 i_2921787(.A(n_325381730), .B(n_324881725), .Z(n_4395));
	notech_nand2 i_2821786(.A(n_326481741), .B(n_325981736), .Z(n_4396));
	notech_nand2 i_2721785(.A(n_327581752), .B(n_327081747), .Z(n_4397));
	notech_and4 i_3021916(.A(n_328081757), .B(n_328281759), .C(n_301681494),
		 .D(n_327981756), .Z(n_4398));
	notech_and4 i_3017596(.A(n_328481761), .B(n_328681763), .C(n_329181768),
		 .D(n_301281490), .Z(n_4399));
	notech_or4 i_8055846(.A(n_32396), .B(n_59120), .C(n_63700), .D(n_61940),
		 .Z(n_27930));
	notech_and4 i_145129801(.A(n_318481661), .B(n_318381660), .C(n_317981656
		), .D(n_318281659), .Z(n_440082450));
	notech_nor2 i_46829(.A(n_1849), .B(n_28082), .Z(n_365728697));
	notech_and2 i_180653089(.A(n_27920), .B(n_58523), .Z(n_365128691));
	notech_or4 i_77953088(.A(n_32396), .B(n_61846), .C(n_63800), .D(n_309960727
		), .Z(n_364350916));
	notech_and2 i_183653087(.A(n_2033), .B(n_59515), .Z(n_364150918));
	notech_or4 i_31316(.A(n_61725), .B(n_61890), .C(n_4401), .D(n_61859), .Z
		(n_28082));
	notech_nand2 i_11707(.A(pipe_mul[1]), .B(n_30935), .Z(n_4401));
	notech_and3 i_177053084(.A(n_32590), .B(n_1817), .C(n_332081797), .Z(n_363850921
		));
	notech_ao4 i_58053082(.A(n_61846), .B(n_30357), .C(n_60453), .D(n_19548)
		, .Z(n_353728636));
	notech_nao3 i_85565313(.A(n_30300), .B(\opa_12[12] ), .C(n_376064291), .Z
		(n_260666999));
	notech_or4 i_61692306(.A(n_61917), .B(n_61903), .C(n_61890), .D(n_348171367
		), .Z(n_1840));
	notech_and2 i_141237604(.A(n_2112), .B(n_2111), .Z(n_4402));
	notech_or4 i_85865310(.A(n_61940), .B(n_31623), .C(n_30319), .D(n_323578244
		), .Z(n_260366996));
	notech_or4 i_84165327(.A(n_63716), .B(n_57387), .C(n_63732), .D(n_58312)
		, .Z(n_259866991));
	notech_mux2 i_311649(.S(n_61284), .A(n_520), .B(add_len_pc32[2]), .Z(\add_len_pc[2] 
		));
	notech_mux2 i_411650(.S(n_61284), .A(n_521), .B(add_len_pc32[3]), .Z(\add_len_pc[3] 
		));
	notech_mux2 i_511651(.S(n_61284), .A(n_522), .B(add_len_pc32[4]), .Z(\add_len_pc[4] 
		));
	notech_nand2 i_520675(.A(n_366582115), .B(n_365882108), .Z(n_4408));
	notech_nand2 i_420674(.A(n_367982129), .B(n_367282122), .Z(n_4409));
	notech_nand2 i_320673(.A(n_369482143), .B(n_368782136), .Z(n_4410));
	notech_and4 i_421314(.A(n_370682155), .B(n_370582154), .C(n_371082159), 
		.D(n_370482153), .Z(n_4411));
	notech_nand2 i_2021778(.A(n_372282171), .B(n_371782166), .Z(n_4412));
	notech_nand2 i_1921777(.A(n_373382182), .B(n_372882177), .Z(n_4413));
	notech_nand2 i_1821776(.A(n_374482193), .B(n_373982188), .Z(n_4414));
	notech_nand2 i_1721775(.A(n_375582204), .B(n_375082199), .Z(n_4415));
	notech_nand2 i_417570(.A(n_376882214), .B(n_376282210), .Z(n_4416));
	notech_mux2 i_1011656(.S(n_61284), .A(n_527), .B(add_len_pc32[9]), .Z(\add_len_pc[9] 
		));
	notech_nao3 i_29641(.A(instrc[117]), .B(n_286063762), .C(n_62442065), .Z
		(n_4418));
	notech_nor2 i_29642(.A(n_62442065), .B(n_29891), .Z(n_442082451));
	notech_nao3 i_29643(.A(instrc[117]), .B(n_286063762), .C(n_29888), .Z(n_442182452
		));
	notech_nand2 i_1020680(.A(n_3813), .B(n_3807), .Z(n_4422));
	notech_nand2 i_3221790(.A(n_382482255), .B(n_381982250), .Z(n_4423));
	notech_nor2 i_202643364(.A(n_4337), .B(n_61628), .Z(n_4424));
	notech_nao3 i_57543338(.A(n_315760785), .B(n_61628), .C(n_315560783), .Z
		(n_25682));
	notech_nor2 i_5807(.A(n_4432), .B(n_57218), .Z(n_4425));
	notech_and4 i_93929171(.A(n_394582334), .B(n_3944), .C(n_3940), .D(n_3943
		), .Z(n_4427));
	notech_and4 i_94029172(.A(n_3959), .B(n_395882339), .C(n_3954), .D(n_3957
		), .Z(n_4428));
	notech_nand2 i_3016220(.A(n_3977), .B(n_397282345), .Z(n_4429));
	notech_and4 i_1416204(.A(n_398482352), .B(n_398382351), .C(n_3994), .D(n_398282350
		), .Z(n_4430));
	notech_nand3 i_416194(.A(n_4023), .B(n_4014), .C(n_4019), .Z(n_4431));
	notech_and3 i_11143320(.A(n_31604), .B(n_31605), .C(n_31606), .Z(n_4432)
		);
	notech_nao3 i_84465324(.A(n_30300), .B(\opa_12[11] ), .C(n_376064291), .Z
		(n_259566988));
	notech_and4 i_68043307(.A(n_25433), .B(n_397882347), .C(n_386982298), .D
		(n_4000), .Z(n_4433));
	notech_or4 i_74243303(.A(n_61890), .B(n_32397), .C(n_25680), .D(n_61725)
		, .Z(n_61516490));
	notech_ao3 i_74643299(.A(n_383482265), .B(n_382882259), .C(n_30418), .Z(n_4434
		));
	notech_nao3 i_86343292(.A(instrc[107]), .B(n_32243), .C(n_382582256), .Z
		(n_61716492));
	notech_or4 i_95143290(.A(instrc[123]), .B(instrc[121]), .C(n_318160809),
		 .D(n_61816493), .Z(n_58116456));
	notech_or4 i_9397(.A(n_32275), .B(n_318160809), .C(n_61816493), .D(n_4432
		), .Z(n_4435));
	notech_ao4 i_82743293(.A(n_25682), .B(n_30330), .C(n_61816493), .D(n_57412
		), .Z(n_4436));
	notech_ao4 i_55043319(.A(n_316760795), .B(n_61628), .C(n_25649), .D(n_30361
		), .Z(n_4437));
	notech_and2 i_177343278(.A(n_383482265), .B(n_383382264), .Z(n_4438));
	notech_and2 i_75543295(.A(n_61516490), .B(n_397882347), .Z(n_443982453)
		);
	notech_ao4 i_160143294(.A(n_28098), .B(n_339661024), .C(n_4025), .D(n_32397
		), .Z(n_4440));
	notech_and2 i_943323(.A(n_396682342), .B(n_383582266), .Z(n_4441));
	notech_ao3 i_75340141(.A(n_27823), .B(n_30364), .C(n_4086), .Z(n_4442)
		);
	notech_and4 i_161940138(.A(n_27843), .B(n_57656), .C(n_336260990), .D(n_30420
		), .Z(n_4443));
	notech_ao4 i_148340136(.A(n_25670), .B(n_4086), .C(n_57206), .D(n_30701)
		, .Z(n_4444));
	notech_or2 i_165640135(.A(n_4442), .B(n_23845), .Z(n_4445));
	notech_and2 i_78140108(.A(n_406282377), .B(n_4039), .Z(n_23845));
	notech_and2 i_64840134(.A(n_24142), .B(n_4035), .Z(n_4446));
	notech_ao4 i_55540133(.A(n_32590), .B(n_61628), .C(n_4086), .D(n_30364),
		 .Z(n_4447));
	notech_and2 i_139040128(.A(n_406382378), .B(n_4033), .Z(n_4448));
	notech_or2 i_19150(.A(n_23847), .B(opc[3]), .Z(n_444982454));
	notech_and3 i_145440116(.A(n_27843), .B(n_57657), .C(n_336260990), .Z(n_4450
		));
	notech_or4 i_60040111(.A(n_309960727), .B(n_29534), .C(n_32646), .D(n_63800
		), .Z(n_25428));
	notech_or4 i_211140110(.A(n_63818), .B(n_63800), .C(n_32394), .D(n_60159
		), .Z(n_4452));
	notech_or4 i_74140109(.A(n_4086), .B(n_19548), .C(n_27823), .D(n_56930),
		 .Z(n_23847));
	notech_ao4 i_153140107(.A(n_29534), .B(n_32627), .C(n_30701), .D(n_30700
		), .Z(n_4453));
	notech_and4 i_517155(.A(n_4079), .B(n_4078), .C(n_4083), .D(n_407782385)
		, .Z(n_4454));
	notech_or4 i_84765321(.A(n_61940), .B(n_31622), .C(n_30319), .D(n_323578244
		), .Z(n_259266985));
	notech_and4 i_51236(.A(n_331260940), .B(n_4265), .C(n_4263), .D(n_4249),
		 .Z(n_445582455));
	notech_and4 i_48755(.A(n_4277), .B(n_4286), .C(n_4172), .D(n_4272), .Z(n_4456
		));
	notech_and3 i_55160(.A(n_4160), .B(n_415982411), .C(n_4111), .Z(n_4457)
		);
	notech_and4 i_47561(.A(n_2112), .B(n_415482406), .C(n_4467), .D(n_2111),
		 .Z(n_4458));
	notech_or4 i_9808(.A(n_61917), .B(n_61903), .C(n_61890), .D(n_30341), .Z
		(n_4459));
	notech_or4 i_62637704(.A(n_61917), .B(n_61903), .C(n_61890), .D(n_4107),
		 .Z(n_4460));
	notech_or4 i_62037703(.A(n_32383), .B(n_32575), .C(n_60175), .D(n_61628)
		, .Z(n_4461));
	notech_or4 i_74337702(.A(n_314960777), .B(n_28008), .C(n_61630), .D(n_60159
		), .Z(n_4462));
	notech_and3 i_8518(.A(n_61087), .B(n_61679), .C(n_411982393), .Z(n_4463)
		);
	notech_nao3 i_29491(.A(instrc[99]), .B(n_30785), .C(n_30449), .Z(n_4464)
		);
	notech_nand2 i_152637616(.A(n_33164), .B(n_33174), .Z(n_29232));
	notech_and2 i_152937615(.A(n_33160), .B(n_33179), .Z(n_29229));
	notech_or4 i_170737612(.A(n_59560), .B(n_348471370), .C(n_415382405), .D
		(n_2091), .Z(n_4465));
	notech_or2 i_175637607(.A(instrc[125]), .B(n_33175), .Z(n_4466));
	notech_and4 i_194237455(.A(n_415782409), .B(n_4296), .C(n_4090), .D(n_4089
		), .Z(n_4467));
	notech_and4 i_79337601(.A(n_4148), .B(n_4150), .C(n_4304), .D(n_414982402
		), .Z(n_4468));
	notech_and4 i_126938(.A(n_4134), .B(n_4324), .C(n_4471), .D(n_4323), .Z(n_4469
		));
	notech_ao4 i_68337531(.A(read_ack), .B(n_19603), .C(n_71912476), .D(n_324671211
		), .Z(n_4470));
	notech_nao3 i_5879(.A(n_19698), .B(n_4098), .C(n_32484), .Z(n_4471));
	notech_and4 i_33312(.A(n_32506), .B(n_61630), .C(n_61087), .D(n_4338), .Z
		(n_26086));
	notech_and2 i_9892319(.A(n_4327), .B(n_1840), .Z(n_22481));
	notech_and3 i_142192320(.A(n_4330), .B(n_4345), .C(n_4335), .Z(n_22474)
		);
	notech_and4 i_36931(.A(n_32386), .B(n_3455), .C(n_4337), .D(n_1850), .Z(n_22467
		));
	notech_and2 i_159792322(.A(n_30867), .B(n_4328), .Z(n_1830));
	notech_or2 i_75865410(.A(n_444668030), .B(n_3910), .Z(n_258366976));
	notech_or2 i_76565403(.A(n_331760945), .B(n_3610), .Z(n_257766970));
	notech_or2 i_71965449(.A(n_444668030), .B(n_3907), .Z(n_257066963));
	notech_or2 i_72665442(.A(n_331760945), .B(n_3609), .Z(n_256466957));
	notech_or2 i_70565463(.A(n_444668030), .B(n_431067894), .Z(n_255766950)
		);
	notech_or2 i_71265456(.A(n_331760945), .B(n_430767891), .Z(n_255166944)
		);
	notech_or2 i_60565563(.A(n_331660944), .B(n_336160989), .Z(n_253466927)
		);
	notech_or4 i_55465614(.A(n_63716), .B(n_57388), .C(n_63732), .D(n_58348)
		, .Z(n_253366926));
	notech_or2 i_55765611(.A(n_57252), .B(n_33248), .Z(n_253066923));
	notech_or4 i_56065608(.A(n_192776985), .B(n_58279), .C(n_61940), .D(n_31626
		), .Z(n_252766920));
	notech_or4 i_52365645(.A(n_63716), .B(n_57388), .C(n_63732), .D(n_58321)
		, .Z(n_252266915));
	notech_or2 i_52665642(.A(n_57252), .B(n_33250), .Z(n_251966912));
	notech_or4 i_52965639(.A(n_192776985), .B(n_58279), .C(n_61940), .D(n_31623
		), .Z(n_251666909));
	notech_nand2 i_48665679(.A(opb[15]), .B(n_57129), .Z(n_250766900));
	notech_or2 i_49365672(.A(n_3610), .B(n_328860916), .Z(n_250066893));
	notech_nand2 i_45865707(.A(opb[12]), .B(n_57129), .Z(n_249366886));
	notech_or2 i_46565700(.A(n_3609), .B(n_328860916), .Z(n_248666879));
	notech_nand2 i_44465721(.A(opb[11]), .B(n_57129), .Z(n_247966872));
	notech_or2 i_45165714(.A(n_430767891), .B(n_328860916), .Z(n_247266865)
		);
	notech_or2 i_28465873(.A(n_55955), .B(n_30997), .Z(n_245766851));
	notech_or2 i_25665901(.A(n_55955), .B(n_30991), .Z(n_244166836));
	notech_or2 i_24165916(.A(n_55955), .B(n_30989), .Z(n_242466821));
	notech_or2 i_12766030(.A(n_331460942), .B(n_31474), .Z(n_242166819));
	notech_or4 i_13266025(.A(n_332160949), .B(n_61940), .C(nbus_11271[2]), .D
		(n_56003), .Z(n_241666815));
	notech_nor2 i_13766020(.A(n_326460892), .B(n_26272), .Z(n_241166811));
	notech_nor2 i_9666060(.A(n_3690), .B(n_57393), .Z(n_240366803));
	notech_nor2 i_9966057(.A(n_323978248), .B(n_33248), .Z(n_240066800));
	notech_nao3 i_10266054(.A(n_63774), .B(opc_10[15]), .C(n_333978345), .Z(n_239766797
		));
	notech_ao3 i_10366053(.A(opa[15]), .B(n_30351), .C(n_60194), .Z(n_239466794
		));
	notech_nor2 i_7866078(.A(n_368667786), .B(n_57393), .Z(n_239366793));
	notech_nor2 i_8166075(.A(n_323978248), .B(n_33250), .Z(n_239066790));
	notech_nao3 i_8466072(.A(n_63770), .B(opc_10[12]), .C(n_333978345), .Z(n_238766787
		));
	notech_ao3 i_8566071(.A(n_61016), .B(n_30351), .C(n_60196), .Z(n_238466784
		));
	notech_or2 i_128566153(.A(n_439367977), .B(n_28555), .Z(n_28260));
	notech_ao4 i_170567653(.A(n_56411), .B(n_58312), .C(n_61679), .D(n_32603
		), .Z(n_238366783));
	notech_ao4 i_170067658(.A(n_56411), .B(n_58321), .C(n_61679), .D(n_32604
		), .Z(n_238266782));
	notech_ao4 i_168367673(.A(n_56411), .B(n_58348), .C(n_61679), .D(n_32607
		), .Z(n_238166781));
	notech_ao4 i_146667872(.A(n_59114), .B(n_32951), .C(n_56387), .D(n_32953
		), .Z(n_237966779));
	notech_ao4 i_145267886(.A(n_59114), .B(n_32954), .C(n_56387), .D(n_32956
		), .Z(n_237766777));
	notech_ao3 i_119468128(.A(n_213666546), .B(n_213766547), .C(n_237366773)
		, .Z(n_237566775));
	notech_or4 i_119268130(.A(n_213366543), .B(n_213466544), .C(n_213566545)
		, .D(n_237066770), .Z(n_237366773));
	notech_or4 i_118968133(.A(n_213066540), .B(n_30500), .C(n_213166541), .D
		(n_213266542), .Z(n_237066770));
	notech_ao3 i_117468148(.A(n_212566535), .B(n_212666536), .C(n_236466764)
		, .Z(n_236666766));
	notech_or4 i_117268150(.A(n_212266532), .B(n_212366533), .C(n_212466534)
		, .D(n_236166761), .Z(n_236466764));
	notech_or4 i_116968153(.A(n_211966529), .B(n_30498), .C(n_212066530), .D
		(n_212166531), .Z(n_236166761));
	notech_ao3 i_111668206(.A(n_211466524), .B(n_211566525), .C(n_235566755)
		, .Z(n_235766757));
	notech_or4 i_111268208(.A(n_211166521), .B(n_211266522), .C(n_211366523)
		, .D(n_235266752), .Z(n_235566755));
	notech_or4 i_110968211(.A(n_210866518), .B(n_30497), .C(n_210966519), .D
		(n_211066520), .Z(n_235266752));
	notech_ao4 i_99668317(.A(n_327360901), .B(n_28742), .C(n_327160899), .D(n_28743
		), .Z(n_234966749));
	notech_or4 i_99368320(.A(n_210066511), .B(n_209866509), .C(n_234366743),
		 .D(n_209966510), .Z(n_234666746));
	notech_nao3 i_99068323(.A(n_209466506), .B(n_234266742), .C(n_30917), .Z
		(n_234366743));
	notech_ao4 i_98968324(.A(n_28855), .B(n_33168), .C(n_99942440), .D(n_28860
		), .Z(n_234266742));
	notech_ao4 i_97668337(.A(n_28742), .B(n_3753), .C(n_28743), .D(n_3752), 
		.Z(n_234066740));
	notech_or4 i_97268340(.A(n_208766500), .B(n_208566498), .C(n_233466734),
		 .D(n_208666499), .Z(n_233766737));
	notech_nand3 i_96968343(.A(n_233366733), .B(n_208266495), .C(n_310067477
		), .Z(n_233466734));
	notech_ao4 i_96868344(.A(n_28855), .B(n_33258), .C(n_28860), .D(n_431067894
		), .Z(n_233366733));
	notech_ao4 i_95468357(.A(n_28742), .B(n_3689), .C(n_28743), .D(n_3688), 
		.Z(n_233166731));
	notech_or4 i_94768360(.A(n_207166489), .B(n_206966487), .C(n_232566725),
		 .D(n_207066488), .Z(n_232866728));
	notech_nand3 i_94368363(.A(n_232466724), .B(n_206666484), .C(n_310167478
		), .Z(n_232566725));
	notech_ao4 i_94268364(.A(n_28855), .B(n_33250), .C(n_28860), .D(n_3907),
		 .Z(n_232466724));
	notech_ao4 i_88668415(.A(n_28742), .B(n_3693), .C(n_28743), .D(n_3692), 
		.Z(n_2322));
	notech_or4 i_88268418(.A(n_206066478), .B(n_205866476), .C(n_231666717),
		 .D(n_205966477), .Z(n_231966720));
	notech_nand3 i_87968421(.A(n_231566716), .B(n_205566473), .C(n_310267479
		), .Z(n_231666717));
	notech_ao4 i_87668422(.A(n_28855), .B(n_33248), .C(n_28860), .D(n_3910),
		 .Z(n_231566716));
	notech_and4 i_72568566(.A(n_231166712), .B(n_231066711), .C(n_205366471)
		, .D(n_230866709), .Z(n_231366714));
	notech_ao4 i_71968572(.A(n_446068044), .B(n_33258), .C(n_431067894), .D(n_445968043
		), .Z(n_231166712));
	notech_ao4 i_71868573(.A(n_4418), .B(n_3752), .C(n_442182452), .D(n_3751
		), .Z(n_231066711));
	notech_nor2 i_71768574(.A(n_204366462), .B(n_30500), .Z(n_230866709));
	notech_ao4 i_72168570(.A(n_57141), .B(n_433367917), .C(n_62442065), .D(n_3750
		), .Z(n_230666707));
	notech_ao4 i_72068571(.A(n_62642067), .B(n_58312), .C(n_62742068), .D(n_58974
		), .Z(n_230566706));
	notech_and4 i_70568586(.A(n_230266703), .B(n_230166702), .C(n_204166460)
		, .D(n_229966700), .Z(n_230466705));
	notech_ao4 i_69968592(.A(n_446068044), .B(n_33250), .C(n_3907), .D(n_445968043
		), .Z(n_230266703));
	notech_ao4 i_69868593(.A(n_4418), .B(n_3688), .C(n_442182452), .D(n_368767787
		), .Z(n_230166702));
	notech_nor2 i_69768594(.A(n_203166451), .B(n_30498), .Z(n_229966700));
	notech_ao4 i_70168590(.A(n_57141), .B(n_309867475), .C(n_62442065), .D(n_368667786
		), .Z(n_229766698));
	notech_ao4 i_70068591(.A(n_62642067), .B(n_58321), .C(n_62742068), .D(n_59050
		), .Z(n_229666697));
	notech_and4 i_64768644(.A(n_229366694), .B(n_229266693), .C(n_202966449)
		, .D(n_229066691), .Z(n_229566696));
	notech_ao4 i_64168650(.A(n_446068044), .B(n_33248), .C(n_3910), .D(n_445968043
		), .Z(n_229366694));
	notech_ao4 i_64068651(.A(n_4418), .B(n_3692), .C(n_442182452), .D(n_3691
		), .Z(n_229266693));
	notech_nor2 i_63968652(.A(n_202066440), .B(n_30497), .Z(n_229066691));
	notech_ao4 i_64368648(.A(n_57141), .B(n_309967476), .C(n_62442065), .D(n_3690
		), .Z(n_228866689));
	notech_ao4 i_64268649(.A(n_62642067), .B(n_58348), .C(n_62742068), .D(n_59068
		), .Z(n_228766688));
	notech_nand3 i_62568666(.A(n_228266683), .B(n_201566435), .C(n_201666436
		), .Z(n_228466685));
	notech_and4 i_62368668(.A(n_327860906), .B(n_201066432), .C(n_201466434)
		, .D(n_201166433), .Z(n_228266683));
	notech_and4 i_53368755(.A(n_227766678), .B(n_227666677), .C(n_200166426)
		, .D(n_227466675), .Z(n_227966680));
	notech_ao4 i_52768761(.A(n_304744481), .B(n_33168), .C(n_99942440), .D(n_304644480
		), .Z(n_227766678));
	notech_ao4 i_52668762(.A(n_327160899), .B(n_30075), .C(n_327260900), .D(n_30078
		), .Z(n_227666677));
	notech_nor2 i_52568763(.A(n_199066417), .B(n_30917), .Z(n_227466675));
	notech_ao4 i_52968759(.A(n_57122), .B(n_326960897), .C(n_327060898), .D(n_72542166
		), .Z(n_227266673));
	notech_ao4 i_52868760(.A(n_72742168), .B(n_58294), .C(n_4924), .D(n_59032
		), .Z(n_227166672));
	notech_and4 i_51368775(.A(n_226866669), .B(n_226766668), .C(n_198866415)
		, .D(n_226566666), .Z(n_227066671));
	notech_ao4 i_50768781(.A(n_304744481), .B(n_33258), .C(n_304644480), .D(n_431067894
		), .Z(n_226866669));
	notech_ao4 i_50668782(.A(n_30075), .B(n_3752), .C(n_30078), .D(n_3751), 
		.Z(n_226766668));
	notech_nor2 i_50568783(.A(n_197966406), .B(n_30500), .Z(n_226566666));
	notech_ao4 i_50968779(.A(n_57122), .B(n_433367917), .C(n_72542166), .D(n_3750
		), .Z(n_226366664));
	notech_ao4 i_50868780(.A(n_72742168), .B(n_58312), .C(n_4924), .D(n_58974
		), .Z(n_226266663));
	notech_and4 i_49368795(.A(n_225966660), .B(n_225866659), .C(n_197766404)
		, .D(n_225666657), .Z(n_226166662));
	notech_ao4 i_48768801(.A(n_304744481), .B(n_33250), .C(n_304644480), .D(n_3907
		), .Z(n_225966660));
	notech_ao4 i_48668802(.A(n_30075), .B(n_3688), .C(n_30078), .D(n_368767787
		), .Z(n_225866659));
	notech_nor2 i_48568803(.A(n_196866395), .B(n_30498), .Z(n_225666657));
	notech_ao4 i_48968799(.A(n_57122), .B(n_309867475), .C(n_72542166), .D(n_368667786
		), .Z(n_225466655));
	notech_ao4 i_48868800(.A(n_72742168), .B(n_58321), .C(n_4924), .D(n_59050
		), .Z(n_225366654));
	notech_and4 i_42968853(.A(n_225066651), .B(n_224966650), .C(n_196666393)
		, .D(n_224766648), .Z(n_225266653));
	notech_ao4 i_42368859(.A(n_304744481), .B(n_33248), .C(n_304644480), .D(n_3910
		), .Z(n_225066651));
	notech_ao4 i_42268860(.A(n_30075), .B(n_3692), .C(n_30078), .D(n_3691), 
		.Z(n_224966650));
	notech_nor2 i_42168861(.A(n_195766384), .B(n_30497), .Z(n_224766648));
	notech_ao4 i_42568857(.A(n_57122), .B(n_309967476), .C(n_72542166), .D(n_3690
		), .Z(n_224566646));
	notech_ao4 i_42468858(.A(n_72742168), .B(n_58348), .C(n_4924), .D(n_59068
		), .Z(n_224466645));
	notech_ao3 i_40868874(.A(n_224066641), .B(n_195366380), .C(n_195466381),
		 .Z(n_224266643));
	notech_and4 i_40668876(.A(n_327860906), .B(n_194966376), .C(n_223866639)
		, .D(n_195266379), .Z(n_224066641));
	notech_ao4 i_40468878(.A(n_323960867), .B(n_33169), .C(n_101142452), .D(n_323860866
		), .Z(n_223866639));
	notech_nand3 i_38568895(.A(n_193966366), .B(n_223166632), .C(n_194266369
		), .Z(n_223366634));
	notech_ao3 i_38268898(.A(n_222966630), .B(n_193766364), .C(n_193866365),
		 .Z(n_223166632));
	notech_and4 i_38068900(.A(n_222766628), .B(n_193666363), .C(n_326860896)
		, .D(n_193366360), .Z(n_222966630));
	notech_ao4 i_37868902(.A(n_323960867), .B(n_33167), .C(n_100842449), .D(n_323860866
		), .Z(n_222766628));
	notech_ao4 i_38468896(.A(n_326360891), .B(n_30391), .C(n_326760895), .D(n_30390
		), .Z(n_222566626));
	notech_nand3 i_36168919(.A(n_192666353), .B(n_222066621), .C(n_192966356
		), .Z(n_222266623));
	notech_ao3 i_35868922(.A(n_221866619), .B(n_192466351), .C(n_192566352),
		 .Z(n_222066621));
	notech_and4 i_35668924(.A(n_221666617), .B(n_192366350), .C(n_325860886)
		, .D(n_192066347), .Z(n_221866619));
	notech_ao4 i_35468926(.A(n_323960867), .B(n_33166), .C(n_100542446), .D(n_323860866
		), .Z(n_221666617));
	notech_ao4 i_36068920(.A(n_325360881), .B(n_30391), .C(n_325760885), .D(n_30390
		), .Z(n_221466615));
	notech_and4 i_31568965(.A(n_221166612), .B(n_221066611), .C(n_191766344)
		, .D(n_220866609), .Z(n_221366614));
	notech_ao4 i_30968971(.A(n_442168005), .B(n_33168), .C(n_99942440), .D(n_442268006
		), .Z(n_221166612));
	notech_ao4 i_30868972(.A(n_327160899), .B(n_445668040), .C(n_327260900),
		 .D(n_445868042), .Z(n_221066611));
	notech_and2 i_30768973(.A(n_327460902), .B(n_190866335), .Z(n_220866609)
		);
	notech_ao4 i_31168969(.A(n_326960897), .B(n_57170), .C(n_91142352), .D(n_327060898
		), .Z(n_220666607));
	notech_ao4 i_31068970(.A(n_91442355), .B(n_58294), .C(n_91542356), .D(n_59032
		), .Z(n_220566606));
	notech_and4 i_27369005(.A(n_220266603), .B(n_220166602), .C(n_219966600)
		, .D(n_190666333), .Z(n_220466605));
	notech_ao4 i_26569011(.A(n_442168005), .B(n_33258), .C(n_431067894), .D(n_442268006
		), .Z(n_220266603));
	notech_ao4 i_26469012(.A(n_445668040), .B(n_3752), .C(n_445868042), .D(n_3751
		), .Z(n_220166602));
	notech_and2 i_26369013(.A(n_189766324), .B(n_310067477), .Z(n_219966600)
		);
	notech_ao4 i_26869009(.A(n_57170), .B(n_433367917), .C(n_91142352), .D(n_3750
		), .Z(n_219766598));
	notech_ao4 i_26669010(.A(n_91442355), .B(n_58312), .C(n_91542356), .D(n_58974
		), .Z(n_219666597));
	notech_and4 i_24869025(.A(n_219366594), .B(n_219266593), .C(n_219066591)
		, .D(n_189566322), .Z(n_219566596));
	notech_ao4 i_24169031(.A(n_442168005), .B(n_33250), .C(n_3907), .D(n_442268006
		), .Z(n_219366594));
	notech_ao4 i_24069032(.A(n_445668040), .B(n_3688), .C(n_445868042), .D(n_368767787
		), .Z(n_219266593));
	notech_and2 i_23969033(.A(n_188666313), .B(n_310167478), .Z(n_219066591)
		);
	notech_ao4 i_24369029(.A(n_57170), .B(n_309867475), .C(n_91142352), .D(n_368667786
		), .Z(n_218866589));
	notech_ao4 i_24269030(.A(n_91442355), .B(n_58321), .C(n_91542356), .D(n_59050
		), .Z(n_218766588));
	notech_ao4 i_20369068(.A(n_31487), .B(n_90742348), .C(n_377064301), .D(n_57170
		), .Z(n_218466585));
	notech_ao4 i_20269069(.A(n_91542356), .B(\nbus_11290[14] ), .C(n_442168005
		), .D(n_33215), .Z(n_218366584));
	notech_and3 i_20469067(.A(n_218166582), .B(n_377364304), .C(n_187866305)
		, .Z(n_218266583));
	notech_ao4 i_20069070(.A(n_97342414), .B(n_442268006), .C(n_377164302), 
		.D(n_445668040), .Z(n_218166582));
	notech_and4 i_18269083(.A(n_217666578), .B(n_217566577), .C(n_217266575)
		, .D(n_187366300), .Z(n_217966580));
	notech_ao4 i_17669089(.A(n_442168005), .B(n_33248), .C(n_3910), .D(n_442268006
		), .Z(n_217666578));
	notech_ao4 i_17569090(.A(n_445668040), .B(n_3692), .C(n_445868042), .D(n_3691
		), .Z(n_217566577));
	notech_and2 i_17469091(.A(n_186466291), .B(n_310267479), .Z(n_217266575)
		);
	notech_ao4 i_17869087(.A(n_57170), .B(n_309967476), .C(n_91142352), .D(n_3690
		), .Z(n_217066573));
	notech_ao4 i_17769088(.A(n_91442355), .B(n_58348), .C(n_91542356), .D(n_59068
		), .Z(n_216966572));
	notech_nand2 i_1227351(.A(n_238366783), .B(n_216566568), .Z(n_216866571)
		);
	notech_nao3 i_170467654(.A(n_3499), .B(n_60605), .C(n_56428), .Z(n_216566568
		));
	notech_nand2 i_1327352(.A(n_238266782), .B(n_215866564), .Z(n_216466567)
		);
	notech_nao3 i_169967659(.A(n_3500), .B(n_60605), .C(n_56428), .Z(n_215866564
		));
	notech_nand2 i_1627355(.A(n_238166781), .B(n_215366560), .Z(n_215766563)
		);
	notech_nao3 i_168267674(.A(n_3503), .B(n_60605), .C(n_56428), .Z(n_215366560
		));
	notech_nand3 i_1327480(.A(n_237966779), .B(n_215166558), .C(n_214566555)
		, .Z(n_215266559));
	notech_or2 i_146467874(.A(n_309892426), .B(n_59050), .Z(n_215166558));
	notech_nao3 i_146567873(.A(n_3564), .B(opb[31]), .C(n_56428), .Z(n_214566555
		));
	notech_nand3 i_1627483(.A(n_237766777), .B(n_214366553), .C(n_214066550)
		, .Z(n_214466554));
	notech_or2 i_145067888(.A(n_309892426), .B(n_59068), .Z(n_214366553));
	notech_nao3 i_145167887(.A(n_3567), .B(opb[31]), .C(n_56429), .Z(n_214066550
		));
	notech_nand3 i_1221610(.A(n_213866548), .B(n_237566775), .C(n_212966539)
		, .Z(n_213966549));
	notech_or2 i_118368139(.A(n_26935), .B(n_33258), .Z(n_213866548));
	notech_nand2 i_118168141(.A(n_30522), .B(opa[11]), .Z(n_213766547));
	notech_or4 i_118268140(.A(n_162262654), .B(n_57407), .C(n_26951), .D(n_431067894
		), .Z(n_213666546));
	notech_and3 i_118468138(.A(n_63770), .B(opc[11]), .C(n_26823), .Z(n_213566545
		));
	notech_ao3 i_118668136(.A(opa[11]), .B(n_26822), .C(n_60196), .Z(n_213466544
		));
	notech_nor2 i_117968143(.A(n_303844472), .B(n_3750), .Z(n_213366543));
	notech_ao3 i_118568137(.A(n_63790), .B(opc_10[11]), .C(n_26821), .Z(n_213266542
		));
	notech_and2 i_117868144(.A(n_305144485), .B(opd[11]), .Z(n_213166541));
	notech_nor2 i_117768145(.A(n_57091), .B(n_433367917), .Z(n_213066540));
	notech_nand2 i_118068142(.A(n_30523), .B(opb[11]), .Z(n_212966539));
	notech_nand3 i_1321611(.A(n_212766537), .B(n_236666766), .C(n_211866528)
		, .Z(n_212866538));
	notech_or2 i_116368159(.A(n_26935), .B(n_33250), .Z(n_212766537));
	notech_nand2 i_116168161(.A(n_30522), .B(opa[12]), .Z(n_212666536));
	notech_or4 i_116268160(.A(n_162262654), .B(n_57407), .C(n_26951), .D(n_3907
		), .Z(n_212566535));
	notech_and3 i_116468158(.A(n_63770), .B(opc[12]), .C(n_26823), .Z(n_212466534
		));
	notech_ao3 i_116668156(.A(opa[12]), .B(n_26822), .C(n_60196), .Z(n_212366533
		));
	notech_nor2 i_115968163(.A(n_303844472), .B(n_368667786), .Z(n_212266532
		));
	notech_ao3 i_116568157(.A(n_63768), .B(opc_10[12]), .C(n_26821), .Z(n_212166531
		));
	notech_and2 i_115868164(.A(n_305144485), .B(opd[12]), .Z(n_212066530));
	notech_nor2 i_115768165(.A(n_57091), .B(n_309867475), .Z(n_211966529));
	notech_nand2 i_116068162(.A(n_30523), .B(opb[12]), .Z(n_211866528));
	notech_nand3 i_1621614(.A(n_211666526), .B(n_235766757), .C(n_210766517)
		, .Z(n_211766527));
	notech_or2 i_110368217(.A(n_26935), .B(n_33248), .Z(n_211666526));
	notech_nand2 i_110168219(.A(n_30522), .B(opa[15]), .Z(n_211566525));
	notech_or4 i_110268218(.A(n_162262654), .B(n_57407), .C(n_26951), .D(n_3910
		), .Z(n_211466524));
	notech_and3 i_110468216(.A(n_63770), .B(opc[15]), .C(n_26823), .Z(n_211366523
		));
	notech_ao3 i_110668214(.A(opa[15]), .B(n_26822), .C(n_60196), .Z(n_211266522
		));
	notech_nor2 i_109968221(.A(n_303844472), .B(n_3690), .Z(n_211166521));
	notech_ao3 i_110568215(.A(n_63770), .B(opc_10[15]), .C(n_26821), .Z(n_211066520
		));
	notech_and2 i_109868222(.A(n_305144485), .B(opd[15]), .Z(n_210966519));
	notech_nor2 i_109768223(.A(n_57091), .B(n_309967476), .Z(n_210866518));
	notech_nand2 i_110068220(.A(n_30523), .B(opb[15]), .Z(n_210766517));
	notech_or4 i_1021160(.A(n_210166512), .B(n_234666746), .C(n_210266513), 
		.D(n_30575), .Z(n_210666516));
	notech_nor2 i_98468329(.A(n_302944463), .B(n_58294), .Z(n_210266513));
	notech_and2 i_98368330(.A(opb[9]), .B(n_30631), .Z(n_210166512));
	notech_nor2 i_98268331(.A(n_327060898), .B(n_303744471), .Z(n_210066511)
		);
	notech_and2 i_98168332(.A(n_305044484), .B(opd[9]), .Z(n_209966510));
	notech_ao3 i_98668327(.A(n_63792), .B(opc_10[9]), .C(n_28741), .Z(n_209866509
		));
	notech_or4 i_97868335(.A(n_336660994), .B(n_30719), .C(n_340361031), .D(n_32217
		), .Z(n_209466506));
	notech_or4 i_1221162(.A(n_208866501), .B(n_233766737), .C(n_209066502), 
		.D(n_30580), .Z(n_209366505));
	notech_nor2 i_96368349(.A(n_302944463), .B(n_58312), .Z(n_209066502));
	notech_and2 i_96268350(.A(n_30631), .B(opb[11]), .Z(n_208866501));
	notech_nor2 i_96168351(.A(n_303744471), .B(n_3750), .Z(n_208766500));
	notech_and2 i_96068352(.A(n_305044484), .B(opd[11]), .Z(n_208666499));
	notech_ao3 i_96568347(.A(n_63770), .B(opc_10[11]), .C(n_28741), .Z(n_208566498
		));
	notech_or2 i_95668355(.A(n_57195), .B(n_433367917), .Z(n_208266495));
	notech_or4 i_1321163(.A(n_207266490), .B(n_232866728), .C(n_207766491), 
		.D(n_30583), .Z(n_208066494));
	notech_nor2 i_93568369(.A(n_302944463), .B(n_58321), .Z(n_207766491));
	notech_and2 i_93468370(.A(n_30631), .B(opb[12]), .Z(n_207266490));
	notech_nor2 i_93368371(.A(n_303744471), .B(n_368667786), .Z(n_207166489)
		);
	notech_and2 i_93268372(.A(n_305044484), .B(opd[12]), .Z(n_207066488));
	notech_ao3 i_93768367(.A(n_63770), .B(opc_10[12]), .C(n_28741), .Z(n_206966487
		));
	notech_or2 i_92968375(.A(n_57195), .B(n_309867475), .Z(n_206666484));
	notech_or4 i_1621166(.A(n_206166479), .B(n_231966720), .C(n_206266480), 
		.D(n_30586), .Z(n_206566483));
	notech_nor2 i_87068427(.A(n_302944463), .B(nbus_11273[15]), .Z(n_206266480
		));
	notech_and2 i_86968428(.A(n_30631), .B(opb[15]), .Z(n_206166479));
	notech_nor2 i_86868429(.A(n_303744471), .B(n_3690), .Z(n_206066478));
	notech_and2 i_86768430(.A(n_305044484), .B(opd[15]), .Z(n_205966477));
	notech_ao3 i_87368425(.A(n_63792), .B(opc_10[15]), .C(n_28741), .Z(n_205866476
		));
	notech_or2 i_86368433(.A(n_57195), .B(n_309967476), .Z(n_205566473));
	notech_nand3 i_1220970(.A(n_230666707), .B(n_230566706), .C(n_231366714)
		, .Z(n_205466472));
	notech_or2 i_71668575(.A(n_62142062), .B(n_31484), .Z(n_205366471));
	notech_ao3 i_70768584(.A(opa[11]), .B(n_442082451), .C(n_60196), .Z(n_204366462
		));
	notech_nand3 i_1320971(.A(n_229766698), .B(n_229666697), .C(n_230466705)
		, .Z(n_204266461));
	notech_or2 i_69668595(.A(n_62142062), .B(n_31485), .Z(n_204166460));
	notech_ao3 i_68768604(.A(opa[12]), .B(n_442082451), .C(n_60196), .Z(n_203166451
		));
	notech_nand3 i_1620974(.A(n_228866689), .B(n_228766688), .C(n_229566696)
		, .Z(n_203066450));
	notech_or2 i_63868653(.A(n_62142062), .B(n_31488), .Z(n_202966449));
	notech_ao3 i_62968662(.A(opa[15]), .B(n_442082451), .C(n_60196), .Z(n_202066440
		));
	notech_or4 i_120831(.A(n_201766437), .B(n_228466685), .C(n_201866438), .D
		(n_200866430), .Z(n_201966439));
	notech_ao3 i_61468676(.A(n_30483), .B(\opa_12[0] ), .C(n_304344477), .Z(n_201866438
		));
	notech_and2 i_61968672(.A(opb[0]), .B(n_200766429), .Z(n_201766437));
	notech_nao3 i_61668674(.A(n_63792), .B(opc[0]), .C(n_29994), .Z(n_201666436
		));
	notech_or2 i_61568675(.A(n_30196), .B(n_101142452), .Z(n_201566435));
	notech_nao3 i_61868673(.A(n_30212), .B(n_30483), .C(n_327760905), .Z(n_201466434
		));
	notech_or2 i_61368677(.A(n_305244486), .B(n_31472), .Z(n_201166433));
	notech_or2 i_61268678(.A(n_57122), .B(n_327560903), .Z(n_201066432));
	notech_ao4 i_61068680(.A(n_304244476), .B(n_33214), .C(n_30077), .D(n_30428
		), .Z(n_200966431));
	notech_and2 i_62068671(.A(n_200966431), .B(opa[0]), .Z(n_200866430));
	notech_nand2 i_60968681(.A(n_304644480), .B(n_291167288), .Z(n_200766429
		));
	notech_nand3 i_1020840(.A(n_227266673), .B(n_227166672), .C(n_227966680)
		, .Z(n_200266427));
	notech_or2 i_52468764(.A(n_4922), .B(n_31482), .Z(n_200166426));
	notech_ao3 i_51568773(.A(n_61007), .B(n_30076), .C(n_60196), .Z(n_199066417
		));
	notech_nand3 i_1220842(.A(n_226366664), .B(n_226266663), .C(n_227066671)
		, .Z(n_198966416));
	notech_or2 i_50468784(.A(n_4922), .B(n_31484), .Z(n_198866415));
	notech_ao3 i_49568793(.A(opa[11]), .B(n_30076), .C(n_60196), .Z(n_197966406
		));
	notech_nand3 i_1320843(.A(n_225466655), .B(n_225366654), .C(n_226166662)
		, .Z(n_197866405));
	notech_or2 i_48468804(.A(n_4922), .B(n_31485), .Z(n_197766404));
	notech_ao3 i_47568813(.A(opa[12]), .B(n_30076), .C(n_60196), .Z(n_196866395
		));
	notech_nand3 i_1620846(.A(n_224566646), .B(n_224466645), .C(n_225266653)
		, .Z(n_196766394));
	notech_or2 i_42068862(.A(n_4922), .B(n_31488), .Z(n_196666393));
	notech_ao3 i_41168871(.A(opa[15]), .B(n_30076), .C(n_60196), .Z(n_195766384
		));
	notech_nand3 i_120735(.A(n_195566382), .B(n_224266643), .C(n_194666373),
		 .Z(n_195666383));
	notech_nand2 i_39968883(.A(n_194566372), .B(opa[0]), .Z(n_195566382));
	notech_and4 i_40168881(.A(n_323660864), .B(n_63758), .C(opc[0]), .D(n_30515
		), .Z(n_195466381));
	notech_nand2 i_39768885(.A(opd[0]), .B(n_30630), .Z(n_195366380));
	notech_nao3 i_39868884(.A(n_63792), .B(opc_10[0]), .C(n_30393), .Z(n_195266379
		));
	notech_or2 i_39368888(.A(n_327560903), .B(n_57168), .Z(n_194966376));
	notech_nor2 i_86169351(.A(n_3608), .B(n_30429), .Z(n_194866375));
	notech_nand2 i_39268889(.A(n_442268006), .B(n_292067297), .Z(n_194766374
		));
	notech_nand2 i_40068882(.A(opb[0]), .B(n_194766374), .Z(n_194666373));
	notech_ao4 i_39068891(.A(n_32697), .B(n_31327), .C(n_3608), .D(n_30429),
		 .Z(n_194566372));
	notech_or4 i_320737(.A(n_194366370), .B(n_193266359), .C(n_223366634), .D
		(n_30607), .Z(n_194466371));
	notech_ao3 i_37268908(.A(n_30395), .B(n_32266), .C(n_326560893), .Z(n_194366370
		));
	notech_or4 i_37068910(.A(n_60196), .B(n_323660864), .C(n_303944473), .D(nbus_11273
		[2]), .Z(n_194266369));
	notech_or4 i_37168909(.A(n_60175), .B(n_303944473), .C(nbus_11273[2]), .D
		(n_32266), .Z(n_193966366));
	notech_nor2 i_36968911(.A(n_326160889), .B(n_303944473), .Z(n_193866365)
		);
	notech_nand2 i_36868912(.A(opd[2]), .B(n_30630), .Z(n_193766364));
	notech_nao3 i_37568905(.A(n_63770), .B(opc_10[2]), .C(n_30393), .Z(n_193666363
		));
	notech_or2 i_36568915(.A(n_326060888), .B(n_57164), .Z(n_193366360));
	notech_ao3 i_37668904(.A(n_30395), .B(n_57517), .C(n_326460892), .Z(n_193266359
		));
	notech_or4 i_720741(.A(n_193066357), .B(n_191966346), .C(n_222266623), .D
		(n_30608), .Z(n_193166358));
	notech_ao3 i_34868932(.A(n_30395), .B(n_32266), .C(n_325560883), .Z(n_193066357
		));
	notech_or4 i_34668934(.A(n_63716), .B(n_61938), .C(nbus_11273[6]), .D(n_30578
		), .Z(n_192966356));
	notech_or4 i_34768933(.A(n_60177), .B(n_303944473), .C(nbus_11273[6]), .D
		(n_32266), .Z(n_192666353));
	notech_nor2 i_34568935(.A(n_325160879), .B(n_303944473), .Z(n_192566352)
		);
	notech_nand2 i_34468936(.A(opd[6]), .B(n_30630), .Z(n_192466351));
	notech_nao3 i_35168929(.A(n_63792), .B(opc_10[6]), .C(n_30393), .Z(n_192366350
		));
	notech_or2 i_34168939(.A(n_325060878), .B(n_57164), .Z(n_192066347));
	notech_ao3 i_35268928(.A(n_30395), .B(n_57512), .C(n_325460882), .Z(n_191966346
		));
	notech_nand3 i_1020744(.A(n_220666607), .B(n_220566606), .C(n_221366614)
		, .Z(n_191866345));
	notech_or2 i_30668974(.A(n_90742348), .B(n_31482), .Z(n_191766344));
	notech_or4 i_29768983(.A(n_63716), .B(n_445768041), .C(n_61938), .D(n_58294
		), .Z(n_190866335));
	notech_nand3 i_1220746(.A(n_219766598), .B(n_219666597), .C(n_220466605)
		, .Z(n_190766334));
	notech_or2 i_26269014(.A(n_90742348), .B(n_31484), .Z(n_190666333));
	notech_or4 i_25169023(.A(n_91142352), .B(n_323660864), .C(n_60196), .D(n_58312
		), .Z(n_189766324));
	notech_nand3 i_1320747(.A(n_218866589), .B(n_218766588), .C(n_219566596)
		, .Z(n_189666323));
	notech_or2 i_23869034(.A(n_90742348), .B(n_31485), .Z(n_189566322));
	notech_or4 i_22969043(.A(n_91142352), .B(n_323660864), .C(n_60194), .D(n_58321
		), .Z(n_188666313));
	notech_and4 i_1520749(.A(n_218466585), .B(n_218366584), .C(n_218266583),
		 .D(n_187666303), .Z(n_188566312));
	notech_nao3 i_18669079(.A(n_63740), .B(opc_10[14]), .C(n_445868042), .Z(n_187866305
		));
	notech_ao4 i_18469081(.A(n_32697), .B(n_31327), .C(n_3608), .D(n_30484),
		 .Z(n_187766304));
	notech_nand2 i_19769072(.A(n_187766304), .B(opa[14]), .Z(n_187666303));
	notech_nand3 i_1620750(.A(n_217066573), .B(n_216966572), .C(n_217966580)
		, .Z(n_187466301));
	notech_or2 i_17369092(.A(n_90742348), .B(n_31488), .Z(n_187366300));
	notech_or4 i_16469101(.A(n_91142352), .B(n_323660864), .C(n_60194), .D(n_58348
		), .Z(n_186466291));
	notech_or4 i_54576(.A(n_61917), .B(n_61903), .C(n_316160789), .D(n_177266204
		), .Z(n_186266289));
	notech_ao4 i_31371667(.A(n_30823), .B(n_57524), .C(n_30786), .D(n_58279)
		, .Z(n_185966286));
	notech_or4 i_22513(.A(n_177166203), .B(n_177066202), .C(n_176966201), .D
		(n_176866200), .Z(n_185866285));
	notech_or4 i_32371657(.A(n_2580), .B(n_32159), .C(n_32161), .D(n_1850), 
		.Z(n_184766277));
	notech_nao3 i_1571949(.A(instrc[124]), .B(n_180666238), .C(tcmp), .Z(n_184666276
		));
	notech_nand2 i_4471920(.A(n_436867952), .B(n_31249), .Z(n_184166271));
	notech_and4 i_21671763(.A(n_183166263), .B(n_183466266), .C(n_176466196)
		, .D(n_176166193), .Z(n_183866268));
	notech_ao4 i_21471765(.A(n_183366265), .B(n_30923), .C(n_174866184), .D(n_3594
		), .Z(n_183466266));
	notech_nand3 i_21171768(.A(n_33164), .B(instrc[104]), .C(instrc[107]), .Z
		(n_183366265));
	notech_ao4 i_21271767(.A(n_111445606), .B(n_57489), .C(n_57136), .D(n_114845640
		), .Z(n_183166263));
	notech_or4 i_18271786(.A(n_32484), .B(instrc[102]), .C(n_61680), .D(n_33142
		), .Z(n_183066262));
	notech_nao3 i_18671782(.A(instrc[89]), .B(instrc[91]), .C(n_30334), .Z(n_182966261
		));
	notech_or4 i_17271796(.A(n_182366255), .B(n_173566173), .C(n_173466172),
		 .D(n_30620), .Z(n_182666258));
	notech_ao4 i_16971799(.A(n_375564286), .B(n_30234), .C(n_30240), .D(n_30266
		), .Z(n_182466256));
	notech_or4 i_16871800(.A(n_30621), .B(n_172566167), .C(n_172666168), .D(n_30623
		), .Z(n_182366255));
	notech_ao4 i_16571803(.A(n_30257), .B(n_338661014), .C(n_57164), .D(n_114845640
		), .Z(n_181966251));
	notech_or4 i_13771830(.A(n_170666150), .B(n_170766151), .C(n_170866152),
		 .D(n_181166243), .Z(n_181466246));
	notech_or4 i_13471833(.A(n_312671105), .B(n_170466148), .C(n_170566149),
		 .D(n_30670), .Z(n_181166243));
	notech_and3 i_127871960(.A(instrc[125]), .B(instrc[127]), .C(instrc[126]
		), .Z(n_180666238));
	notech_nao3 i_11271852(.A(n_179966231), .B(n_169066134), .C(n_169166135)
		, .Z(n_180266234));
	notech_ao4 i_10271862(.A(n_30823), .B(n_57444), .C(n_30815), .D(n_3345),
		 .Z(n_179966231));
	notech_ao3 i_54649(.A(n_30614), .B(n_30520), .C(n_179666228), .Z(n_179766229
		));
	notech_ao3 i_34171639(.A(n_32514), .B(n_30377), .C(n_186266289), .Z(n_179666228
		));
	notech_and3 i_34071640(.A(n_19680), .B(n_30650), .C(eval_flag), .Z(n_179566227
		));
	notech_or2 i_5671908(.A(n_339461022), .B(n_250947001), .Z(n_179466226)
		);
	notech_nand3 i_33871642(.A(n_242146913), .B(n_240546897), .C(n_179466226
		), .Z(n_179366225));
	notech_and4 i_33271648(.A(n_56747), .B(n_178766219), .C(n_178866220), .D
		(n_178966221), .Z(n_179266224));
	notech_nao3 i_33371647(.A(n_180666238), .B(n_322360851), .C(n_56766), .Z
		(n_178966221));
	notech_nand3 i_33171649(.A(n_57638), .B(n_63730), .C(n_30315), .Z(n_178866220
		));
	notech_or4 i_32971651(.A(n_32323), .B(n_30904), .C(n_61938), .D(n_58279)
		, .Z(n_178766219));
	notech_nand2 i_32571655(.A(eval_flag), .B(n_178266214), .Z(n_178666218)
		);
	notech_ao3 i_32471656(.A(n_32388), .B(eval_flag), .C(n_60194), .Z(n_178566217
		));
	notech_ao4 i_32071660(.A(tcmp), .B(n_184766277), .C(n_178066212), .D(n_184666276
		), .Z(n_178466216));
	notech_or2 i_32671654(.A(eval_flag), .B(n_178466216), .Z(n_178366215));
	notech_nao3 i_31971661(.A(n_3457), .B(n_1850), .C(n_1854), .Z(n_178266214
		));
	notech_ao4 i_5771907(.A(n_60196), .B(n_30305), .C(n_32397), .D(n_32390),
		 .Z(n_178066212));
	notech_nao3 i_3971925(.A(instrc[104]), .B(instrc[106]), .C(n_3347), .Z(n_177666208
		));
	notech_nao3 i_1371951(.A(n_180666238), .B(instrc[124]), .C(n_30839), .Z(n_177366205
		));
	notech_and4 i_31271668(.A(n_185966286), .B(n_177666208), .C(n_177366205)
		, .D(n_30613), .Z(n_177266204));
	notech_ao3 i_30771673(.A(instrc[90]), .B(instrc[88]), .C(n_3346), .Z(n_177166203
		));
	notech_ao3 i_30571675(.A(instrc[98]), .B(instrc[97]), .C(n_159462626), .Z
		(n_177066202));
	notech_ao3 i_30871672(.A(instrc[102]), .B(instrc[103]), .C(n_1462), .Z(n_176966201
		));
	notech_ao3 i_30671674(.A(instrc[94]), .B(instrc[92]), .C(n_3345), .Z(n_176866200
		));
	notech_and4 i_53512(.A(n_183866268), .B(n_176566197), .C(n_176666198), .D
		(n_30632), .Z(n_176766199));
	notech_nand3 i_20871771(.A(instrc[117]), .B(n_286063762), .C(n_175166187
		), .Z(n_176666198));
	notech_or2 i_20671772(.A(n_1460), .B(n_175066186), .Z(n_176566197));
	notech_nao3 i_20271773(.A(n_32481), .B(n_32353), .C(n_174966185), .Z(n_176466196
		));
	notech_or4 i_19971775(.A(n_323160859), .B(n_30552), .C(n_33162), .D(n_33153
		), .Z(n_176166193));
	notech_ao4 i_20971770(.A(n_241746909), .B(n_174766183), .C(n_174066176),
		 .D(n_29890), .Z(n_175266188));
	notech_nao3 i_18771781(.A(n_323060858), .B(n_174666182), .C(n_322960857)
		, .Z(n_175166187));
	notech_ao4 i_18371785(.A(n_159662628), .B(n_182966261), .C(n_159562627),
		 .D(n_3345), .Z(n_175066186));
	notech_ao4 i_17971789(.A(n_183066262), .B(n_1462), .C(n_29572), .D(n_159462626
		), .Z(n_174966185));
	notech_ao4 i_17771791(.A(n_57638), .B(n_2810), .C(n_30798), .D(n_32224),
		 .Z(n_174866184));
	notech_ao4 i_19071778(.A(n_321860846), .B(n_30547), .C(n_340461032), .D(n_339561023
		), .Z(n_174766183));
	notech_nand3 i_18871780(.A(n_321860846), .B(n_57130), .C(n_63730), .Z(n_174666182
		));
	notech_ao3 i_17571793(.A(n_322360851), .B(n_30344), .C(n_3402), .Z(n_174066176
		));
	notech_ao3 i_54018(.A(n_173666174), .B(n_30619), .C(n_172066162), .Z(n_173966175
		));
	notech_nand3 i_16171807(.A(n_339961027), .B(n_30727), .C(n_171966161), .Z
		(n_173666174));
	notech_and4 i_15571812(.A(instrc[94]), .B(instrc[92]), .C(n_30869), .D(n_30666
		), .Z(n_173566173));
	notech_ao3 i_15371814(.A(n_30869), .B(n_143360301), .C(n_375364284), .Z(n_173466172
		));
	notech_or4 i_16371805(.A(n_322660854), .B(n_1460), .C(n_30751), .D(n_33139
		), .Z(n_172766169));
	notech_ao3 i_16071808(.A(n_55831), .B(n_63730), .C(n_171866160), .Z(n_172666168
		));
	notech_nor2 i_15471813(.A(n_30249), .B(n_30248), .Z(n_172566167));
	notech_ao4 i_16271806(.A(n_241746909), .B(n_171766159), .C(n_171466156),
		 .D(n_30725), .Z(n_172066162));
	notech_nao3 i_14871819(.A(n_323060858), .B(n_171666158), .C(n_322960857)
		, .Z(n_171966161));
	notech_ao4 i_14671821(.A(n_57638), .B(n_2810), .C(n_30798), .D(n_32220),
		 .Z(n_171866160));
	notech_ao4 i_15171816(.A(n_321860846), .B(n_30547), .C(n_339561023), .D(n_2829
		), .Z(n_171766159));
	notech_nand3 i_14971818(.A(n_321860846), .B(n_57164), .C(n_63730), .Z(n_171666158
		));
	notech_ao3 i_14471823(.A(n_322360851), .B(n_30436), .C(n_30266), .Z(n_171466156
		));
	notech_or4 i_54249(.A(n_170966153), .B(n_171066154), .C(n_170266146), .D
		(n_181466246), .Z(n_171366155));
	notech_ao4 i_13071836(.A(n_241746909), .B(n_169566139), .C(n_168666130),
		 .D(n_30308), .Z(n_171066154));
	notech_and4 i_12971837(.A(instrc[119]), .B(instrc[118]), .C(n_56820), .D
		(n_169966143), .Z(n_170966153));
	notech_and3 i_12871838(.A(n_61087), .B(n_61680), .C(n_169866142), .Z(n_170866152
		));
	notech_ao3 i_12771839(.A(n_63794), .B(n_58274), .C(n_169766141), .Z(n_170766151
		));
	notech_ao3 i_12671840(.A(n_30869), .B(n_32481), .C(n_30867), .Z(n_170666150
		));
	notech_and2 i_12371841(.A(fepc), .B(n_61859), .Z(n_170566149));
	notech_nor2 i_12271842(.A(n_114845640), .B(n_57097), .Z(n_170466148));
	notech_or4 i_12171843(.A(n_169466138), .B(n_169366137), .C(n_169666140),
		 .D(n_180266234), .Z(n_170366147));
	notech_and4 i_13171835(.A(n_30869), .B(n_32481), .C(n_32353), .D(n_170366147
		), .Z(n_170266146));
	notech_nao3 i_11071854(.A(n_323060858), .B(n_169266136), .C(n_322960857)
		, .Z(n_169966143));
	notech_nand3 i_10971855(.A(n_349871383), .B(n_32181), .C(n_57019), .Z(n_169866142
		));
	notech_ao4 i_10071864(.A(n_57638), .B(n_2810), .C(n_30798), .D(n_32311),
		 .Z(n_169766141));
	notech_ao3 i_12071844(.A(n_180666238), .B(n_33162), .C(n_30839), .Z(n_169666140
		));
	notech_ao4 i_11871846(.A(n_321860846), .B(n_30547), .C(instrc[112]), .D(n_2821
		), .Z(n_169566139));
	notech_and4 i_11571849(.A(instrc[98]), .B(instrc[97]), .C(instrc[99]), .D
		(n_436767951), .Z(n_169466138));
	notech_nor2 i_11471850(.A(n_30835), .B(n_3347), .Z(n_169366137));
	notech_nand3 i_11171853(.A(n_321860846), .B(n_57097), .C(n_63730), .Z(n_169266136
		));
	notech_and4 i_10771857(.A(instrc[102]), .B(instrc[101]), .C(instrc[103])
		, .D(n_30450), .Z(n_169166135));
	notech_nao3 i_10671858(.A(instrc[90]), .B(n_33160), .C(n_3346), .Z(n_169066134
		));
	notech_ao3 i_9771867(.A(n_180666238), .B(n_436567949), .C(n_57521), .Z(n_168666130
		));
	notech_ao4 i_132973208(.A(n_3910), .B(n_292192264), .C(n_292292265), .D(n_31309
		), .Z(n_168566129));
	notech_ao4 i_133073207(.A(n_293792280), .B(n_31276), .C(n_57436), .D(n_30997
		), .Z(n_168466128));
	notech_ao4 i_133573202(.A(n_3907), .B(n_292192264), .C(n_292292265), .D(n_31306
		), .Z(n_168366127));
	notech_ao4 i_133673201(.A(n_293792280), .B(n_31273), .C(n_57436), .D(n_30991
		), .Z(n_168266126));
	notech_ao4 i_133773200(.A(n_431067894), .B(n_292192264), .C(n_292292265)
		, .D(n_31305), .Z(n_168166125));
	notech_ao4 i_133873199(.A(n_293792280), .B(n_31272), .C(n_57436), .D(n_30989
		), .Z(n_168066124));
	notech_ao4 i_137373164(.A(n_30744), .B(n_31018), .C(n_28747367), .D(n_31286
		), .Z(n_167966123));
	notech_ao4 i_137473163(.A(n_29047370), .B(n_33172), .C(n_29347373), .D(n_31319
		), .Z(n_167866122));
	notech_or4 i_63674523(.A(n_30842), .B(n_30552), .C(n_33153), .D(instrc[
		124]), .Z(n_28747367));
	notech_or2 i_66674517(.A(n_165766101), .B(n_340261030), .Z(n_29047370)
		);
	notech_or4 i_16586(.A(instrc[125]), .B(n_33153), .C(n_33175), .D(n_340261030
		), .Z(n_29347373));
	notech_nand2 i_574496(.A(n_4466), .B(instrc[124]), .Z(n_167466118));
	notech_and4 i_59873918(.A(n_37407), .B(n_79112547), .C(n_167466118), .D(instrc
		[127]), .Z(n_165766101));
	notech_ao3 i_8684466(.A(nbus_11273[3]), .B(nbus_11273[4]), .C(n_27833), 
		.Z(n_27831));
	notech_or4 i_100584465(.A(n_32663), .B(n_2952), .C(n_30899), .D(n_30901)
		, .Z(n_32575));
	notech_or4 i_130784463(.A(opa[0]), .B(opa[1]), .C(opa[2]), .D(opa[3]), .Z
		(n_27832));
	notech_nand3 i_125684461(.A(nbus_11273[0]), .B(nbus_11273[1]), .C(nbus_11273
		[2]), .Z(n_27833));
	notech_nand2 i_121784460(.A(nbus_11273[0]), .B(n_58229), .Z(n_27834));
	notech_nao3 i_26825(.A(n_32646), .B(n_63800), .C(n_61797), .Z(n_32573)
		);
	notech_nand2 i_1421772(.A(n_374564276), .B(n_373964270), .Z(n_391564446)
		);
	notech_or4 i_212584456(.A(n_60177), .B(n_32646), .C(n_63800), .D(n_32394
		), .Z(n_391464445));
	notech_or4 i_212184455(.A(n_32391), .B(n_63730), .C(n_61959), .D(n_32394
		), .Z(n_391364444));
	notech_or2 i_147537596(.A(n_390364434), .B(n_390464435), .Z(n_391264443)
		);
	notech_or4 i_146237597(.A(n_32275), .B(n_32250), .C(n_365964190), .D(n_390464435
		), .Z(n_391164442));
	notech_ao4 i_27537598(.A(n_30719), .B(n_32342), .C(n_57679), .D(n_32314)
		, .Z(n_23760));
	notech_or4 i_54237599(.A(instrc[119]), .B(instrc[118]), .C(instrc[117]),
		 .D(instrc[116]), .Z(n_23763));
	notech_ao4 i_25537600(.A(n_30316), .B(n_32342), .C(n_32314), .D(n_57638)
		, .Z(n_391064441));
	notech_and2 i_32337605(.A(n_390164432), .B(n_390264433), .Z(n_25094));
	notech_or2 i_117237613(.A(instrc[125]), .B(instrc[126]), .Z(n_79112547)
		);
	notech_or4 i_185737625(.A(n_60196), .B(n_32576), .C(n_32628), .D(n_32184
		), .Z(n_32181));
	notech_nand3 i_31737547(.A(n_61087), .B(n_61630), .C(n_30524), .Z(n_32195
		));
	notech_or2 i_120437691(.A(n_26618), .B(n_26398), .Z(n_390964440));
	notech_nao3 i_120537692(.A(n_57436), .B(n_30903), .C(n_26398), .Z(n_390864439
		));
	notech_nor2 i_7255(.A(n_390364434), .B(n_23759), .Z(n_390664437));
	notech_or4 i_7253(.A(n_32275), .B(n_32250), .C(n_365964190), .D(n_23759)
		, .Z(n_390564436));
	notech_ao4 i_26537759(.A(n_30723), .B(n_32342), .C(n_32314), .D(n_57657)
		, .Z(n_390464435));
	notech_and2 i_182037498(.A(n_372964260), .B(n_60159), .Z(n_390364434));
	notech_nao3 i_62537775(.A(n_30367), .B(n_316260790), .C(n_61890), .Z(n_390264433
		));
	notech_or4 i_57037776(.A(n_61917), .B(n_61903), .C(n_61890), .D(n_391464445
		), .Z(n_390164432));
	notech_or4 i_40037780(.A(instrc[113]), .B(instrc[114]), .C(n_2830), .D(n_30316
		), .Z(n_390064431));
	notech_and4 i_50056(.A(n_371864249), .B(n_372064251), .C(n_371664247), .D
		(n_369464225), .Z(n_389964430));
	notech_ao3 i_149040075(.A(nbus_11273[4]), .B(nbus_11273[5]), .C(n_27832)
		, .Z(n_105014667));
	notech_and2 i_176840067(.A(nbus_11273[6]), .B(n_105014667), .Z(n_27829)
		);
	notech_nand2 i_20879(.A(n_58225), .B(opa[0]), .Z(n_389864429));
	notech_nand2 i_20877(.A(nbus_11273[4]), .B(nbus_11273[3]), .Z(n_389764428
		));
	notech_and4 i_1116201(.A(n_364564176), .B(n_364464175), .C(n_365564186),
		 .D(n_364364174), .Z(n_389664427));
	notech_and3 i_98643288(.A(n_61959), .B(n_63758), .C(n_61680), .Z(n_25665
		));
	notech_or4 i_3221630(.A(n_293885352), .B(n_332463896), .C(n_352764059), 
		.D(n_30677), .Z(n_389564426));
	notech_nand2 i_1120681(.A(n_352364055), .B(n_351764049), .Z(n_389464425)
		);
	notech_nand2 i_1420684(.A(n_351164043), .B(n_350564037), .Z(n_389364424)
		);
	notech_mux2 i_1411660(.S(n_61284), .A(n_531), .B(add_len_pc32[13]), .Z(\add_len_pc[13] 
		));
	notech_mux2 i_1111657(.S(n_61286), .A(n_528), .B(add_len_pc32[10]), .Z(\add_len_pc[10] 
		));
	notech_nand2 i_421602(.A(n_3289), .B(n_3284), .Z(n_389064421));
	notech_or4 i_1721615(.A(n_264585062), .B(n_3147), .C(n_3273), .D(n_30702
		), .Z(n_388964420));
	notech_or4 i_1821616(.A(n_263485051), .B(n_3155), .C(n_3259), .D(n_30703
		), .Z(n_388864419));
	notech_or4 i_1921617(.A(n_262385040), .B(n_3164), .C(n_3247), .D(n_30704
		), .Z(n_388764418));
	notech_or4 i_2021618(.A(n_261285029), .B(n_3172), .C(n_3240), .D(n_30705
		), .Z(n_388664417));
	notech_nand2 i_421154(.A(n_3233), .B(n_3226), .Z(n_388564416));
	notech_or4 i_2021170(.A(n_261285029), .B(n_3193), .C(n_3210), .D(n_30706
		), .Z(n_388464415));
	notech_ao3 i_115346476(.A(n_3295), .B(n_28855), .C(n_3296), .Z(n_388364414
		));
	notech_and3 i_115446477(.A(n_3294), .B(n_3293), .C(n_28860), .Z(n_388264413
		));
	notech_and2 i_112849782(.A(n_58664), .B(n_3133), .Z(n_131426641));
	notech_ao3 i_114549772(.A(n_23747), .B(n_391264443), .C(n_390664437), .Z
		(n_131526642));
	notech_and3 i_114649771(.A(n_390564436), .B(n_23750), .C(n_391164442), .Z
		(n_131626643));
	notech_or2 i_132549730(.A(n_3132), .B(n_23763), .Z(n_388164412));
	notech_or4 i_35656(.A(instrc[113]), .B(instrc[114]), .C(n_2830), .D(n_57251
		), .Z(n_388064411));
	notech_or4 i_129437746(.A(n_32275), .B(n_365964190), .C(n_391064441), .D
		(n_32250), .Z(n_387964410));
	notech_or2 i_129837747(.A(n_391064441), .B(n_390364434), .Z(n_387864409)
		);
	notech_nao3 i_132849728(.A(instrc[116]), .B(n_188662913), .C(n_3130), .Z
		(n_387764408));
	notech_or2 i_32466(.A(n_57251), .B(n_57091), .Z(n_387664407));
	notech_nao3 i_1749708(.A(n_26957), .B(n_63758), .C(n_164562677), .Z(n_387564406
		));
	notech_or4 i_1153057(.A(instrc[115]), .B(instrc[112]), .C(n_340461032), 
		.D(n_57256), .Z(n_25090));
	notech_nand3 i_1053058(.A(n_63744), .B(n_25121), .C(n_382064351), .Z(n_25110
		));
	notech_and4 i_117553090(.A(n_385664387), .B(n_256963516), .C(n_382864359
		), .D(n_30697), .Z(n_365228692));
	notech_and4 i_117453091(.A(n_385864389), .B(n_2570), .C(n_382664357), .D
		(n_30689), .Z(n_365328693));
	notech_and3 i_114453092(.A(n_385464385), .B(n_257363519), .C(n_383064361
		), .Z(n_365428694));
	notech_and3 i_113053093(.A(n_58664), .B(n_30693), .C(n_383464365), .Z(n_365528695
		));
	notech_and2 i_112953094(.A(n_30695), .B(n_30640), .Z(n_365628696));
	notech_and3 i_5155875(.A(nbus_11273[6]), .B(n_105014667), .C(nbus_11273[
		7]), .Z(n_96629667));
	notech_or4 i_2721625(.A(n_30574), .B(n_286963771), .C(n_295563853), .D(n_30716
		), .Z(n_387464405));
	notech_or4 i_2821626(.A(n_217484594), .B(n_287763778), .C(n_294863846), 
		.D(n_30717), .Z(n_387364404));
	notech_or4 i_2921627(.A(n_288563786), .B(n_216384583), .C(n_294163839), 
		.D(n_30718), .Z(n_387264403));
	notech_and4 i_3021628(.A(n_222077272), .B(n_293563833), .C(n_289363794),
		 .D(n_293463832), .Z(n_387164402));
	notech_or2 i_6455862(.A(n_30368), .B(n_27835), .Z(n_27827));
	notech_nand3 i_81455934(.A(n_57544), .B(n_386664397), .C(n_286763769), .Z
		(n_29419));
	notech_or4 i_54855916(.A(n_292663824), .B(n_292363821), .C(n_291963817),
		 .D(n_291663814), .Z(n_27798));
	notech_or4 i_87955980(.A(n_318060808), .B(n_2577), .C(n_286263764), .D(n_386764398
		), .Z(n_29540));
	notech_and2 i_97255977(.A(n_60159), .B(n_290763807), .Z(n_386964400));
	notech_or2 i_87055984(.A(n_386964400), .B(n_386764398), .Z(n_29550));
	notech_or4 i_39155989(.A(n_61823), .B(n_30309), .C(n_57638), .D(n_57057)
		, .Z(n_386864399));
	notech_ao4 i_28455991(.A(n_30719), .B(n_32211), .C(n_57679), .D(n_32314)
		, .Z(n_29560));
	notech_ao4 i_27455993(.A(n_30723), .B(n_32211), .C(n_32314), .D(n_57657)
		, .Z(n_386764398));
	notech_ao4 i_26455995(.A(n_32211), .B(n_30316), .C(n_32314), .D(n_57638)
		, .Z(n_386664397));
	notech_ao4 i_25455996(.A(n_30721), .B(n_32211), .C(n_32314), .D(n_30698)
		, .Z(n_29553));
	notech_and2 i_43755987(.A(n_386864399), .B(n_286363765), .Z(n_386464395)
		);
	notech_and4 i_110846497(.A(n_116342604), .B(n_391064441), .C(n_23759), .D
		(n_366264193), .Z(n_386364394));
	notech_and2 i_44346496(.A(n_390064431), .B(n_3311), .Z(n_386264393));
	notech_and2 i_126346498(.A(n_391164442), .B(n_335260980), .Z(n_386164392
		));
	notech_and2 i_126446499(.A(n_335160979), .B(n_3312), .Z(n_386064391));
	notech_or4 i_149660662(.A(n_32269), .B(n_384764378), .C(n_384964380), .D
		(instrc[120]), .Z(n_385864389));
	notech_nand2 i_150560664(.A(n_382964360), .B(n_30504), .Z(n_385664387)
		);
	notech_nand2 i_149160666(.A(n_30504), .B(n_25121), .Z(n_385464385));
	notech_and4 i_143729646(.A(n_349464028), .B(n_349364027), .C(n_348964023
		), .D(n_349264026), .Z(n_385364384));
	notech_or4 i_39960693(.A(instrc[113]), .B(instrc[114]), .C(n_2845), .D(n_32308
		), .Z(n_385264383));
	notech_or4 i_32260694(.A(n_60196), .B(n_32383), .C(n_61797), .D(n_61630)
		, .Z(n_385164382));
	notech_ao4 i_29460700(.A(n_32308), .B(n_32204), .C(n_2848), .D(n_57638),
		 .Z(n_385064381));
	notech_ao4 i_27660701(.A(n_57553), .B(n_32219), .C(n_57679), .D(n_32314)
		, .Z(n_384964380));
	notech_ao4 i_24660704(.A(n_30721), .B(n_32219), .C(n_32314), .D(n_30698)
		, .Z(n_384864379));
	notech_ao4 i_96060670(.A(n_63776), .B(n_61959), .C(n_32397), .D(n_25121)
		, .Z(n_384764378));
	notech_nor2 i_7360705(.A(n_384764378), .B(n_58597), .Z(n_91234596));
	notech_and4 i_1117577(.A(n_285263754), .B(n_285163753), .C(n_285063752),
		 .D(n_285563757), .Z(n_384664377));
	notech_and4 i_1121897(.A(n_284063742), .B(n_283963741), .C(n_260663549),
		 .D(n_284363745), .Z(n_384564376));
	notech_and4 i_1421900(.A(n_282963731), .B(n_282863730), .C(n_261763559),
		 .D(n_283263734), .Z(n_384464375));
	notech_or4 i_1121833(.A(n_262863569), .B(n_282163723), .C(n_30734), .D(n_30735
		), .Z(n_384364374));
	notech_nand2 i_521603(.A(n_281263714), .B(n_280763709), .Z(n_384264373)
		);
	notech_nand2 i_521155(.A(n_280163703), .B(n_279663699), .Z(n_384164372)
		);
	notech_or4 i_1121161(.A(n_266163600), .B(n_30747), .C(n_278863692), .D(n_30740
		), .Z(n_384064371));
	notech_nand2 i_520995(.A(n_278163685), .B(n_277563679), .Z(n_383964370)
		);
	notech_or4 i_1121001(.A(n_268663623), .B(n_30747), .C(n_2767), .D(n_30745
		), .Z(n_383864369));
	notech_or4 i_1120841(.A(n_269663633), .B(n_30747), .C(n_2758), .D(n_30746
		), .Z(n_383764368));
	notech_ao4 i_28660715(.A(n_32290), .B(n_32204), .C(n_2848), .D(n_30698),
		 .Z(n_87434558));
	notech_ao3 i_179660668(.A(n_28557), .B(n_33152), .C(instrc[118]), .Z(n_25121
		));
	notech_nand3 i_32537660(.A(n_61091), .B(n_61630), .C(n_19680), .Z(n_32186
		));
	notech_nao3 i_120160724(.A(n_58574), .B(n_30647), .C(n_256463511), .Z(n_383564366
		));
	notech_nao3 i_8868(.A(n_382064351), .B(n_58601), .C(n_384764378), .Z(n_383464365
		));
	notech_ao4 i_29060714(.A(n_32288), .B(n_32204), .C(n_57679), .D(n_2848),
		 .Z(n_24733));
	notech_and2 i_198960733(.A(n_382064351), .B(n_382964360), .Z(n_383364364
		));
	notech_or4 i_195660734(.A(n_30368), .B(n_27835), .C(n_26028), .D(n_27798
		), .Z(n_383264363));
	notech_or4 i_189060735(.A(instrc[123]), .B(instrc[121]), .C(n_318160809)
		, .D(n_256763514), .Z(n_24735));
	notech_and2 i_182260737(.A(n_273763668), .B(n_60159), .Z(n_383164362));
	notech_nand2 i_147860742(.A(n_30495), .B(n_25121), .Z(n_383064361));
	notech_nand2 i_1360706(.A(n_273063661), .B(n_60159), .Z(n_382964360));
	notech_nand2 i_147660743(.A(n_382964360), .B(n_30495), .Z(n_382864359)
		);
	notech_ao4 i_26660702(.A(n_30723), .B(n_32219), .C(n_32314), .D(n_57657)
		, .Z(n_382764358));
	notech_or4 i_146560746(.A(n_32269), .B(n_384764378), .C(instrc[120]), .D
		(n_382764358), .Z(n_382664357));
	notech_nao3 i_120060725(.A(n_32241), .B(n_30647), .C(n_256463511), .Z(n_382564356
		));
	notech_or4 i_39860777(.A(instrc[115]), .B(instrc[112]), .C(n_58716), .D(n_30316
		), .Z(n_382264353));
	notech_nand3 i_38760779(.A(n_335960987), .B(n_61091), .C(n_61680), .Z(n_382164352
		));
	notech_nand2 i_25660789(.A(n_258463528), .B(n_116542606), .Z(n_382064351
		));
	notech_nand3 i_24160790(.A(n_336560993), .B(n_61091), .C(n_61680), .Z(n_381964350
		));
	notech_or4 i_6730375(.A(opa[7]), .B(n_30270), .C(n_27835), .D(n_27798), 
		.Z(n_381864349));
	notech_and3 i_138360747(.A(n_382164352), .B(n_383564366), .C(n_272463655
		), .Z(n_381764348));
	notech_and3 i_138260748(.A(n_381964350), .B(n_379564326), .C(n_382564356
		), .Z(n_381664347));
	notech_ao3 i_111060765(.A(n_328560913), .B(n_256463511), .C(n_258063525)
		, .Z(n_381564346));
	notech_ao4 i_123460757(.A(n_335660984), .B(n_273463665), .C(n_24733), .D
		(n_383164362), .Z(n_381464345));
	notech_ao4 i_123360758(.A(n_57672), .B(n_273363664), .C(n_24733), .D(n_24735
		), .Z(n_381364344));
	notech_ao3 i_45460770(.A(n_385264383), .B(n_24717), .C(n_2583), .Z(n_381264343
		));
	notech_ao3 i_43963406(.A(n_385264383), .B(n_24716), .C(n_2583), .Z(n_381164342
		));
	notech_and2 i_123163384(.A(n_379464325), .B(n_332360951), .Z(n_381064341
		));
	notech_and2 i_123263383(.A(n_379564326), .B(n_332660954), .Z(n_380964340
		));
	notech_and2 i_197055965(.A(n_290663806), .B(instrc[117]), .Z(n_29557));
	notech_ao4 i_29860717(.A(n_32292), .B(n_32204), .C(n_2848), .D(n_57657),
		 .Z(n_380864339));
	notech_and2 i_106563390(.A(n_24733), .B(n_256463511), .Z(n_380764338));
	notech_or4 i_54460716(.A(instrc[119]), .B(instrc[118]), .C(n_57696), .D(n_33152
		), .Z(n_24736));
	notech_and4 i_816998(.A(n_255663503), .B(n_255563502), .C(n_256063507), 
		.D(n_255463501), .Z(n_380664337));
	notech_nand2 i_1117001(.A(n_254663493), .B(n_254063487), .Z(n_380564336)
		);
	notech_nand2 i_1417004(.A(n_253363480), .B(n_252763474), .Z(n_380464335)
		);
	notech_and4 i_1421836(.A(n_251663463), .B(n_251563462), .C(n_239563392),
		 .D(n_251963466), .Z(n_380364334));
	notech_nand2 i_221600(.A(n_251063457), .B(n_250563453), .Z(n_380264333)
		);
	notech_nand2 i_621604(.A(n_250063448), .B(n_249563443), .Z(n_380164332)
		);
	notech_or4 i_3121629(.A(n_2428), .B(n_170584161), .C(n_248663434), .D(n_30750
		), .Z(n_380064331));
	notech_nand2 i_221152(.A(n_248263430), .B(n_247763425), .Z(n_379964330)
		);
	notech_nand2 i_621156(.A(n_2472), .B(n_2467), .Z(n_379864329));
	notech_or4 i_50260769(.A(instrc[113]), .B(instrc[114]), .C(n_2845), .D(n_32292
		), .Z(n_24717));
	notech_and3 i_81363362(.A(n_57544), .B(n_379064321), .C(n_234763344), .Z
		(n_29758));
	notech_and2 i_100863363(.A(n_32259), .B(n_30658), .Z(n_29890));
	notech_or4 i_201560731(.A(n_32275), .B(n_318160809), .C(n_380864339), .D
		(n_256763514), .Z(n_379564326));
	notech_or2 i_201860730(.A(n_383164362), .B(n_380864339), .Z(n_379464325)
		);
	notech_and2 i_97363395(.A(n_2460), .B(n_60159), .Z(n_379364324));
	notech_or4 i_50760713(.A(instrc[113]), .B(instrc[114]), .C(n_2845), .D(n_32288
		), .Z(n_24716));
	notech_or4 i_39063410(.A(n_61823), .B(n_30309), .C(n_57637), .D(n_57130)
		, .Z(n_379264323));
	notech_ao4 i_28163414(.A(n_57553), .B(n_32224), .C(n_57672), .D(n_32314)
		, .Z(n_29888));
	notech_ao4 i_27163415(.A(n_30723), .B(n_32224), .C(n_57566), .D(n_57657)
		, .Z(n_379164322));
	notech_ao4 i_26163416(.A(n_32224), .B(n_30316), .C(n_57562), .D(n_57633)
		, .Z(n_379064321));
	notech_ao4 i_25163417(.A(n_30721), .B(n_32224), .C(n_57562), .D(n_30698)
		, .Z(n_29887));
	notech_ao3 i_11963418(.A(n_30727), .B(n_57696), .C(instrc[118]), .Z(n_29891
		));
	notech_ao4 i_124037723(.A(n_335660984), .B(n_273463665), .C(n_338061008)
		, .D(n_329360921), .Z(n_378964320));
	notech_ao4 i_123937722(.A(n_57672), .B(n_273363664), .C(n_338061008), .D
		(n_26618), .Z(n_378864319));
	notech_and3 i_138637724(.A(n_382164352), .B(n_390864439), .C(n_368764218
		), .Z(n_378764318));
	notech_and4 i_138737725(.A(n_381964350), .B(n_331260940), .C(n_390964440
		), .D(n_332560953), .Z(n_378664317));
	notech_ao3 i_111637721(.A(n_26398), .B(n_328560913), .C(n_276660615), .Z
		(n_378564316));
	notech_and3 i_44137720(.A(n_337861006), .B(n_26603), .C(n_275360602), .Z
		(n_378464315));
	notech_nor2 i_81855985(.A(n_29419), .B(n_30282), .Z(n_378364314));
	notech_nand2 i_1121769(.A(n_232363320), .B(n_231663314), .Z(n_378264313)
		);
	notech_nand2 i_1121513(.A(n_230963308), .B(n_230363302), .Z(n_378164312)
		);
	notech_nand2 i_1421516(.A(n_229763296), .B(n_229163290), .Z(n_378064311)
		);
	notech_nand2 i_1121353(.A(n_228563284), .B(n_228063279), .Z(n_377964310)
		);
	notech_and4 i_1421356(.A(n_227263271), .B(n_227463273), .C(n_227163270),
		 .D(n_216963169), .Z(n_377864309));
	notech_nand2 i_1121321(.A(n_226663265), .B(n_226063259), .Z(n_377764308)
		);
	notech_nand2 i_1421324(.A(n_225463253), .B(n_224863247), .Z(n_377664307)
		);
	notech_nand2 i_1121065(.A(n_224263241), .B(n_223763236), .Z(n_377564306)
		);
	notech_or4 i_1421004(.A(n_221463213), .B(n_30559), .C(n_223063229), .D(n_222863227
		), .Z(n_377464305));
	notech_or4 i_42655988(.A(n_32184), .B(n_29534), .C(\opcode[0] ), .D(n_61824
		), .Z(n_29533));
	notech_and2 i_43463407(.A(n_379264323), .B(n_234363340), .Z(n_54741988)
		);
	notech_and2 i_81763400(.A(n_29758), .B(n_29888), .Z(n_94542386));
	notech_and4 i_92543352(.A(n_363764168), .B(n_363664167), .C(n_363264163)
		, .D(n_363564166), .Z(n_97342414));
	notech_or4 i_45471526(.A(n_61892), .B(n_113283588), .C(n_61725), .D(n_61859
		), .Z(n_113183587));
	notech_and4 i_45271528(.A(n_1804), .B(n_1803), .C(n_1801), .D(n_1802), .Z
		(n_113283588));
	notech_or4 i_45371527(.A(n_4401), .B(n_1861), .C(n_61861), .D(n_61630), 
		.Z(n_113383589));
	notech_and4 i_52439(.A(n_344281909), .B(n_113383589), .C(n_341381880), .D
		(n_113183587), .Z(\nbus_11337[16] ));
	notech_or4 i_45871522(.A(n_61890), .B(n_61725), .C(n_61861), .D(n_214984569
		), .Z(n_113483590));
	notech_and4 i_52437(.A(n_344281909), .B(n_341381880), .C(n_344381910), .D
		(n_113483590), .Z(\nbus_11337[0] ));
	notech_nand2 i_51571465(.A(opz[0]), .B(n_113683592), .Z(n_113583591));
	notech_nand2 i_51271468(.A(n_58691), .B(n_57218), .Z(n_113683592));
	notech_nao3 i_51471466(.A(n_345785866), .B(instrc[104]), .C(n_339561023)
		, .Z(n_113883594));
	notech_nao3 i_52371457(.A(n_345785866), .B(instrc[105]), .C(n_339561023)
		, .Z(n_114283598));
	notech_nao3 i_7071894(.A(instrc[115]), .B(instrc[114]), .C(instrc[112]),
		 .Z(n_114683602));
	notech_nao3 i_53271448(.A(instrc[106]), .B(n_345785866), .C(n_339561023)
		, .Z(n_114783603));
	notech_nand2 i_53971441(.A(n_59558), .B(n_32311), .Z(n_114883604));
	notech_or2 i_53871442(.A(n_345585864), .B(n_32260), .Z(n_114983605));
	notech_nor2 i_54271438(.A(n_345585864), .B(n_32274), .Z(n_115083606));
	notech_nor2 i_54471436(.A(n_345585864), .B(n_32276), .Z(n_115183607));
	notech_and2 i_54771433(.A(imm[7]), .B(n_115383609), .Z(n_115283608));
	notech_nand2 i_54671434(.A(n_57057), .B(n_57230), .Z(n_115383609));
	notech_and2 i_55571425(.A(imm[11]), .B(n_32203), .Z(n_115483610));
	notech_and2 i_55771423(.A(imm[12]), .B(n_32203), .Z(n_115583611));
	notech_and2 i_55971421(.A(imm[13]), .B(n_32203), .Z(n_115683612));
	notech_and2 i_56171419(.A(imm[14]), .B(n_32203), .Z(n_115783613));
	notech_nand2 i_106870915(.A(add_src[14]), .B(n_30668), .Z(n_115983615)
		);
	notech_ao4 i_106770916(.A(n_4424), .B(n_349385901), .C(n_4347), .D(n_115783613
		), .Z(n_116883624));
	notech_nao3 i_1512909(.A(n_130783763), .B(n_115983615), .C(n_116883624),
		 .Z(n_21377));
	notech_nand2 i_108770896(.A(add_src[13]), .B(n_30668), .Z(n_116983625)
		);
	notech_ao4 i_108670897(.A(n_4424), .B(n_349385901), .C(n_4347), .D(n_115683612
		), .Z(n_117883634));
	notech_nao3 i_1412908(.A(n_131583771), .B(n_116983625), .C(n_117883634),
		 .Z(n_21372));
	notech_nand2 i_110670877(.A(add_src[12]), .B(n_30668), .Z(n_117983635)
		);
	notech_ao4 i_110570878(.A(n_4424), .B(n_349385901), .C(n_4347), .D(n_115583611
		), .Z(n_118883644));
	notech_nao3 i_1312907(.A(n_132383779), .B(n_117983635), .C(n_118883644),
		 .Z(n_21367));
	notech_nand2 i_112570858(.A(add_src[11]), .B(n_30668), .Z(n_118983645)
		);
	notech_ao4 i_112470859(.A(n_4424), .B(n_349385901), .C(n_4347), .D(n_115483610
		), .Z(n_119883654));
	notech_nao3 i_1212906(.A(n_133183787), .B(n_118983645), .C(n_119883654),
		 .Z(n_21362));
	notech_nand2 i_120170782(.A(add_src[7]), .B(n_30668), .Z(n_119983655));
	notech_ao4 i_120070783(.A(n_4424), .B(n_349385901), .C(n_57024), .D(n_115283608
		), .Z(n_120883664));
	notech_nao3 i_812902(.A(n_133983795), .B(n_119983655), .C(n_120883664), 
		.Z(n_21342));
	notech_nand2 i_122170763(.A(add_src[6]), .B(n_30668), .Z(n_120983665));
	notech_ao4 i_122070764(.A(n_4424), .B(n_349385901), .C(n_348285890), .D(n_115183607
		), .Z(n_121883674));
	notech_nao3 i_712901(.A(n_134783803), .B(n_120983665), .C(n_121883674), 
		.Z(n_21337));
	notech_or4 i_123270752(.A(n_301560644), .B(n_301960648), .C(n_61706), .D
		(opd[4]), .Z(n_121983675));
	notech_nand2 i_123170753(.A(n_344885857), .B(n_121983675), .Z(n_122283678
		));
	notech_ao4 i_123370751(.A(n_31476), .B(n_135683812), .C(n_56983), .D(n_344485853
		), .Z(n_122383679));
	notech_or2 i_124570739(.A(n_347085879), .B(n_31513), .Z(n_123283688));
	notech_or4 i_124970735(.A(n_351885926), .B(n_348485892), .C(opd[4]), .D(opd
		[5]), .Z(n_123383689));
	notech_nand2 i_124770737(.A(opd[5]), .B(n_122283678), .Z(n_123483690));
	notech_ao4 i_124670738(.A(n_115083606), .B(n_348285890), .C(n_4424), .D(n_345385862
		), .Z(n_123583691));
	notech_nor2 i_124870736(.A(n_122383679), .B(n_31477), .Z(n_123683692));
	notech_or4 i_612900(.A(n_123583691), .B(n_123683692), .C(n_136083816), .D
		(n_30446), .Z(n_21332));
	notech_nor2 i_127570709(.A(n_33518), .B(n_345285861), .Z(n_123783693));
	notech_or4 i_127470710(.A(n_32184), .B(n_32628), .C(n_26637), .D(n_61630
		), .Z(n_124983705));
	notech_nao3 i_412898(.A(n_137283828), .B(n_136583821), .C(n_123783693), 
		.Z(n_21322));
	notech_or2 i_130270683(.A(n_350785915101152), .B(n_345285861), .Z(n_125083706
		));
	notech_nand2 i_129070695(.A(n_348485892), .B(n_349485902), .Z(n_125183707
		));
	notech_or4 i_130170684(.A(n_32184), .B(n_32391), .C(n_26637), .D(n_61628
		), .Z(n_126283718));
	notech_nand2 i_130370682(.A(n_125183707), .B(n_58802), .Z(n_126383719)
		);
	notech_nand3 i_312897(.A(n_137983835), .B(n_138383839), .C(n_125083706),
		 .Z(n_21317));
	notech_or2 i_132770658(.A(n_350685914101151), .B(n_345285861), .Z(n_126483720
		));
	notech_or4 i_131670669(.A(n_19707), .B(n_61706), .C(n_31472), .D(opd[1])
		, .Z(n_126583721));
	notech_and4 i_212896(.A(n_138683842), .B(n_138583841), .C(n_139483850), 
		.D(n_126483720), .Z(n_21312));
	notech_nor2 i_134970636(.A(n_350585913101150), .B(n_345285861), .Z(n_127683732
		));
	notech_nor2 i_134870637(.A(n_4352), .B(nbus_11273[0]), .Z(n_128583741)
		);
	notech_or4 i_112895(.A(n_140483860), .B(n_127683732), .C(n_30452), .D(n_30451
		), .Z(n_21307));
	notech_ao4 i_51671464(.A(n_345585864), .B(n_32267), .C(n_58716), .D(n_2845
		), .Z(n_128983745));
	notech_ao4 i_52471456(.A(n_58707), .B(n_2829), .C(n_57104), .D(n_57211),
		 .Z(n_129283748));
	notech_ao4 i_52571455(.A(n_345585864), .B(n_32270), .C(n_31605), .D(n_58691
		), .Z(n_129483750));
	notech_ao4 i_53371447(.A(n_2829), .B(n_2845), .C(n_56898), .D(n_57211), 
		.Z(n_129683752));
	notech_ao4 i_53471446(.A(n_345585864), .B(n_32271), .C(n_31606), .D(n_58691
		), .Z(n_129883754));
	notech_ao4 i_106970914(.A(n_2129), .B(n_32895), .C(n_2128), .D(n_32866),
		 .Z(n_130183757));
	notech_ao4 i_107070913(.A(n_4353), .B(nbus_11271[14]), .C(n_4349), .D(n_33497
		), .Z(n_130283758));
	notech_ao4 i_107170912(.A(n_24142), .B(n_33499), .C(n_4350), .D(n_33498)
		, .Z(n_130483760));
	notech_ao4 i_107270911(.A(n_2127), .B(n_31522), .C(n_4352), .D(nbus_11273
		[14]), .Z(n_130583761));
	notech_and4 i_107570908(.A(n_130583761), .B(n_130483760), .C(n_130283758
		), .D(n_130183757), .Z(n_130783763));
	notech_ao4 i_108870895(.A(n_2129), .B(n_32894), .C(n_2128), .D(n_32865),
		 .Z(n_130983765));
	notech_ao4 i_108970894(.A(n_4350), .B(n_33501), .C(n_4349), .D(n_33500),
		 .Z(n_131083766));
	notech_ao4 i_109070893(.A(n_4353), .B(nbus_11271[13]), .C(n_24142), .D(n_33502
		), .Z(n_131283768));
	notech_ao4 i_109170892(.A(n_2127), .B(n_31521), .C(n_4352), .D(nbus_11273
		[13]), .Z(n_131383769));
	notech_and4 i_109470889(.A(n_131383769), .B(n_131283768), .C(n_131083766
		), .D(n_130983765), .Z(n_131583771));
	notech_ao4 i_110770876(.A(n_2129), .B(n_32893), .C(n_2128), .D(n_32864),
		 .Z(n_131783773));
	notech_ao4 i_110870875(.A(n_4350), .B(n_33504), .C(n_4349), .D(n_33503),
		 .Z(n_131883774));
	notech_ao4 i_110970874(.A(n_4353), .B(nbus_11271[12]), .C(n_24142), .D(n_33505
		), .Z(n_132083776));
	notech_ao4 i_111070873(.A(n_2127), .B(n_31520), .C(n_4352), .D(n_58321),
		 .Z(n_132183777));
	notech_and4 i_111370870(.A(n_132183777), .B(n_132083776), .C(n_131883774
		), .D(n_131783773), .Z(n_132383779));
	notech_ao4 i_112670857(.A(n_2129), .B(n_32892), .C(n_2128), .D(n_32863),
		 .Z(n_132583781));
	notech_ao4 i_112770856(.A(n_4353), .B(nbus_11271[11]), .C(n_4349), .D(n_33506
		), .Z(n_132683782));
	notech_ao4 i_112870855(.A(n_24142), .B(n_33508), .C(n_4350), .D(n_33507)
		, .Z(n_132883784));
	notech_ao4 i_112970854(.A(n_2127), .B(n_31519), .C(n_4352), .D(n_58312),
		 .Z(n_132983785));
	notech_and4 i_113270851(.A(n_132983785), .B(n_132883784), .C(n_132683782
		), .D(n_132583781), .Z(n_133183787));
	notech_ao4 i_120270781(.A(n_2129), .B(n_32888), .C(n_2128), .D(n_32859),
		 .Z(n_133383789));
	notech_ao4 i_120370780(.A(n_4353), .B(nbus_11271[7]), .C(n_4349), .D(n_33509
		), .Z(n_133483790));
	notech_ao4 i_120470779(.A(n_24142), .B(n_33511), .C(n_4350), .D(n_33510)
		, .Z(n_133683792));
	notech_ao4 i_120570778(.A(n_2127), .B(n_31515), .C(n_4352), .D(nbus_11273
		[7]), .Z(n_133783793));
	notech_and4 i_120870775(.A(n_133783793), .B(n_133683792), .C(n_133483790
		), .D(n_133383789), .Z(n_133983795));
	notech_ao4 i_122270762(.A(n_2129), .B(n_32887), .C(n_2128), .D(n_32858),
		 .Z(n_134183797));
	notech_ao4 i_122370761(.A(n_4353), .B(nbus_11271[6]), .C(n_4349), .D(n_33512
		), .Z(n_134283798));
	notech_ao4 i_122470760(.A(n_24142), .B(n_33514), .C(n_4350), .D(n_33513)
		, .Z(n_134483800));
	notech_ao4 i_122570759(.A(n_2127), .B(n_31514), .C(n_4352), .D(nbus_11273
		[6]), .Z(n_134583801));
	notech_and4 i_122870756(.A(n_134583801), .B(n_134483800), .C(n_134283798
		), .D(n_134183797), .Z(n_134783803));
	notech_ao4 i_125170733(.A(n_2128), .B(n_32857), .C(n_344785856), .D(n_32322
		), .Z(n_134983805));
	notech_ao4 i_125270732(.A(n_4349), .B(n_33515), .C(n_2129), .D(n_32886),
		 .Z(n_135183807));
	notech_ao4 i_125370731(.A(n_33516), .B(n_4350), .C(n_4353), .D(nbus_11271
		[5]), .Z(n_135283808));
	notech_and4 i_125870726(.A(n_135283808), .B(n_135183807), .C(n_134983805
		), .D(n_123283688), .Z(n_135483810));
	notech_or2 i_123670748(.A(n_347185880), .B(opd[5]), .Z(n_135683812));
	notech_ao4 i_125470730(.A(n_4352), .B(nbus_11273[5]), .C(n_24142), .D(n_33517
		), .Z(n_135883814));
	notech_nand3 i_125970725(.A(n_135883814), .B(n_123383689), .C(n_123483690
		), .Z(n_136083816));
	notech_ao4 i_128270703(.A(n_347085879), .B(n_31511), .C(n_4352), .D(nbus_11273
		[3]), .Z(n_136283818));
	notech_ao4 i_127670708(.A(n_351885926), .B(n_348485892), .C(n_344785856)
		, .D(n_32320), .Z(n_136383819));
	notech_and3 i_128670699(.A(n_124983705), .B(n_136383819), .C(n_136283818
		), .Z(n_136583821));
	notech_ao4 i_127770707(.A(n_2128), .B(n_32856), .C(n_347185880), .D(opd[
		3]), .Z(n_136683822));
	notech_ao4 i_127970706(.A(n_4349), .B(n_33519), .C(n_2129), .D(n_32884),
		 .Z(n_136783823));
	notech_ao4 i_128070705(.A(n_4350), .B(n_33520), .C(n_4353), .D(nbus_11271
		[3]), .Z(n_136983825));
	notech_ao4 i_128170704(.A(n_31476), .B(n_349085898), .C(n_24142), .D(n_33521
		), .Z(n_137083826));
	notech_and4 i_128770698(.A(n_137083826), .B(n_136983825), .C(n_136783823
		), .D(n_136683822), .Z(n_137283828));
	notech_ao4 i_130470681(.A(n_344785856), .B(n_32318), .C(n_58802), .D(n_348885896
		), .Z(n_137483830));
	notech_ao4 i_130570680(.A(n_2129), .B(n_32883), .C(n_2128), .D(n_32855),
		 .Z(n_137683832));
	notech_ao4 i_130670679(.A(n_4353), .B(nbus_11271[2]), .C(n_4349), .D(n_33523
		), .Z(n_137783833));
	notech_and4 i_131270673(.A(n_137783833), .B(n_137683832), .C(n_137483830
		), .D(n_126283718), .Z(n_137983835));
	notech_ao4 i_130770678(.A(n_24142), .B(n_33525), .C(n_4350), .D(n_33524)
		, .Z(n_138083836));
	notech_ao4 i_130870677(.A(n_31510), .B(n_347085879), .C(n_4352), .D(nbus_11273
		[2]), .Z(n_138183837));
	notech_and3 i_131370672(.A(n_138183837), .B(n_138083836), .C(n_126383719
		), .Z(n_138383839));
	notech_ao4 i_133270653(.A(n_24142), .B(n_33529), .C(n_4350), .D(n_33528)
		, .Z(n_138583841));
	notech_ao4 i_133370652(.A(n_347085879), .B(n_31509), .C(n_4352), .D(n_58225
		), .Z(n_138683842));
	notech_and2 i_132870657(.A(n_348485892), .B(n_126583721), .Z(n_138883844
		));
	notech_ao4 i_132970656(.A(n_344785856), .B(n_32316), .C(n_31473), .D(n_348685894
		), .Z(n_138983845));
	notech_ao4 i_133070655(.A(n_2129), .B(n_32882), .C(n_2128), .D(n_32854),
		 .Z(n_139183847));
	notech_ao4 i_133170654(.A(n_4353), .B(nbus_11271[1]), .C(n_4349), .D(n_33527
		), .Z(n_139283848));
	notech_and4 i_133770648(.A(n_139283848), .B(n_139183847), .C(n_138983845
		), .D(n_138883844), .Z(n_139483850));
	notech_ao4 i_135370632(.A(n_4350), .B(n_33532), .C(n_4353), .D(nbus_11271
		[0]), .Z(n_139683852));
	notech_ao4 i_135470631(.A(n_347085879), .B(n_31508), .C(n_24142), .D(n_33533
		), .Z(n_139783853));
	notech_ao4 i_135170634(.A(n_2128), .B(n_32853), .C(n_344785856), .D(n_32313
		), .Z(n_140183857));
	notech_ao4 i_135270633(.A(n_4349), .B(n_33531), .C(n_2129), .D(n_32881),
		 .Z(n_140283858));
	notech_nand2 i_135670629(.A(n_140283858), .B(n_140183857), .Z(n_140383859
		));
	notech_or4 i_135870627(.A(n_348385891), .B(n_128583741), .C(n_344385852)
		, .D(n_140383859), .Z(n_140483860));
	notech_mux2 i_6266094(.S(n_32273), .A(n_141283868), .B(n_141083866), .Z(n_140683862
		));
	notech_and2 i_6366093(.A(n_28240), .B(n_390864439), .Z(n_140783863));
	notech_and3 i_6466092(.A(n_331360941), .B(n_331260940), .C(n_390964440),
		 .Z(n_140883864));
	notech_ao4 i_4366113(.A(n_60177), .B(\nbus_11290[1] ), .C(n_30920), .D(n_30788
		), .Z(n_141083866));
	notech_ao4 i_4266114(.A(n_60177), .B(n_58225), .C(n_30919), .D(n_30788),
		 .Z(n_141283868));
	notech_and3 i_6066096(.A(n_382164352), .B(n_329260920), .C(n_330260930),
		 .Z(n_141583871));
	notech_and4 i_6166095(.A(n_381964350), .B(n_331260940), .C(n_329460922),
		 .D(n_330160929), .Z(n_141683872));
	notech_mux2 i_5466102(.S(n_32544), .A(n_141983875), .B(n_142183877), .Z(n_141783873
		));
	notech_ao4 i_3966117(.A(n_60177), .B(n_58225), .C(n_30919), .D(n_28555),
		 .Z(n_141983875));
	notech_ao4 i_3866118(.A(n_60170), .B(n_59001), .C(n_30920), .D(n_28555),
		 .Z(n_142183877));
	notech_nand3 i_59065578(.A(n_61091), .B(n_61628), .C(read_data[1]), .Z(n_142483880
		));
	notech_ao4 i_5266104(.A(n_32697), .B(n_31362), .C(n_163396015), .D(n_30906
		), .Z(n_142583881));
	notech_and2 i_5366103(.A(n_332960957), .B(n_329660924), .Z(n_142683882)
		);
	notech_ao4 i_4866108(.A(n_32697), .B(n_30731), .C(n_29419), .D(n_30283),
		 .Z(n_142783883));
	notech_and3 i_4966107(.A(n_442368007), .B(n_29533), .C(n_29540), .Z(n_142883884
		));
	notech_nand2 i_7566081(.A(tsc[24]), .B(n_30615), .Z(n_142983885));
	notech_or2 i_7466082(.A(n_131426641), .B(n_60519), .Z(n_143283888));
	notech_or2 i_6966087(.A(n_387964410), .B(n_58893), .Z(n_143783893));
	notech_or2 i_26965888(.A(n_55955), .B(n_30995), .Z(n_145683912));
	notech_nao3 i_26665891(.A(n_19612), .B(read_data[14]), .C(n_35412112), .Z
		(n_145983915));
	notech_or4 i_26365894(.A(n_56003), .B(n_378564316), .C(n_61938), .D(nbus_11271
		[14]), .Z(n_146283918));
	notech_nand3 i_74965419(.A(n_1640), .B(n_171160315), .C(n_1736), .Z(n_148583941
		));
	notech_or2 i_74665422(.A(n_444668030), .B(n_97342414), .Z(n_148883944)
		);
	notech_nand2 i_74365425(.A(sav_edi[14]), .B(n_61861), .Z(n_149183947));
	notech_or2 i_77765391(.A(n_337361001), .B(nbus_11271[30]), .Z(n_149483950
		));
	notech_or2 i_77465394(.A(n_122826555), .B(n_33194), .Z(n_149783953));
	notech_nand3 i_77165397(.A(n_55904), .B(n_171160315), .C(n_1767), .Z(n_150083956
		));
	notech_or2 i_76865400(.A(n_5750), .B(n_122226549), .Z(n_150383959));
	notech_and4 i_97865190(.A(n_29557), .B(n_30282), .C(n_63758), .D(opc_10[
		14]), .Z(n_150483960));
	notech_or2 i_97365195(.A(n_445268036), .B(n_31487), .Z(n_151183967));
	notech_or2 i_99665172(.A(n_443168015), .B(n_60519), .Z(n_151283968));
	notech_or2 i_99165177(.A(n_443368017), .B(n_58893), .Z(n_151983975));
	notech_ao4 i_186564328(.A(n_118426511), .B(n_33171), .C(n_118526512), .D
		(n_106826395), .Z(n_152083976));
	notech_ao4 i_186464329(.A(n_443468018), .B(n_364628688), .C(n_443268016)
		, .D(n_58429), .Z(n_152283978));
	notech_and3 i_186764326(.A(n_152083976), .B(n_152283978), .C(n_151983975
		), .Z(n_152383979));
	notech_ao4 i_186264331(.A(n_443568019), .B(n_31942), .C(n_305744491), .D
		(n_31500), .Z(n_152483980));
	notech_ao4 i_184964344(.A(\nbus_11290[14] ), .B(n_142883884), .C(nbus_11273
		[14]), .D(n_30455), .Z(n_152783983));
	notech_ao4 i_184864345(.A(n_57612), .B(n_33215), .C(n_57057), .D(n_377064301
		), .Z(n_152983985));
	notech_nand3 i_185164342(.A(n_152783983), .B(n_152983985), .C(n_151183967
		), .Z(n_153083986));
	notech_ao4 i_184664347(.A(n_29418), .B(n_377164302), .C(n_57611), .D(n_97342414
		), .Z(n_153183987));
	notech_ao4 i_165864534(.A(n_57001), .B(n_31538), .C(n_61091), .D(n_30859
		), .Z(n_153483990));
	notech_ao4 i_165664536(.A(n_55884), .B(n_33539), .C(n_331060938), .D(n_31506
		), .Z(n_153683992));
	notech_and4 i_166064532(.A(n_153683992), .B(n_153483990), .C(n_150083956
		), .D(n_150383959), .Z(n_153883994));
	notech_ao4 i_165364539(.A(n_122726554), .B(\nbus_11283[30] ), .C(n_122626553
		), .D(\nbus_11290[30] ), .Z(n_153983995));
	notech_ao4 i_165164541(.A(n_337461002), .B(n_318771158), .C(n_5758), .D(n_122926556
		), .Z(n_154183997));
	notech_and4 i_165564537(.A(n_154183997), .B(n_153983995), .C(n_149483950
		), .D(n_149783953), .Z(n_154383999));
	notech_ao4 i_163664556(.A(\nbus_11290[14] ), .B(n_142683882), .C(nbus_11273
		[14]), .D(n_30454), .Z(n_154484000));
	notech_ao4 i_163464558(.A(n_444568029), .B(n_33215), .C(n_444868032), .D
		(n_31487), .Z(n_154684002));
	notech_and4 i_163864554(.A(n_154684002), .B(n_154484000), .C(n_148883944
		), .D(n_149183947), .Z(n_154884004));
	notech_ao4 i_163164561(.A(n_28365), .B(n_377264303), .C(n_28367), .D(n_377164302
		), .Z(n_154984005));
	notech_ao4 i_162964563(.A(n_331760945), .B(n_385364384), .C(n_333260960)
		, .D(n_33538), .Z(n_155184007));
	notech_and3 i_163064562(.A(n_169684152), .B(n_155184007), .C(n_160684062
		), .Z(n_155284008));
	notech_ao4 i_149464696(.A(n_28260), .B(n_30896), .C(n_28558), .D(n_141783873
		), .Z(n_155484010));
	notech_ao4 i_149364697(.A(n_59001), .B(n_436967953), .C(n_58225), .D(n_437067954
		), .Z(n_155584011));
	notech_ao4 i_149164699(.A(n_55884), .B(n_33537), .C(n_61091), .D(n_30833
		), .Z(n_155784013));
	notech_ao4 i_149064700(.A(n_439467978), .B(n_56956), .C(n_333260960), .D
		(n_33536), .Z(n_155884014));
	notech_and4 i_149664694(.A(n_155884014), .B(n_155784013), .C(n_155584011
		), .D(n_155484010), .Z(n_156084016));
	notech_ao4 i_148764703(.A(n_30891), .B(n_439367977), .C(n_331660944), .D
		(n_334060968), .Z(n_156184017));
	notech_ao4 i_148664704(.A(n_439667980), .B(n_334360971), .C(n_439567979)
		, .D(n_33103), .Z(n_156284018));
	notech_ao4 i_148464706(.A(n_28252), .B(n_30916), .C(n_28251), .D(n_30914
		), .Z(n_156584021));
	notech_and3 i_148564705(.A(n_169484150), .B(n_142483880), .C(n_156584021
		), .Z(n_156684022));
	notech_ao4 i_122064963(.A(n_141683872), .B(n_59041), .C(n_58339), .D(n_141583871
		), .Z(n_157084026));
	notech_ao4 i_121964964(.A(n_378464315), .B(n_31487), .C(n_61087), .D(n_30793
		), .Z(n_157184027));
	notech_ao4 i_121764966(.A(n_97342414), .B(n_378864319), .C(n_378964320),
		 .D(n_33215), .Z(n_157384029));
	notech_and4 i_122264961(.A(n_146283918), .B(n_157384029), .C(n_157184027
		), .D(n_157084026), .Z(n_157584031));
	notech_ao4 i_121464969(.A(n_385364384), .B(n_331560943), .C(n_377264303)
		, .D(n_26396), .Z(n_157684032));
	notech_ao4 i_121064971(.A(n_55975), .B(n_32073), .C(n_55966), .D(n_33535
		), .Z(n_157884034));
	notech_and4 i_121664967(.A(n_157884034), .B(n_157684032), .C(n_145683912
		), .D(n_145983915), .Z(n_158084036));
	notech_ao4 i_107565094(.A(n_58225), .B(n_140783863), .C(n_338061008), .D
		(n_140683862), .Z(n_158184037));
	notech_ao4 i_107465095(.A(n_61087), .B(n_30777), .C(n_140883864), .D(n_59001
		), .Z(n_158284038));
	notech_ao4 i_107265097(.A(n_331460942), .B(n_56956), .C(n_55946), .D(n_31509
		), .Z(n_158484040));
	notech_ao4 i_107165098(.A(n_30891), .B(n_332160949), .C(n_334060968), .D
		(n_26603), .Z(n_158584041));
	notech_and4 i_107765092(.A(n_158584041), .B(n_158484040), .C(n_158284038
		), .D(n_158184037), .Z(n_158784043));
	notech_ao4 i_106865101(.A(n_334360971), .B(n_332460952), .C(n_332260950)
		, .D(n_33103), .Z(n_158884044));
	notech_ao4 i_106765102(.A(n_30914), .B(n_26268), .C(n_30896), .D(n_26278
		), .Z(n_158984045));
	notech_ao4 i_106465104(.A(n_55966), .B(n_33534), .C(n_30916), .D(n_26271
		), .Z(n_159184047));
	notech_ao4 i_106365105(.A(n_55955), .B(n_30969), .C(n_55975), .D(n_32060
		), .Z(n_159284048));
	notech_and4 i_107065099(.A(n_159284048), .B(n_159184047), .C(n_158984045
		), .D(n_158884044), .Z(n_159484050));
	notech_ao4 i_103565133(.A(n_131526642), .B(n_33171), .C(n_106826395), .D
		(n_131626643), .Z(n_159584051));
	notech_ao4 i_103465134(.A(n_388064411), .B(n_364628688), .C(n_387864409)
		, .D(n_58429), .Z(n_159784053));
	notech_ao4 i_103165137(.A(n_31942), .B(n_388164412), .C(n_31500), .D(n_390064431
		), .Z(n_159984055));
	notech_and4 i_103365135(.A(n_443068014), .B(n_159984055), .C(n_143283888
		), .D(n_142983885), .Z(n_160284058));
	notech_nand3 i_12263237(.A(n_61091), .B(n_61628), .C(read_data[14]), .Z(n_160684062
		));
	notech_nor2 i_14363216(.A(n_177284202), .B(n_333060958), .Z(n_160884064)
		);
	notech_and3 i_14463215(.A(n_332960957), .B(n_163784093), .C(n_332860956)
		, .Z(n_160984065));
	notech_mux2 i_14063219(.S(n_32244), .A(n_161484070), .B(n_161284068), .Z
		(n_161084066));
	notech_ao4 i_10363254(.A(n_60163), .B(n_59005), .C(n_29557), .D(n_30920)
		, .Z(n_161284068));
	notech_ao4 i_10263255(.A(n_60169), .B(n_58225), .C(n_30919), .D(n_29557)
		, .Z(n_161484070));
	notech_nand2 i_23963120(.A(tsc[30]), .B(n_30615), .Z(n_161784073));
	notech_nao3 i_23863121(.A(opc_10[30]), .B(n_63758), .C(n_388164412), .Z(n_162084076
		));
	notech_or2 i_23363126(.A(n_387964410), .B(\nbus_11290[30] ), .Z(n_162584081
		));
	notech_or2 i_65562728(.A(n_336760995), .B(n_331660944), .Z(n_163084086)
		);
	notech_or4 i_65262731(.A(n_28551), .B(n_61938), .C(n_31611), .D(n_30441)
		, .Z(n_163384089));
	notech_nand3 i_64962734(.A(n_171160315), .B(n_1708), .C(n_1640), .Z(n_163684092
		));
	notech_or4 i_65962724(.A(n_2382), .B(n_2383), .C(n_165695997), .D(n_28552
		), .Z(n_163784093));
	notech_ao3 i_71162672(.A(opc_10[30]), .B(n_63780), .C(n_28869), .Z(n_163984095
		));
	notech_or2 i_70662677(.A(n_28863), .B(\nbus_11290[30] ), .Z(n_164684102)
		);
	notech_or2 i_75762626(.A(n_386464395), .B(n_56956), .Z(n_165184107));
	notech_or2 i_75462629(.A(n_29540), .B(n_334360971), .Z(n_165484110));
	notech_or2 i_75162632(.A(n_30280), .B(n_57057), .Z(n_165784113));
	notech_or2 i_77962604(.A(n_57362), .B(n_58992), .Z(n_166584121));
	notech_ao3 i_84762542(.A(opc_10[30]), .B(n_63782), .C(n_444068024), .Z(n_166684122
		));
	notech_or2 i_84262547(.A(n_443868022), .B(n_58992), .Z(n_167384129));
	notech_ao3 i_88462507(.A(opc_10[30]), .B(n_63780), .C(n_443568019), .Z(n_167484130
		));
	notech_or2 i_87962512(.A(n_443368017), .B(n_58992), .Z(n_168184137));
	notech_ao3 i_92062472(.A(opc_10[30]), .B(n_63780), .C(n_442768011), .Z(n_168284138
		));
	notech_or2 i_91462477(.A(n_442568009), .B(n_58992), .Z(n_168984145));
	notech_nor2 i_92362469(.A(n_30693), .B(n_58992), .Z(n_169384149));
	notech_ao4 i_31256(.A(n_331360941), .B(n_59005), .C(n_28240), .D(n_58225
		), .Z(n_169484150));
	notech_ao4 i_8563272(.A(n_59041), .B(n_381964350), .C(n_58339), .D(n_382164352
		), .Z(n_169684152));
	notech_ao4 i_167561740(.A(n_117626503), .B(n_33194), .C(n_117726504), .D
		(n_5758), .Z(n_169784153));
	notech_ao4 i_167461741(.A(n_442968013), .B(n_5750), .C(n_442668010), .D(\nbus_11283[30] 
		), .Z(n_169984155));
	notech_nand3 i_167761738(.A(n_169784153), .B(n_169984155), .C(n_168984145
		), .Z(n_170084156));
	notech_ao4 i_167261743(.A(n_442868012), .B(nbus_11271[30]), .C(n_327960907
		), .D(n_31506), .Z(n_170184157));
	notech_ao4 i_167961736(.A(n_30697), .B(n_33194), .C(n_30689), .D(n_5758)
		, .Z(n_170284158));
	notech_ao4 i_167861737(.A(n_61702), .B(n_31538), .C(n_30695), .D(\nbus_11283[30] 
		), .Z(n_170484160));
	notech_nao3 i_52263349(.A(n_170284158), .B(n_170484160), .C(n_169384149)
		, .Z(n_170584161));
	notech_ao4 i_164861767(.A(n_118426511), .B(n_33194), .C(n_118526512), .D
		(n_5758), .Z(n_171284164));
	notech_ao4 i_164761768(.A(n_5750), .B(n_443468018), .C(\nbus_11283[30] )
		, .D(n_443268016), .Z(n_171484166));
	notech_nand3 i_165061765(.A(n_171284164), .B(n_171484166), .C(n_168184137
		), .Z(n_171584167));
	notech_ao4 i_164561770(.A(nbus_11271[30]), .B(n_443168015), .C(n_305744491
		), .D(n_31506), .Z(n_171684168));
	notech_ao4 i_162061795(.A(n_119226519), .B(n_33194), .C(n_119326520), .D
		(n_5758), .Z(n_171984171));
	notech_ao4 i_161961796(.A(n_443968023), .B(n_5750), .C(n_443768021), .D(n_58483
		), .Z(n_172184173));
	notech_nand3 i_162261793(.A(n_171984171), .B(n_172184173), .C(n_167384129
		), .Z(n_172284174));
	notech_ao4 i_161761798(.A(n_443668020), .B(nbus_11271[30]), .C(n_379264323
		), .D(n_31506), .Z(n_172584175));
	notech_ao4 i_153761877(.A(n_57319), .B(n_33194), .C(n_57320), .D(n_5758)
		, .Z(n_172884178));
	notech_ao4 i_153661878(.A(n_303822063), .B(n_5750), .C(n_57363), .D(n_58483
		), .Z(n_173084180));
	notech_and3 i_153961875(.A(n_172884178), .B(n_173084180), .C(n_166584121
		), .Z(n_173184181));
	notech_ao4 i_153361880(.A(n_303922064), .B(nbus_11271[30]), .C(n_386864399
		), .D(n_31506), .Z(n_173284182));
	notech_ao4 i_153261881(.A(n_61702), .B(n_31538), .C(n_299122016), .D(n_318771158
		), .Z(n_173384183));
	notech_ao4 i_151761896(.A(n_29342), .B(n_30896), .C(n_29560), .D(n_161084066
		), .Z(n_173784185));
	notech_ao4 i_151561898(.A(n_194884375), .B(n_59001), .C(n_58225), .D(n_439767981
		), .Z(n_174784187));
	notech_and4 i_151961894(.A(n_174784187), .B(n_173784185), .C(n_165484110
		), .D(n_165784113), .Z(n_174984189));
	notech_ao4 i_151261901(.A(n_29333), .B(n_30914), .C(n_29550), .D(n_33103
		), .Z(n_175084190));
	notech_ao4 i_151061903(.A(n_378364314), .B(n_30891), .C(n_29334), .D(n_30916
		), .Z(n_175284192));
	notech_and4 i_151461899(.A(n_30274), .B(n_175284192), .C(n_175084190), .D
		(n_165184107), .Z(n_175484194));
	notech_ao4 i_147761936(.A(n_388364414), .B(n_33194), .C(n_388264413), .D
		(n_5758), .Z(n_175584195));
	notech_ao4 i_147661937(.A(n_28852), .B(n_5750), .C(n_28874), .D(n_58483)
		, .Z(n_175784197));
	notech_nand3 i_147961934(.A(n_175584195), .B(n_175784197), .C(n_164684102
		), .Z(n_175884198));
	notech_ao4 i_147461939(.A(n_28867), .B(n_60611), .C(n_28854), .D(n_31506
		), .Z(n_176584199));
	notech_ao4 i_139762015(.A(n_32697), .B(n_31362), .C(n_30906), .D(n_30633
		), .Z(n_177284202));
	notech_ao4 i_139362019(.A(\nbus_11290[0] ), .B(n_160984065), .C(n_58238)
		, .D(n_160884064), .Z(n_177484204));
	notech_ao4 i_139162021(.A(n_327660904), .B(n_28251), .C(n_333260960), .D
		(n_33540), .Z(n_177684206));
	notech_and4 i_139562017(.A(n_163384089), .B(n_177684206), .C(n_177484204
		), .D(n_163684092), .Z(n_177884208));
	notech_ao4 i_138862024(.A(n_439567979), .B(n_33169), .C(n_101142452), .D
		(n_439667980), .Z(n_177984209));
	notech_ao4 i_138662026(.A(n_61091), .B(n_30832), .C(n_439467978), .D(n_31472
		), .Z(n_178184211));
	notech_and3 i_138762025(.A(n_169576761), .B(n_178184211), .C(n_116976235
		), .Z(n_178284212));
	notech_ao4 i_102462372(.A(n_131526642), .B(n_33194), .C(n_5758), .D(n_131626643
		), .Z(n_178484214));
	notech_ao4 i_102362373(.A(n_5750), .B(n_388064411), .C(n_58483), .D(n_387864409
		), .Z(n_178684216));
	notech_ao4 i_102062376(.A(n_60611), .B(n_131426641), .C(n_390064431), .D
		(n_31506), .Z(n_178884218));
	notech_and4 i_102262374(.A(n_178884218), .B(n_162084076), .C(n_30502), .D
		(n_161784073), .Z(n_179184221));
	notech_or2 i_173060647(.A(n_57383), .B(n_58601), .Z(n_179284222));
	notech_or4 i_173160646(.A(instrc[123]), .B(n_318060808), .C(n_57383), .D
		(instrc[120]), .Z(n_179384223));
	notech_nao3 i_173360645(.A(n_30553), .B(n_58592), .C(n_57383), .Z(n_179484224
		));
	notech_or4 i_173460644(.A(instrc[123]), .B(n_318060808), .C(n_188084307)
		, .D(instrc[120]), .Z(n_179584225));
	notech_and3 i_5760583(.A(n_385664387), .B(n_256963516), .C(n_30640), .Z(n_179684226
		));
	notech_and4 i_5860582(.A(n_385864389), .B(n_2570), .C(n_383464365), .D(n_58664
		), .Z(n_179784227));
	notech_and2 i_5560585(.A(n_192684353), .B(n_180084230), .Z(n_179884228)
		);
	notech_mux2 i_5660584(.S(n_58601), .A(n_30919), .B(n_30920), .Z(n_179984229
		));
	notech_nao3 i_24860397(.A(opa[1]), .B(n_58592), .C(n_60163), .Z(n_180084230
		));
	notech_ao3 i_5360587(.A(n_382864359), .B(n_256963516), .C(n_383364364), 
		.Z(n_180584233));
	notech_and4 i_5460586(.A(n_58664), .B(n_382664357), .C(n_383464365), .D(n_185684283
		), .Z(n_180684234));
	notech_nand2 i_77759928(.A(n_382064351), .B(n_25121), .Z(n_180784235));
	notech_nand2 i_79459911(.A(n_115942600), .B(n_32219), .Z(n_180884236));
	notech_or4 i_23160412(.A(instrc[115]), .B(instrc[112]), .C(n_58716), .D(n_327560903
		), .Z(n_181184239));
	notech_or2 i_22860415(.A(n_101142452), .B(n_382664357), .Z(n_181484242)
		);
	notech_nand2 i_22560418(.A(tsc[32]), .B(n_30615), .Z(n_181784245));
	notech_or4 i_24260402(.A(n_63716), .B(n_188084307), .C(n_61938), .D(n_58225
		), .Z(n_182284250));
	notech_or2 i_23860405(.A(n_334360971), .B(n_382664357), .Z(n_182584253)
		);
	notech_nand2 i_41260261(.A(n_30354), .B(opd[14]), .Z(n_184784274));
	notech_nao3 i_41160262(.A(n_63794), .B(opc[14]), .C(n_441868002), .Z(n_185084277
		));
	notech_or4 i_40560267(.A(n_58592), .B(n_384764378), .C(n_384964380), .D(n_97342414
		), .Z(n_185584282));
	notech_or4 i_41460259(.A(n_32269), .B(n_384764378), .C(instrc[120]), .D(n_384864379
		), .Z(n_185684283));
	notech_nand2 i_206763373(.A(n_61630), .B(read_data[30]), .Z(n_185884285)
		);
	notech_or2 i_43760239(.A(n_25110), .B(n_60611), .Z(n_186184288));
	notech_nao3 i_43360242(.A(opc_10[30]), .B(n_63758), .C(n_365428694), .Z(n_186484291
		));
	notech_or4 i_43060245(.A(n_58716), .B(n_58707), .C(n_57256), .D(n_5750),
		 .Z(n_186784294));
	notech_or4 i_49960198(.A(n_57438), .B(n_26063), .C(n_58550), .D(n_31074)
		, .Z(n_187284299));
	notech_or2 i_49360201(.A(n_5783), .B(n_31477), .Z(n_187584302));
	notech_or2 i_108060766(.A(n_57383), .B(n_25121), .Z(n_188084307));
	notech_ao4 i_125459479(.A(n_150969547), .B(n_31068), .C(n_151069548), .D
		(n_31067), .Z(n_188184308));
	notech_ao4 i_125159480(.A(n_57027), .B(n_33104), .C(n_57068), .D(n_187176929
		), .Z(n_188284309));
	notech_ao4 i_124959482(.A(n_57438), .B(n_31047), .C(n_57036), .D(n_334660974
		), .Z(n_188484311));
	notech_and4 i_125659477(.A(n_188484311), .B(n_188284309), .C(n_188184308
		), .D(n_187584302), .Z(n_188684313));
	notech_ao4 i_124459485(.A(n_143469472), .B(n_31071), .C(n_143769475), .D
		(n_31048), .Z(n_188784314));
	notech_ao4 i_124259487(.A(n_143569473), .B(n_31075), .C(n_143369471), .D
		(n_31072), .Z(n_188984316));
	notech_and4 i_124859483(.A(n_187576933), .B(n_188984316), .C(n_188784314
		), .D(n_187284299), .Z(n_189184318));
	notech_ao4 i_116559556(.A(n_365628696), .B(n_58483), .C(n_56030), .D(n_32581
		), .Z(n_189284319));
	notech_ao4 i_116359558(.A(n_365528695), .B(n_58992), .C(n_382264353), .D
		(n_31506), .Z(n_189484321));
	notech_and4 i_116759554(.A(n_189484321), .B(n_189284319), .C(n_186484291
		), .D(n_186784294), .Z(n_189684323));
	notech_ao4 i_116059561(.A(n_365228692), .B(n_33194), .C(n_5758), .D(n_365328693
		), .Z(n_189784324));
	notech_and4 i_116259559(.A(n_55802), .B(n_186184288), .C(n_189784324), .D
		(n_185884285), .Z(n_190084327));
	notech_ao4 i_114259579(.A(n_180684234), .B(n_59041), .C(n_58339), .D(n_180584233
		), .Z(n_190484331));
	notech_ao4 i_114159580(.A(n_385464385), .B(n_377264303), .C(n_385664387)
		, .D(n_33215), .Z(n_190684333));
	notech_ao4 i_113859583(.A(n_56030), .B(n_32566), .C(n_57178), .D(n_377064301
		), .Z(n_190884335));
	notech_and4 i_114059581(.A(n_190884335), .B(n_186576923), .C(n_184784274
		), .D(n_185084277), .Z(n_191184338));
	notech_ao4 i_102459682(.A(n_31075), .B(n_179484224), .C(n_31074), .D(n_179584225
		), .Z(n_191284339));
	notech_ao4 i_102359683(.A(n_31071), .B(n_179284222), .C(n_179384223), .D
		(n_31072), .Z(n_191384340));
	notech_ao4 i_102159685(.A(n_56030), .B(n_32556), .C(n_187176929), .D(n_57174
		), .Z(n_191584342));
	notech_ao4 i_102059686(.A(n_382864359), .B(n_33104), .C(n_31068), .D(n_383064361
		), .Z(n_191684343));
	notech_and4 i_102659680(.A(n_191684343), .B(n_191584342), .C(n_191384340
		), .D(n_191284339), .Z(n_191884345));
	notech_ao4 i_101759689(.A(n_31067), .B(n_57260), .C(n_334660974), .D(n_382664357
		), .Z(n_191984346));
	notech_ao4 i_101659690(.A(n_31048), .B(n_188084307), .C(n_31047), .D(n_57383
		), .Z(n_192084347));
	notech_ao4 i_101459692(.A(n_58664), .B(\nbus_11290[4] ), .C(n_58051), .D
		(n_31477), .Z(n_192284349));
	notech_ao3 i_101559691(.A(n_187576933), .B(n_192284349), .C(n_335060978)
		, .Z(n_192484351));
	notech_ao4 i_99959707(.A(n_58592), .B(n_334260970), .C(n_179984229), .D(n_25121
		), .Z(n_192684353));
	notech_ao4 i_99659710(.A(n_441567999), .B(n_59001), .C(n_384964380), .D(n_179884228
		), .Z(n_192784354));
	notech_ao4 i_99559711(.A(n_56030), .B(n_32553), .C(n_58225), .D(n_440567989
		), .Z(n_192884355));
	notech_ao4 i_99359713(.A(n_382864359), .B(n_33103), .C(n_30916), .D(n_383064361
		), .Z(n_193084357));
	notech_and4 i_99859708(.A(n_193084357), .B(n_192884355), .C(n_192784354)
		, .D(n_182584253), .Z(n_193284359));
	notech_ao4 i_99059716(.A(n_30891), .B(n_57383), .C(n_30914), .D(n_57260)
		, .Z(n_193384360));
	notech_ao4 i_98859718(.A(n_57174), .B(n_30280), .C(n_56956), .D(n_58051)
		, .Z(n_193584362));
	notech_and4 i_99259714(.A(n_193584362), .B(n_193384360), .C(n_30274), .D
		(n_182284250), .Z(n_193784364));
	notech_ao4 i_98459722(.A(n_179784227), .B(\nbus_11290[0] ), .C(n_58238),
		 .D(n_179684226), .Z(n_193984366));
	notech_ao4 i_98259724(.A(n_382864359), .B(n_33169), .C(n_327760905), .D(n_383064361
		), .Z(n_194184368));
	notech_and4 i_98659720(.A(n_194184368), .B(n_193984366), .C(n_181484242)
		, .D(n_181784245), .Z(n_194384370));
	notech_ao4 i_97959727(.A(n_58051), .B(n_31472), .C(n_327660904), .D(n_57260
		), .Z(n_194484371));
	notech_and4 i_98159725(.A(n_327860906), .B(n_55802), .C(n_181184239), .D
		(n_194484371), .Z(n_194784374));
	notech_and2 i_98155933(.A(n_442368007), .B(n_29533), .Z(n_194884375));
	notech_or4 i_8255844(.A(n_32589), .B(n_28008), .C(n_63780), .D(n_61959),
		 .Z(n_194984376));
	notech_ao4 i_10355823(.A(n_32697), .B(n_30731), .C(n_29419), .D(n_30282)
		, .Z(n_195184378));
	notech_and3 i_10455822(.A(n_442368007), .B(n_29533), .C(n_57611), .Z(n_195284379
		));
	notech_and4 i_9555831(.A(n_284331524), .B(n_194984376), .C(n_27930), .D(n_215184571
		), .Z(n_195384380));
	notech_nand2 i_11755809(.A(tsc[26]), .B(n_30615), .Z(n_195484381));
	notech_or2 i_11655810(.A(n_131426641), .B(nbus_11271[26]), .Z(n_195784384
		));
	notech_nao3 i_11155815(.A(n_57395), .B(opd[26]), .C(n_58691), .Z(n_196284389
		));
	notech_nand2 i_12655800(.A(tsc[27]), .B(n_30615), .Z(n_196384390));
	notech_or2 i_12555801(.A(n_131426641), .B(nbus_11271[27]), .Z(n_196684393
		));
	notech_nao3 i_12055806(.A(n_57395), .B(opd[27]), .C(n_58691), .Z(n_197184398
		));
	notech_nand2 i_15755791(.A(tsc[28]), .B(n_30615), .Z(n_197284399));
	notech_or2 i_14155792(.A(n_131426641), .B(nbus_11271[28]), .Z(n_197584402
		));
	notech_nao3 i_12955797(.A(n_57395), .B(opd[28]), .C(n_58696), .Z(n_198084407
		));
	notech_or2 i_21855730(.A(n_25110), .B(nbus_11271[26]), .Z(n_198484411)
		);
	notech_nao3 i_21355735(.A(n_57395), .B(opd[26]), .C(n_57174), .Z(n_198984416
		));
	notech_nand2 i_22855720(.A(tsc[59]), .B(n_30615), .Z(n_199284419));
	notech_or2 i_22555723(.A(n_365528695), .B(\nbus_11290[27] ), .Z(n_199584422
		));
	notech_nao3 i_22255726(.A(n_57397), .B(opd[27]), .C(n_57174), .Z(n_199884425
		));
	notech_or2 i_23655712(.A(n_25110), .B(nbus_11271[28]), .Z(n_200284429)
		);
	notech_nand3 i_23155717(.A(n_57395), .B(n_32219), .C(opd[28]), .Z(n_200784434
		));
	notech_nand3 i_55155415(.A(n_55904), .B(n_171160315), .C(n_1759), .Z(n_201184437
		));
	notech_or2 i_54755418(.A(n_122726554), .B(\nbus_11283[26] ), .Z(n_201484440
		));
	notech_or2 i_54455421(.A(n_122826555), .B(n_33198), .Z(n_201784443));
	notech_nand2 i_54155424(.A(sav_edi[26]), .B(n_61861), .Z(n_202084446));
	notech_nand3 i_56355403(.A(n_55904), .B(n_171160315), .C(n_1761), .Z(n_202384449
		));
	notech_or2 i_56055406(.A(n_122726554), .B(\nbus_11283[27] ), .Z(n_202684452
		));
	notech_or2 i_55755409(.A(n_122826555), .B(n_33195), .Z(n_202984455));
	notech_nand2 i_55455412(.A(sav_edi[27]), .B(n_61861), .Z(n_203384458));
	notech_nand3 i_57555391(.A(n_55904), .B(n_171160315), .C(n_1763), .Z(n_203684461
		));
	notech_or2 i_57255394(.A(n_122726554), .B(\nbus_11283[28] ), .Z(n_203984464
		));
	notech_or2 i_56955397(.A(n_122826555), .B(n_33196), .Z(n_204284467));
	notech_nand2 i_56655400(.A(sav_edi[28]), .B(n_61861), .Z(n_204584470));
	notech_nor2 i_61155355(.A(n_28867), .B(nbus_11271[28]), .Z(n_204684471)
		);
	notech_nao3 i_60655360(.A(n_57395), .B(opd[28]), .C(n_57195), .Z(n_205384478
		));
	notech_or2 i_65955307(.A(n_327560903), .B(n_57057), .Z(n_205484479));
	notech_nao3 i_65455312(.A(n_63794), .B(opc[0]), .C(n_29333), .Z(n_206184486
		));
	notech_nao3 i_67855288(.A(n_57395), .B(opd[26]), .C(n_57057), .Z(n_206984494
		));
	notech_nand3 i_69455272(.A(n_57378), .B(n_32211), .C(opd[28]), .Z(n_207784502
		));
	notech_nor2 i_73155235(.A(n_443668020), .B(nbus_11271[28]), .Z(n_207884503
		));
	notech_and3 i_72655240(.A(n_57378), .B(n_32224), .C(opd[28]), .Z(n_208584510
		));
	notech_nor2 i_74755219(.A(n_443168015), .B(nbus_11271[26]), .Z(n_208684511
		));
	notech_nao3 i_74255224(.A(n_57378), .B(opd[26]), .C(n_57112), .Z(n_209384518
		));
	notech_nor2 i_75555211(.A(n_443168015), .B(nbus_11271[27]), .Z(n_209484519
		));
	notech_nao3 i_75055216(.A(n_57378), .B(opd[27]), .C(n_57112), .Z(n_210184526
		));
	notech_nor2 i_76355203(.A(n_443168015), .B(n_60564), .Z(n_210284527));
	notech_nand3 i_75855208(.A(n_57378), .B(n_125342694), .C(opd[28]), .Z(n_211184534
		));
	notech_ao3 i_77955187(.A(n_57378), .B(opd[26]), .C(n_57164), .Z(n_211284535
		));
	notech_nao3 i_77455192(.A(n_63770), .B(opc_10[26]), .C(n_442768011), .Z(n_211984542
		));
	notech_ao3 i_81755153(.A(n_57378), .B(opd[27]), .C(n_57164), .Z(n_212084543
		));
	notech_nao3 i_81155158(.A(opc_10[27]), .B(n_63780), .C(n_442768011), .Z(n_213084550
		));
	notech_nor2 i_82155150(.A(n_30693), .B(\nbus_11290[27] ), .Z(n_213484554
		));
	notech_and3 i_83055141(.A(n_57378), .B(n_32220), .C(opd[28]), .Z(n_213584555
		));
	notech_nao3 i_82555146(.A(n_63748), .B(opc_10[28]), .C(n_442768011), .Z(n_214284562
		));
	notech_nor2 i_83355138(.A(n_30693), .B(\nbus_11290[28] ), .Z(n_214784567
		));
	notech_or4 i_100054984(.A(n_61890), .B(n_195384380), .C(n_61718), .D(n_61861
		), .Z(n_214884568));
	notech_ao4 i_180571996(.A(n_27924), .B(n_60159), .C(n_60196), .D(n_32390
		), .Z(n_214984569));
	notech_and4 i_185954138(.A(n_27920), .B(n_27919), .C(n_316760795), .D(n_214984569
		), .Z(n_215184571));
	notech_ao4 i_170854288(.A(n_442868012), .B(n_60564), .C(n_440082450), .D
		(n_442968013), .Z(n_215584575));
	notech_ao4 i_170754289(.A(n_442568009), .B(\nbus_11290[28] ), .C(n_442668010
		), .D(\nbus_11283[28] ), .Z(n_215784577));
	notech_nand3 i_171054286(.A(n_215584575), .B(n_215784577), .C(n_214284562
		), .Z(n_215884578));
	notech_ao4 i_170554291(.A(n_117626503), .B(n_33196), .C(n_4427), .D(n_117726504
		), .Z(n_215984579));
	notech_ao4 i_171254284(.A(n_4427), .B(n_30689), .C(n_30697), .D(n_33196)
		, .Z(n_216084580));
	notech_ao4 i_171154285(.A(n_30695), .B(\nbus_11283[28] ), .C(n_31536), .D
		(n_61702), .Z(n_216284582));
	notech_nao3 i_52055919(.A(n_216084580), .B(n_216284582), .C(n_214784567)
		, .Z(n_216384583));
	notech_ao4 i_169754298(.A(n_442868012), .B(nbus_11271[27]), .C(n_284131522
		), .D(n_442968013), .Z(n_216684586));
	notech_ao4 i_169654299(.A(n_442568009), .B(n_58938), .C(n_442668010), .D
		(\nbus_11283[27] ), .Z(n_216884588));
	notech_nand3 i_170054296(.A(n_216684586), .B(n_216884588), .C(n_213084550
		), .Z(n_216984589));
	notech_ao4 i_169454301(.A(n_117626503), .B(n_33195), .C(n_5711), .D(n_117726504
		), .Z(n_217084590));
	notech_ao4 i_170254294(.A(n_5711), .B(n_30689), .C(n_30697), .D(n_33195)
		, .Z(n_217184591));
	notech_ao4 i_170154295(.A(n_31535), .B(n_61706), .C(n_30695), .D(\nbus_11283[27] 
		), .Z(n_217384593));
	notech_nao3 i_51955920(.A(n_217184591), .B(n_217384593), .C(n_213484554)
		, .Z(n_217484594));
	notech_ao4 i_162754365(.A(n_442868012), .B(nbus_11271[26]), .C(n_284231523
		), .D(n_442968013), .Z(n_217784597));
	notech_ao4 i_162654366(.A(n_442568009), .B(\nbus_11290[26] ), .C(n_442668010
		), .D(\nbus_11283[26] ), .Z(n_217984599));
	notech_nand3 i_162954363(.A(n_217784597), .B(n_217984599), .C(n_211984542
		), .Z(n_218084600));
	notech_ao4 i_162454368(.A(n_117626503), .B(n_33198), .C(n_5720), .D(n_117726504
		), .Z(n_218184601));
	notech_ao4 i_161354379(.A(n_440082450), .B(n_443468018), .C(n_7636), .D(n_443568019
		), .Z(n_218484604));
	notech_ao4 i_161254380(.A(n_4427), .B(n_118526512), .C(n_118426511), .D(n_33196
		), .Z(n_218684606));
	notech_nand3 i_161554377(.A(n_218484604), .B(n_218684606), .C(n_211184534
		), .Z(n_218784607));
	notech_ao4 i_161054382(.A(n_443268016), .B(\nbus_11283[28] ), .C(n_443368017
		), .D(n_58929), .Z(n_218884608));
	notech_ao4 i_160654386(.A(n_284131522), .B(n_443468018), .C(n_172669762)
		, .D(n_443568019), .Z(n_219184611));
	notech_ao4 i_160554387(.A(n_5711), .B(n_118526512), .C(n_118426511), .D(n_33195
		), .Z(n_219384613));
	notech_nand3 i_160854384(.A(n_219184611), .B(n_219384613), .C(n_210184526
		), .Z(n_219484614));
	notech_ao4 i_160354389(.A(n_443268016), .B(\nbus_11283[27] ), .C(n_443368017
		), .D(n_58938), .Z(n_219584615));
	notech_ao4 i_159954393(.A(n_284231523), .B(n_443468018), .C(n_175169787)
		, .D(n_443568019), .Z(n_219884618));
	notech_ao4 i_159854394(.A(n_5720), .B(n_118526512), .C(n_118426511), .D(n_33198
		), .Z(n_220084620));
	notech_nand3 i_160154391(.A(n_219884618), .B(n_220084620), .C(n_209384518
		), .Z(n_220184621));
	notech_ao4 i_159654396(.A(n_443268016), .B(\nbus_11283[26] ), .C(n_443368017
		), .D(\nbus_11290[26] ), .Z(n_220284622));
	notech_ao4 i_158554407(.A(n_440082450), .B(n_443968023), .C(n_7636), .D(n_444068024
		), .Z(n_220584625));
	notech_ao4 i_158454408(.A(n_4427), .B(n_119326520), .C(n_119226519), .D(n_33196
		), .Z(n_220784627));
	notech_nao3 i_158754405(.A(n_220584625), .B(n_220784627), .C(n_208584510
		), .Z(n_220884628));
	notech_ao4 i_158254410(.A(n_443768021), .B(n_58465), .C(n_443868022), .D
		(n_58929), .Z(n_220984629));
	notech_ao4 i_155154441(.A(n_440082450), .B(n_303822063), .C(n_7636), .D(n_299122016
		), .Z(n_221284632));
	notech_ao4 i_155054442(.A(n_4427), .B(n_57320), .C(n_57319), .D(n_33196)
		, .Z(n_221484634));
	notech_and3 i_155354439(.A(n_221284632), .B(n_221484634), .C(n_207784502
		), .Z(n_221584635));
	notech_ao4 i_154854444(.A(n_57363), .B(n_58465), .C(n_57362), .D(n_58929
		), .Z(n_221684636));
	notech_ao4 i_154754445(.A(n_31536), .B(n_61706), .C(n_303922064), .D(n_60564
		), .Z(n_221784637));
	notech_ao4 i_153654455(.A(n_284231523), .B(n_303822063), .C(n_175169787)
		, .D(n_299122016), .Z(n_221984639));
	notech_ao4 i_153554456(.A(n_5720), .B(n_57320), .C(n_57319), .D(n_33198)
		, .Z(n_222184641));
	notech_and3 i_153854453(.A(n_221984639), .B(n_222184641), .C(n_206984494
		), .Z(n_222284642));
	notech_ao4 i_153354458(.A(n_57363), .B(\nbus_11283[26] ), .C(n_57362), .D
		(\nbus_11290[26] ), .Z(n_222384643));
	notech_ao4 i_153254459(.A(n_31534), .B(n_61706), .C(n_303922064), .D(nbus_11271
		[26]), .Z(n_222484644));
	notech_ao4 i_147754513(.A(n_58956), .B(n_195284379), .C(n_58238), .D(n_30463
		), .Z(n_222684646));
	notech_ao4 i_147654514(.A(n_29540), .B(n_101142452), .C(n_29334), .D(n_327760905
		), .Z(n_222884648));
	notech_and3 i_147954511(.A(n_222684646), .B(n_222884648), .C(n_206184486
		), .Z(n_222984649));
	notech_ao4 i_147454516(.A(n_386464395), .B(n_56965), .C(n_29550), .D(n_33169
		), .Z(n_223084650));
	notech_ao4 i_143554555(.A(n_440082450), .B(n_28852), .C(n_7636), .D(n_28869
		), .Z(n_223384653));
	notech_ao4 i_143454556(.A(n_4427), .B(n_388264413), .C(n_388364414), .D(n_33196
		), .Z(n_223584655));
	notech_nand3 i_143754553(.A(n_223384653), .B(n_223584655), .C(n_205384478
		), .Z(n_223684656));
	notech_ao4 i_143254558(.A(n_28874), .B(n_58465), .C(n_28863), .D(n_58929
		), .Z(n_223784657));
	notech_ao4 i_140454586(.A(n_440082450), .B(n_122226549), .C(n_7636), .D(n_337461002
		), .Z(n_224084660));
	notech_ao4 i_140254588(.A(n_57001), .B(n_31536), .C(n_331060938), .D(n_31504
		), .Z(n_224284662));
	notech_and4 i_140654584(.A(n_224284662), .B(n_224084660), .C(n_204284467
		), .D(n_204584470), .Z(n_224484664));
	notech_ao4 i_139954591(.A(n_122626553), .B(n_58929), .C(n_4427), .D(n_122926556
		), .Z(n_224584665));
	notech_ao4 i_139754593(.A(n_55884), .B(n_33543), .C(n_337361001), .D(n_60564
		), .Z(n_224784667));
	notech_and4 i_140154589(.A(n_224784667), .B(n_224584665), .C(n_203684461
		), .D(n_203984464), .Z(n_224984669));
	notech_ao4 i_139454596(.A(n_284131522), .B(n_122226549), .C(n_172669762)
		, .D(n_337461002), .Z(n_225084670));
	notech_ao4 i_139254598(.A(n_57001), .B(n_31535), .C(n_331060938), .D(n_31503
		), .Z(n_225284672));
	notech_and4 i_139654594(.A(n_225284672), .B(n_225084670), .C(n_202984455
		), .D(n_203384458), .Z(n_225484674));
	notech_ao4 i_138954601(.A(n_122626553), .B(n_58938), .C(n_5711), .D(n_122926556
		), .Z(n_225584675));
	notech_ao4 i_138754603(.A(n_55884), .B(n_33542), .C(n_337361001), .D(nbus_11271
		[27]), .Z(n_225784677));
	notech_and4 i_139154599(.A(n_225784677), .B(n_225584675), .C(n_202384449
		), .D(n_202684452), .Z(n_225984679));
	notech_ao4 i_138454606(.A(n_284231523), .B(n_122226549), .C(n_175169787)
		, .D(n_337461002), .Z(n_226084680));
	notech_ao4 i_138254608(.A(n_57001), .B(n_31534), .C(n_331060938), .D(n_31502
		), .Z(n_226284682));
	notech_and4 i_138654604(.A(n_226284682), .B(n_226084680), .C(n_201784443
		), .D(n_202084446), .Z(n_226484684));
	notech_ao4 i_137954611(.A(n_122626553), .B(n_58911), .C(n_5720), .D(n_122926556
		), .Z(n_226584685));
	notech_ao4 i_137754613(.A(n_55884), .B(n_33541), .C(n_337361001), .D(n_60582
		), .Z(n_226784687));
	notech_and4 i_138154609(.A(n_226784687), .B(n_226584685), .C(n_201184437
		), .D(n_201484440), .Z(n_226984689));
	notech_ao4 i_111954869(.A(n_440082450), .B(n_25090), .C(n_7636), .D(n_365428694
		), .Z(n_227084690));
	notech_ao4 i_111854870(.A(n_4427), .B(n_365328693), .C(n_365228692), .D(n_33196
		), .Z(n_227284692));
	notech_and3 i_112154867(.A(n_200784434), .B(n_227084690), .C(n_227284692
		), .Z(n_227384693));
	notech_ao4 i_111554873(.A(n_365628696), .B(n_58465), .C(n_365528695), .D
		(n_58929), .Z(n_227484694));
	notech_ao4 i_111454874(.A(n_31536), .B(n_61706), .C(n_56030), .D(n_32579
		), .Z(n_227684696));
	notech_ao4 i_111154877(.A(n_284131522), .B(n_25090), .C(n_172669762), .D
		(n_365428694), .Z(n_227884698));
	notech_ao4 i_110954879(.A(n_5711), .B(n_365328693), .C(n_365228692), .D(n_33195
		), .Z(n_228084700));
	notech_and4 i_111354875(.A(n_228084700), .B(n_199884425), .C(n_227884698
		), .D(n_199584422), .Z(n_228284702));
	notech_ao4 i_110654882(.A(n_25110), .B(nbus_11271[27]), .C(n_365628696),
		 .D(n_58456), .Z(n_228384703));
	notech_and4 i_110854880(.A(n_55802), .B(n_228384703), .C(n_274331424), .D
		(n_199284419), .Z(n_228684706));
	notech_ao4 i_110254886(.A(n_284231523), .B(n_25090), .C(n_175169787), .D
		(n_365428694), .Z(n_228784707));
	notech_ao4 i_110154887(.A(n_5720), .B(n_365328693), .C(n_365228692), .D(n_33198
		), .Z(n_228984709));
	notech_and3 i_110454884(.A(n_198984416), .B(n_228784707), .C(n_228984709
		), .Z(n_229084710));
	notech_ao4 i_109854890(.A(n_365628696), .B(n_58447), .C(n_365528695), .D
		(n_58911), .Z(n_229184711));
	notech_ao4 i_109754891(.A(n_31534), .B(n_61706), .C(n_56030), .D(n_32578
		), .Z(n_229384713));
	notech_ao4 i_104754941(.A(n_440082450), .B(n_388064411), .C(n_7636), .D(n_388164412
		), .Z(n_229584715));
	notech_ao4 i_104654942(.A(n_4427), .B(n_131626643), .C(n_131526642), .D(n_33196
		), .Z(n_229784717));
	notech_ao4 i_104354945(.A(n_387864409), .B(n_58465), .C(n_387964410), .D
		(n_58929), .Z(n_229984719));
	notech_and4 i_104554943(.A(n_229984719), .B(n_197584402), .C(n_30506), .D
		(n_197284399), .Z(n_230284722));
	notech_ao4 i_103954949(.A(n_284131522), .B(n_388064411), .C(n_172669762)
		, .D(n_388164412), .Z(n_230384723));
	notech_ao4 i_103854950(.A(n_5711), .B(n_131626643), .C(n_131526642), .D(n_33195
		), .Z(n_230584725));
	notech_ao4 i_103554953(.A(n_387864409), .B(n_58456), .C(n_387964410), .D
		(n_58938), .Z(n_230784727));
	notech_and4 i_103754951(.A(n_230784727), .B(n_196684393), .C(n_30507), .D
		(n_196384390), .Z(n_231084730));
	notech_ao4 i_103154957(.A(n_284231523), .B(n_388064411), .C(n_175169787)
		, .D(n_388164412), .Z(n_231184731));
	notech_ao4 i_102954958(.A(n_5720), .B(n_131626643), .C(n_131526642), .D(n_33198
		), .Z(n_231384733));
	notech_ao4 i_102654961(.A(n_387864409), .B(n_58447), .C(n_387964410), .D
		(n_58911), .Z(n_231584735));
	notech_and4 i_102854959(.A(n_231584735), .B(n_195784384), .C(n_65029351)
		, .D(n_195484381), .Z(n_231884738));
	notech_or4 i_80852277(.A(n_58716), .B(n_32217), .C(n_57256), .D(n_363350926
		), .Z(n_231984739));
	notech_nao3 i_80952276(.A(n_63776), .B(opc_10[25]), .C(n_299122016), .Z(n_232684746
		));
	notech_nand3 i_2621016(.A(n_234084760), .B(n_232684746), .C(n_231984739)
		, .Z(n_18674));
	notech_or4 i_85652229(.A(n_58716), .B(n_32217), .C(n_57256), .D(n_3464),
		 .Z(n_232784747));
	notech_nao3 i_85752228(.A(opc_10[22]), .B(n_63758), .C(n_299122016), .Z(n_233484754
		));
	notech_nand3 i_2321013(.A(n_234784767), .B(n_233484754), .C(n_232784747)
		, .Z(n_18656));
	notech_ao4 i_81052275(.A(n_57363), .B(n_58438), .C(n_303922064), .D(n_60510
		), .Z(n_233584755));
	notech_ao4 i_81152274(.A(n_57320), .B(n_101026337), .C(n_57362), .D(n_58920
		), .Z(n_233784757));
	notech_ao4 i_81252273(.A(n_386864399), .B(n_31501), .C(n_57319), .D(n_33172
		), .Z(n_233884758));
	notech_and4 i_81552270(.A(n_233884758), .B(n_233784757), .C(n_233584755)
		, .D(n_350128600), .Z(n_234084760));
	notech_ao4 i_85852227(.A(n_57363), .B(n_58411), .C(n_303922064), .D(n_60537
		), .Z(n_234284762));
	notech_ao4 i_85952226(.A(n_57320), .B(n_59464), .C(n_57362), .D(n_58875)
		, .Z(n_234484764));
	notech_ao4 i_86052225(.A(n_386864399), .B(n_31496), .C(n_57319), .D(n_33284
		), .Z(n_234584765));
	notech_and4 i_86352222(.A(n_234584765), .B(n_234484764), .C(n_234284762)
		, .D(n_350328602), .Z(n_234784767));
	notech_nand2 i_5849671(.A(tsc[16]), .B(n_30615), .Z(n_234984769));
	notech_or2 i_5749672(.A(n_387964410), .B(\nbus_11290[16] ), .Z(n_235284772
		));
	notech_or2 i_5249677(.A(n_5444), .B(n_131626643), .Z(n_235784777));
	notech_and2 i_6749662(.A(tsc[17]), .B(n_30615), .Z(n_235884778));
	notech_nor2 i_6649663(.A(n_387964410), .B(\nbus_11290[17] ), .Z(n_236184781
		));
	notech_nor2 i_6149668(.A(n_5397), .B(n_131626643), .Z(n_236684786));
	notech_nand2 i_7649653(.A(tsc[18]), .B(n_30615), .Z(n_236784787));
	notech_or2 i_7549654(.A(n_387964410), .B(\nbus_11290[18] ), .Z(n_237084790
		));
	notech_or2 i_7049659(.A(n_5436), .B(n_131626643), .Z(n_237584795));
	notech_nand2 i_8549644(.A(tsc[19]), .B(n_30615), .Z(n_237684796));
	notech_or2 i_8449645(.A(n_387964410), .B(\nbus_11290[19] ), .Z(n_237984799
		));
	notech_or2 i_7949650(.A(n_5356), .B(n_131626643), .Z(n_238484804));
	notech_nand2 i_16949561(.A(tsc[48]), .B(n_30615), .Z(n_240184821));
	notech_or2 i_16649564(.A(n_365528695), .B(\nbus_11290[16] ), .Z(n_240484824
		));
	notech_nand3 i_16349567(.A(n_57378), .B(n_32219), .C(opd[16]), .Z(n_240784827
		));
	notech_or2 i_17749553(.A(n_25110), .B(nbus_11271[17]), .Z(n_241184831)
		);
	notech_nand3 i_17249558(.A(n_57378), .B(n_32219), .C(opd[17]), .Z(n_241684836
		));
	notech_nand2 i_18749543(.A(tsc[50]), .B(n_30615), .Z(n_241984839));
	notech_or2 i_18449546(.A(n_365528695), .B(\nbus_11290[18] ), .Z(n_242284842
		));
	notech_nand3 i_18149549(.A(n_57378), .B(n_32219), .C(opd[18]), .Z(n_242584845
		));
	notech_or2 i_19549535(.A(n_25110), .B(nbus_11271[19]), .Z(n_243084849)
		);
	notech_nand3 i_19049540(.A(n_57378), .B(n_32219), .C(opd[19]), .Z(n_243684854
		));
	notech_or2 i_20649524(.A(n_5783), .B(n_58784), .Z(n_244184859));
	notech_or4 i_20349527(.A(n_63716), .B(n_143769475), .C(n_61938), .D(nbus_11273
		[3]), .Z(n_244484862));
	notech_nand3 i_52149231(.A(n_55904), .B(n_171160315), .C(n_1739), .Z(n_245184869
		));
	notech_nand2 i_51849234(.A(sav_edi[16]), .B(n_61861), .Z(n_245484872));
	notech_or2 i_51549237(.A(n_122726554), .B(\nbus_11283[16] ), .Z(n_245784875
		));
	notech_or2 i_51249240(.A(n_320051171), .B(n_122226549), .Z(n_246084878)
		);
	notech_nand3 i_53349219(.A(n_55904), .B(n_171160315), .C(n_1741), .Z(n_246384881
		));
	notech_nand2 i_53049222(.A(sav_edi[17]), .B(n_61858), .Z(n_246684884));
	notech_or2 i_52749225(.A(n_122726554), .B(\nbus_11283[17] ), .Z(n_246984887
		));
	notech_or2 i_52449228(.A(n_319951172), .B(n_122226549), .Z(n_247284890)
		);
	notech_nand3 i_54549207(.A(n_55904), .B(n_171160315), .C(n_1743), .Z(n_247584893
		));
	notech_nand2 i_54249210(.A(sav_edi[18]), .B(n_61858), .Z(n_247884896));
	notech_or2 i_53949213(.A(n_122726554), .B(\nbus_11283[18] ), .Z(n_248184899
		));
	notech_or2 i_53649216(.A(n_319825274), .B(n_122226549), .Z(n_248484902)
		);
	notech_nand3 i_55749195(.A(n_55904), .B(n_171160315), .C(n_1745), .Z(n_248784905
		));
	notech_nand2 i_55449198(.A(sav_edi[19]), .B(n_61858), .Z(n_249084908));
	notech_or2 i_55149201(.A(n_122726554), .B(\nbus_11283[19] ), .Z(n_249384911
		));
	notech_or2 i_54849204(.A(n_319725273), .B(n_122226549), .Z(n_249684914)
		);
	notech_or4 i_60849144(.A(n_63716), .B(n_169676762), .C(n_61938), .D(nbus_11273
		[3]), .Z(n_250584923));
	notech_or4 i_65349099(.A(n_63716), .B(n_29342), .C(n_61938), .D(n_58256)
		, .Z(n_251984936));
	notech_and3 i_75548997(.A(n_57378), .B(n_125342694), .C(opd[16]), .Z(n_252484941
		));
	notech_or2 i_75049002(.A(n_443168015), .B(nbus_11271[16]), .Z(n_253184948
		));
	notech_and3 i_76348989(.A(n_57395), .B(n_125342694), .C(opd[17]), .Z(n_253284949
		));
	notech_or2 i_75848994(.A(n_443168015), .B(nbus_11271[17]), .Z(n_253984956
		));
	notech_and3 i_77148981(.A(n_57395), .B(n_125342694), .C(opd[18]), .Z(n_254084957
		));
	notech_or2 i_76648986(.A(n_443168015), .B(nbus_11271[18]), .Z(n_254784964
		));
	notech_and3 i_77948973(.A(n_57395), .B(n_125342694), .C(opd[19]), .Z(n_254884965
		));
	notech_or2 i_77448978(.A(n_443168015), .B(nbus_11271[19]), .Z(n_255584972
		));
	notech_nor2 i_80448948(.A(n_442868012), .B(nbus_11271[16]), .Z(n_255684973
		));
	notech_nand3 i_79948953(.A(n_57395), .B(n_32220), .C(opd[16]), .Z(n_256384980
		));
	notech_or4 i_80748945(.A(n_335660984), .B(n_61630), .C(n_32317), .D(n_33199
		), .Z(n_256784984));
	notech_nor2 i_81648936(.A(n_442868012), .B(nbus_11271[17]), .Z(n_256884985
		));
	notech_and3 i_81148941(.A(n_57395), .B(n_32220), .C(opd[17]), .Z(n_257584992
		));
	notech_nor2 i_81948933(.A(n_30697), .B(n_33200), .Z(n_257984996));
	notech_nor2 i_82848924(.A(n_442868012), .B(nbus_11271[18]), .Z(n_258084997
		));
	notech_and3 i_82348929(.A(n_57395), .B(n_32220), .C(opd[18]), .Z(n_258785004
		));
	notech_nor2 i_83148921(.A(n_30697), .B(n_33201), .Z(n_259185008));
	notech_nor2 i_84048912(.A(n_442868012), .B(nbus_11271[19]), .Z(n_259285009
		));
	notech_and3 i_83548917(.A(n_57392), .B(n_32220), .C(opd[19]), .Z(n_259985016
		));
	notech_nor2 i_84448909(.A(n_30697), .B(n_33202), .Z(n_260385020));
	notech_ao4 i_190847885(.A(n_319725273), .B(n_442968013), .C(n_232870324)
		, .D(n_442768011), .Z(n_260485021));
	notech_ao4 i_190747886(.A(n_5356), .B(n_117726504), .C(n_117626503), .D(n_33202
		), .Z(n_260685023));
	notech_nao3 i_191047883(.A(n_260485021), .B(n_260685023), .C(n_259985016
		), .Z(n_260785024));
	notech_ao4 i_190547888(.A(n_442668010), .B(\nbus_11283[19] ), .C(n_442568009
		), .D(\nbus_11290[19] ), .Z(n_260885025));
	notech_ao4 i_191247881(.A(n_30693), .B(\nbus_11290[19] ), .C(n_30695), .D
		(\nbus_11283[19] ), .Z(n_260985026));
	notech_ao4 i_191147882(.A(n_61702), .B(n_31527), .C(n_5356), .D(n_30689)
		, .Z(n_261185028));
	notech_nao3 i_51149731(.A(n_260985026), .B(n_261185028), .C(n_260385020)
		, .Z(n_261285029));
	notech_ao4 i_189847895(.A(n_319825274), .B(n_442968013), .C(n_235370349)
		, .D(n_442768011), .Z(n_261585032));
	notech_ao4 i_189747896(.A(n_5436), .B(n_117726504), .C(n_117626503), .D(n_33201
		), .Z(n_261785034));
	notech_nao3 i_190047893(.A(n_261585032), .B(n_261785034), .C(n_258785004
		), .Z(n_261885035));
	notech_ao4 i_189547898(.A(n_442668010), .B(\nbus_11283[18] ), .C(n_442568009
		), .D(\nbus_11290[18] ), .Z(n_261985036));
	notech_ao4 i_190247891(.A(n_30693), .B(\nbus_11290[18] ), .C(n_30695), .D
		(\nbus_11283[18] ), .Z(n_262085037));
	notech_ao4 i_190147892(.A(n_61702), .B(n_31526), .C(n_5436), .D(n_30689)
		, .Z(n_262285039));
	notech_nao3 i_51049732(.A(n_262085037), .B(n_262285039), .C(n_259185008)
		, .Z(n_262385040));
	notech_ao4 i_188847905(.A(n_319951172), .B(n_442968013), .C(n_237870374)
		, .D(n_442768011), .Z(n_262685043));
	notech_ao4 i_188747906(.A(n_5397), .B(n_117726504), .C(n_33200), .D(n_117626503
		), .Z(n_262885045));
	notech_nao3 i_189047903(.A(n_262685043), .B(n_262885045), .C(n_257584992
		), .Z(n_262985046));
	notech_ao4 i_188547908(.A(n_442668010), .B(\nbus_11283[17] ), .C(n_442568009
		), .D(\nbus_11290[17] ), .Z(n_263085047));
	notech_ao4 i_189247901(.A(n_30693), .B(\nbus_11290[17] ), .C(n_30695), .D
		(\nbus_11283[17] ), .Z(n_263185048));
	notech_ao4 i_189147902(.A(n_61702), .B(n_31525), .C(n_5397), .D(n_30689)
		, .Z(n_263385050));
	notech_nao3 i_50949733(.A(n_263185048), .B(n_263385050), .C(n_257984996)
		, .Z(n_263485051));
	notech_ao4 i_187847915(.A(n_320051171), .B(n_442968013), .C(n_240370399)
		, .D(n_442768011), .Z(n_263785054));
	notech_ao4 i_187747916(.A(n_5444), .B(n_117726504), .C(n_117626503), .D(n_33199
		), .Z(n_263985056));
	notech_nand3 i_188047913(.A(n_263785054), .B(n_263985056), .C(n_256384980
		), .Z(n_264085057));
	notech_ao4 i_187547918(.A(n_442668010), .B(\nbus_11283[16] ), .C(n_442568009
		), .D(\nbus_11290[16] ), .Z(n_264185058));
	notech_ao4 i_188247911(.A(n_30693), .B(n_59059), .C(n_30695), .D(\nbus_11283[16] 
		), .Z(n_264285059));
	notech_ao4 i_188147912(.A(n_31524), .B(n_61702), .C(n_5444), .D(n_30689)
		, .Z(n_264485061));
	notech_nand3 i_50849734(.A(n_264285059), .B(n_264485061), .C(n_256784984
		), .Z(n_264585062));
	notech_ao4 i_185747936(.A(n_443268016), .B(\nbus_11283[19] ), .C(n_443368017
		), .D(n_58866), .Z(n_264885065));
	notech_ao4 i_185647937(.A(n_232870324), .B(n_443568019), .C(n_57112), .D
		(n_305478064), .Z(n_265085067));
	notech_nand3 i_185947934(.A(n_264885065), .B(n_265085067), .C(n_255584972
		), .Z(n_265185068));
	notech_ao4 i_185447939(.A(n_118426511), .B(n_33202), .C(n_5356), .D(n_118526512
		), .Z(n_265285069));
	notech_ao4 i_185047943(.A(n_443268016), .B(\nbus_11283[18] ), .C(n_443368017
		), .D(n_59077), .Z(n_265585072));
	notech_or2 i_549720(.A(n_319825274), .B(n_57256), .Z(n_265785074));
	notech_ao4 i_184947944(.A(n_235370349), .B(n_443568019), .C(n_57112), .D
		(n_265785074), .Z(n_265885075));
	notech_nand3 i_185247941(.A(n_265585072), .B(n_265885075), .C(n_254784964
		), .Z(n_265985076));
	notech_ao4 i_184747946(.A(n_118426511), .B(n_33201), .C(n_5436), .D(n_118526512
		), .Z(n_266085077));
	notech_ao4 i_184347950(.A(n_443268016), .B(\nbus_11283[17] ), .C(n_443368017
		), .D(n_59086), .Z(n_266385080));
	notech_or2 i_1249713(.A(n_319951172), .B(n_57256), .Z(n_266585082));
	notech_ao4 i_184247951(.A(n_237870374), .B(n_443568019), .C(n_57112), .D
		(n_266585082), .Z(n_266685083));
	notech_nand3 i_184547948(.A(n_266385080), .B(n_266685083), .C(n_253984956
		), .Z(n_266785084));
	notech_ao4 i_184047953(.A(n_33200), .B(n_118426511), .C(n_5397), .D(n_118526512
		), .Z(n_266885085));
	notech_ao4 i_183647957(.A(n_443268016), .B(\nbus_11283[16] ), .C(n_443368017
		), .D(n_59059), .Z(n_267185088));
	notech_or2 i_749718(.A(n_320051171), .B(n_57256), .Z(n_267385090));
	notech_ao4 i_183547958(.A(n_240370399), .B(n_443568019), .C(n_267385090)
		, .D(n_57112), .Z(n_267485091));
	notech_nand3 i_183847955(.A(n_267185088), .B(n_267485091), .C(n_253184948
		), .Z(n_267585092));
	notech_ao4 i_183347960(.A(n_118426511), .B(n_33199), .C(n_5444), .D(n_118526512
		), .Z(n_267685093));
	notech_ao4 i_175148042(.A(n_74922852), .B(n_29333), .C(n_66222765), .D(n_57057
		), .Z(n_267985096));
	notech_ao4 i_175048043(.A(n_29337), .B(n_75322856), .C(n_29341), .D(n_75222855
		), .Z(n_268085097));
	notech_ao4 i_174848045(.A(n_29340), .B(n_75522858), .C(n_29338), .D(n_75622859
		), .Z(n_268285099));
	notech_and4 i_175348040(.A(n_268285099), .B(n_268085097), .C(n_267985096
		), .D(n_251984936), .Z(n_268485101));
	notech_ao4 i_174548048(.A(n_74522848), .B(n_29334), .C(n_74622849), .D(n_378364314
		), .Z(n_268585102));
	notech_ao4 i_174448049(.A(n_338361011), .B(n_29540), .C(n_386464395), .D
		(n_58784), .Z(n_268685103));
	notech_ao4 i_174248051(.A(n_29533), .B(\nbus_11290[3] ), .C(n_29550), .D
		(n_33118), .Z(n_268885105));
	notech_and4 i_174748046(.A(n_65022753), .B(n_268885105), .C(n_268685103)
		, .D(n_268585102), .Z(n_269085107));
	notech_ao4 i_171148082(.A(n_200477060), .B(n_74922852), .C(n_66222765), 
		.D(n_57604), .Z(n_269185108));
	notech_ao4 i_171048083(.A(n_140076466), .B(n_75322856), .C(n_139976465),
		 .D(n_75222855), .Z(n_269285109));
	notech_ao4 i_170848085(.A(n_139876464), .B(n_75522858), .C(n_140176467),
		 .D(n_75622859), .Z(n_269485111));
	notech_and4 i_171348080(.A(n_269485111), .B(n_269285109), .C(n_269185108
		), .D(n_250584923), .Z(n_269685113));
	notech_ao4 i_170548088(.A(n_200377059), .B(n_74522848), .C(n_57666), .D(n_74622849
		), .Z(n_269785114));
	notech_ao4 i_170448089(.A(n_323278241), .B(n_338361011), .C(n_58044), .D
		(n_58784), .Z(n_269885115));
	notech_ao4 i_170248091(.A(n_279977810), .B(nbus_11271[3]), .C(n_192676984
		), .D(n_33118), .Z(n_270085117));
	notech_and4 i_170748086(.A(n_65022753), .B(n_270085117), .C(n_269885115)
		, .D(n_269785114), .Z(n_270285119));
	notech_ao4 i_166048133(.A(n_232870324), .B(n_337461002), .C(n_337361001)
		, .D(nbus_11271[19]), .Z(n_270385120));
	notech_ao4 i_165848135(.A(n_122826555), .B(n_33202), .C(n_5356), .D(n_122926556
		), .Z(n_270585122));
	notech_and4 i_166248131(.A(n_270585122), .B(n_270385120), .C(n_249384911
		), .D(n_249684914), .Z(n_270785124));
	notech_ao4 i_165548138(.A(n_331060938), .B(n_31492), .C(n_122626553), .D
		(n_58866), .Z(n_270985125));
	notech_ao4 i_165348140(.A(n_55884), .B(n_33547), .C(n_57001), .D(n_31527
		), .Z(n_271185127));
	notech_and4 i_165748136(.A(n_271185127), .B(n_270985125), .C(n_248784905
		), .D(n_249084908), .Z(n_271385129));
	notech_ao4 i_165048143(.A(n_235370349), .B(n_337461002), .C(n_337361001)
		, .D(nbus_11271[18]), .Z(n_271485130));
	notech_ao4 i_164848145(.A(n_122826555), .B(n_33201), .C(n_5436), .D(n_122926556
		), .Z(n_271785132));
	notech_and4 i_165248141(.A(n_271785132), .B(n_271485130), .C(n_248184899
		), .D(n_248484902), .Z(n_271985134));
	notech_ao4 i_164548148(.A(n_331060938), .B(n_31491), .C(n_122626553), .D
		(n_59077), .Z(n_272085135));
	notech_ao4 i_164348150(.A(n_55884), .B(n_33546), .C(n_57001), .D(n_31526
		), .Z(n_272385137));
	notech_and4 i_164748146(.A(n_272385137), .B(n_272085135), .C(n_247584893
		), .D(n_247884896), .Z(n_272585139));
	notech_ao4 i_164048153(.A(n_237870374), .B(n_337461002), .C(n_337361001)
		, .D(nbus_11271[17]), .Z(n_272685140));
	notech_ao4 i_163848155(.A(n_33200), .B(n_122826555), .C(n_5397), .D(n_122926556
		), .Z(n_272885142));
	notech_and4 i_164248151(.A(n_272885142), .B(n_272685140), .C(n_246984887
		), .D(n_247284890), .Z(n_273085144));
	notech_ao4 i_163548158(.A(n_331060938), .B(n_31490), .C(n_122626553), .D
		(n_59086), .Z(n_273185145));
	notech_ao4 i_163348160(.A(n_55884), .B(n_33545), .C(n_57001), .D(n_31525
		), .Z(n_273385147));
	notech_and4 i_163748156(.A(n_273385147), .B(n_273185145), .C(n_246384881
		), .D(n_246684884), .Z(n_273585149));
	notech_ao4 i_163048163(.A(n_240370399), .B(n_337461002), .C(n_337361001)
		, .D(nbus_11271[16]), .Z(n_273685150));
	notech_ao4 i_162848165(.A(n_122826555), .B(n_33199), .C(n_5444), .D(n_122926556
		), .Z(n_273885152));
	notech_and4 i_163248161(.A(n_273885152), .B(n_273685150), .C(n_245784875
		), .D(n_246084878), .Z(n_274085154));
	notech_ao4 i_162548168(.A(n_331060938), .B(n_31489), .C(n_122626553), .D
		(n_59059), .Z(n_274185155));
	notech_ao4 i_162348170(.A(n_55884), .B(n_33544), .C(n_57006), .D(n_31524
		), .Z(n_274385157));
	notech_and4 i_162748166(.A(n_274385157), .B(n_274185155), .C(n_245184869
		), .D(n_245484872), .Z(n_274585159));
	notech_ao4 i_137448413(.A(n_74922852), .B(n_151069548), .C(n_66222765), 
		.D(n_57068), .Z(n_274685160));
	notech_ao4 i_137348414(.A(n_75322856), .B(n_143469472), .C(n_75222855), 
		.D(n_143569473), .Z(n_274785161));
	notech_ao4 i_137148416(.A(n_75522858), .B(n_143669474), .C(n_75622859), 
		.D(n_143369471), .Z(n_274985163));
	notech_and4 i_137648411(.A(n_274985163), .B(n_274785161), .C(n_274685160
		), .D(n_244484862), .Z(n_275185165));
	notech_ao4 i_136848419(.A(n_74522848), .B(n_150969547), .C(n_74622849), 
		.D(n_57438), .Z(n_275285166));
	notech_ao4 i_136648421(.A(n_33118), .B(n_57027), .C(n_338361011), .D(n_57036
		), .Z(n_275485168));
	notech_and4 i_137048417(.A(n_65022753), .B(n_275485168), .C(n_275285166)
		, .D(n_244184859), .Z(n_275685170));
	notech_ao4 i_136348424(.A(n_319725273), .B(n_25090), .C(n_232870324), .D
		(n_365428694), .Z(n_275785171));
	notech_ao4 i_136148425(.A(n_5356), .B(n_365328693), .C(n_365228692), .D(n_33202
		), .Z(n_275985173));
	notech_and3 i_136548422(.A(n_243684854), .B(n_275785171), .C(n_275985173
		), .Z(n_276085174));
	notech_ao4 i_135848428(.A(n_365628696), .B(n_58384), .C(n_365528695), .D
		(n_58866), .Z(n_276185175));
	notech_ao4 i_135748429(.A(n_31527), .B(n_61702), .C(n_56030), .D(n_32569
		), .Z(n_276385177));
	notech_ao4 i_135448432(.A(n_319825274), .B(n_25090), .C(n_235370349), .D
		(n_365428694), .Z(n_276585179));
	notech_ao4 i_135248434(.A(n_5436), .B(n_365328693), .C(n_365228692), .D(n_33201
		), .Z(n_276785181));
	notech_and4 i_135648430(.A(n_276785181), .B(n_242584845), .C(n_276585179
		), .D(n_242284842), .Z(n_276985183));
	notech_ao4 i_134948437(.A(n_25110), .B(nbus_11271[18]), .C(n_365628696),
		 .D(n_58375), .Z(n_277085184));
	notech_and4 i_135148435(.A(n_55802), .B(n_277085184), .C(n_314325220), .D
		(n_241984839), .Z(n_277385187));
	notech_ao4 i_134548441(.A(n_319951172), .B(n_25090), .C(n_237870374), .D
		(n_365428694), .Z(n_277485188));
	notech_ao4 i_134448442(.A(n_5397), .B(n_365328693), .C(n_365228692), .D(n_33200
		), .Z(n_277685190));
	notech_and3 i_134748439(.A(n_241684836), .B(n_277485188), .C(n_277685190
		), .Z(n_277785191));
	notech_ao4 i_134148445(.A(n_365628696), .B(n_58366), .C(n_365528695), .D
		(n_59086), .Z(n_277885192));
	notech_ao4 i_134048446(.A(n_31525), .B(n_61702), .C(n_56030), .D(n_32568
		), .Z(n_278085194));
	notech_ao4 i_133748449(.A(n_320051171), .B(n_25090), .C(n_240370399), .D
		(n_365428694), .Z(n_278285196));
	notech_ao4 i_133548451(.A(n_5444), .B(n_365328693), .C(n_365228692), .D(n_33199
		), .Z(n_278485198));
	notech_and4 i_133948447(.A(n_278485198), .B(n_278285196), .C(n_240484824
		), .D(n_240784827), .Z(n_278685200));
	notech_ao4 i_133248454(.A(n_25110), .B(nbus_11271[16]), .C(n_365628696),
		 .D(n_58357), .Z(n_278785201));
	notech_and4 i_133448452(.A(n_55802), .B(n_278785201), .C(n_314525222), .D
		(n_240184821), .Z(n_279085204));
	notech_ao4 i_132348458(.A(n_74922852), .B(n_57260), .C(n_66222765), .D(n_57174
		), .Z(n_279185205));
	notech_ao4 i_132248459(.A(n_75322856), .B(n_179284222), .C(n_75222855), 
		.D(n_179484224), .Z(n_279285206));
	notech_ao4 i_132048461(.A(n_75522858), .B(n_179584225), .C(n_75622859), 
		.D(n_179384223), .Z(n_279485208));
	notech_ao4 i_131948462(.A(n_74622849), .B(n_57383), .C(n_188084307), .D(n_74822851
		), .Z(n_279585209));
	notech_and4 i_132648456(.A(n_279585209), .B(n_279485208), .C(n_279285206
		), .D(n_279185205), .Z(n_279785211));
	notech_ao4 i_131648465(.A(n_58051), .B(n_58784), .C(n_74522848), .D(n_383064361
		), .Z(n_279885212));
	notech_ao4 i_131548466(.A(n_33118), .B(n_382864359), .C(n_338361011), .D
		(n_382664357), .Z(n_279985213));
	notech_ao4 i_131348468(.A(n_56030), .B(n_32555), .C(n_58664), .D(\nbus_11290[3] 
		), .Z(n_280185215));
	notech_and3 i_131448467(.A(n_65022753), .B(n_55802), .C(n_280185215), .Z
		(n_280385217));
	notech_ao4 i_125548526(.A(n_232870324), .B(n_388164412), .C(n_305478064)
		, .D(n_58691), .Z(n_280585219));
	notech_ao4 i_125448527(.A(n_131426641), .B(nbus_11271[19]), .C(n_131526642
		), .D(n_33202), .Z(n_280785221));
	notech_ao4 i_125148530(.A(n_387864409), .B(n_58384), .C(n_390064431), .D
		(n_31492), .Z(n_280985223));
	notech_and4 i_125348528(.A(n_237984799), .B(n_280985223), .C(n_30510), .D
		(n_237684796), .Z(n_281285226));
	notech_ao4 i_124748534(.A(n_235370349), .B(n_388164412), .C(n_58691), .D
		(n_265785074), .Z(n_281385227));
	notech_ao4 i_124648535(.A(n_131426641), .B(nbus_11271[18]), .C(n_131526642
		), .D(n_33201), .Z(n_281585229));
	notech_ao4 i_124348538(.A(n_387864409), .B(n_58375), .C(n_390064431), .D
		(n_31491), .Z(n_281785231));
	notech_and4 i_124548536(.A(n_237084790), .B(n_281785231), .C(n_30511), .D
		(n_236784787), .Z(n_282085234));
	notech_ao4 i_123948542(.A(n_237870374), .B(n_388164412), .C(n_58691), .D
		(n_266585082), .Z(n_282185235));
	notech_ao4 i_123848543(.A(n_131426641), .B(nbus_11271[17]), .C(n_131526642
		), .D(n_33200), .Z(n_282385237));
	notech_ao4 i_123548546(.A(n_387864409), .B(n_58366), .C(n_390064431), .D
		(n_31490), .Z(n_282585239));
	notech_or4 i_123748544(.A(n_235884778), .B(n_263485051), .C(n_236184781)
		, .D(n_30487), .Z(n_282885242));
	notech_ao4 i_123148550(.A(n_240370399), .B(n_388164412), .C(n_58691), .D
		(n_267385090), .Z(n_282985243));
	notech_ao4 i_123048551(.A(n_131426641), .B(nbus_11271[16]), .C(n_131526642
		), .D(n_33199), .Z(n_283185245));
	notech_ao4 i_122748554(.A(n_387864409), .B(n_58357), .C(n_390064431), .D
		(n_31489), .Z(n_283385247));
	notech_and4 i_122948552(.A(n_283385247), .B(n_234984769), .C(n_235284772
		), .D(n_30513), .Z(n_283685250));
	notech_nand2 i_5546357(.A(tsc[31]), .B(n_30615), .Z(n_283785251));
	notech_or2 i_5446358(.A(n_131426641), .B(nbus_11271[31]), .Z(n_284085254
		));
	notech_nao3 i_4946363(.A(n_57392), .B(opd[31]), .C(n_58691), .Z(n_284585259
		));
	notech_nao3 i_35646062(.A(n_3480), .B(n_61286), .C(n_32186), .Z(n_284885262
		));
	notech_or4 i_34946069(.A(n_61858), .B(n_61702), .C(n_19680), .D(n_31516)
		, .Z(n_285585269));
	notech_or2 i_38646032(.A(n_25110), .B(nbus_11271[31]), .Z(n_286385277)
		);
	notech_nand3 i_38146037(.A(n_57392), .B(n_32219), .C(opd[31]), .Z(n_286885282
		));
	notech_or2 i_42145998(.A(n_55955), .B(n_30983), .Z(n_287185285));
	notech_nand3 i_52945904(.A(n_55904), .B(n_171160315), .C(n_1723), .Z(n_288685300
		));
	notech_or2 i_52145911(.A(n_5269), .B(n_444668030), .Z(n_289385307));
	notech_nand3 i_54145892(.A(n_1769), .B(n_55904), .C(n_171160315), .Z(n_290085314
		));
	notech_or2 i_53845895(.A(n_122726554), .B(\nbus_11283[31] ), .Z(n_290385317
		));
	notech_or2 i_53545898(.A(n_122826555), .B(n_33206), .Z(n_290685320));
	notech_nand2 i_53245901(.A(sav_edi[31]), .B(n_61858), .Z(n_290985323));
	notech_nor2 i_65645781(.A(n_443168015), .B(nbus_11271[31]), .Z(n_291085324
		));
	notech_nand3 i_65145786(.A(n_57392), .B(n_125342694), .C(opd[31]), .Z(n_291785331
		));
	notech_nor2 i_67945758(.A(n_442868012), .B(n_60591), .Z(n_291885332));
	notech_and3 i_67445763(.A(n_57392), .B(n_32220), .C(opd[31]), .Z(n_292585339
		));
	notech_nor2 i_68245755(.A(n_30693), .B(\nbus_11290[31] ), .Z(n_292985343
		));
	notech_ao4 i_174444769(.A(n_300822033), .B(n_442968013), .C(n_262470619)
		, .D(n_442768011), .Z(n_293085344));
	notech_ao4 i_174344770(.A(n_5243), .B(n_117726504), .C(n_117626503), .D(n_33206
		), .Z(n_293285346));
	notech_nao3 i_174644767(.A(n_293085344), .B(n_293285346), .C(n_292585339
		), .Z(n_293385347));
	notech_ao4 i_174144772(.A(n_442668010), .B(n_60458), .C(n_442568009), .D
		(\nbus_11290[31] ), .Z(n_293485348));
	notech_ao4 i_174844765(.A(n_5243), .B(n_30689), .C(n_30697), .D(n_33206)
		, .Z(n_293585349));
	notech_ao4 i_174744766(.A(n_31539), .B(n_61702), .C(n_30695), .D(n_60458
		), .Z(n_293785351));
	notech_nao3 i_52346422(.A(n_293585349), .B(n_293785351), .C(n_292985343)
		, .Z(n_293885352));
	notech_ao4 i_172544788(.A(n_300822033), .B(n_443468018), .C(n_262470619)
		, .D(n_443568019), .Z(n_294185355));
	notech_ao4 i_172444789(.A(n_5243), .B(n_118526512), .C(n_118426511), .D(n_33206
		), .Z(n_294385357));
	notech_nand3 i_172744786(.A(n_294185355), .B(n_294385357), .C(n_291785331
		), .Z(n_294485358));
	notech_ao4 i_172244791(.A(n_443268016), .B(n_60458), .C(n_443368017), .D
		(n_58983), .Z(n_294585359));
	notech_ao4 i_156744942(.A(n_300822033), .B(n_122226549), .C(n_262470619)
		, .D(n_337461002), .Z(n_294885362));
	notech_ao4 i_156544944(.A(n_57006), .B(n_31539), .C(n_331060938), .D(n_31507
		), .Z(n_295085364));
	notech_and4 i_156944940(.A(n_295085364), .B(n_294885362), .C(n_290685320
		), .D(n_290985323), .Z(n_295285366));
	notech_ao4 i_156244947(.A(n_122626553), .B(n_58983), .C(n_5243), .D(n_122926556
		), .Z(n_295385367));
	notech_ao4 i_155944949(.A(n_55884), .B(n_33551), .C(n_337361001), .D(n_60591
		), .Z(n_295585369));
	notech_and4 i_156444945(.A(n_295585369), .B(n_295385367), .C(n_290085314
		), .D(n_290385317), .Z(n_295785371));
	notech_ao4 i_155644952(.A(n_28368), .B(n_266870661), .C(n_266970662), .D
		(n_28367), .Z(n_295885372));
	notech_ao4 i_155544953(.A(n_267170664), .B(n_28365), .C(n_444768031), .D
		(n_267470667), .Z(n_295985373));
	notech_ao4 i_155344955(.A(n_444868032), .B(n_31481), .C(n_300722032), .D
		(n_331760945), .Z(n_296185375));
	notech_and4 i_155844950(.A(n_296185375), .B(n_295985373), .C(n_295885372
		), .D(n_289385307), .Z(n_296385377));
	notech_ao4 i_155044958(.A(n_444468028), .B(\nbus_11290[8] ), .C(n_444568029
		), .D(n_33253), .Z(n_296485378));
	notech_ao4 i_154944959(.A(n_61091), .B(n_30843), .C(n_444368027), .D(nbus_11273
		[8]), .Z(n_296585379));
	notech_ao4 i_154744961(.A(n_55884), .B(n_33550), .C(n_57006), .D(n_31516
		), .Z(n_296785381));
	notech_and4 i_155244956(.A(n_296785381), .B(n_296585379), .C(n_296485378
		), .D(n_288685300), .Z(n_296985383));
	notech_ao4 i_147545031(.A(n_26397), .B(n_266870661), .C(n_266970662), .D
		(n_26394), .Z(n_297085384));
	notech_ao4 i_147345032(.A(n_267170664), .B(n_26396), .C(n_378564316), .D
		(n_267470667), .Z(n_297185385));
	notech_ao4 i_147145034(.A(n_61087), .B(n_30784), .C(n_331560943), .D(n_300722032
		), .Z(n_297385387));
	notech_ao4 i_147045035(.A(n_378464315), .B(n_31481), .C(n_55946), .D(n_31516
		), .Z(n_297485388));
	notech_and4 i_147745029(.A(n_297485388), .B(n_297385387), .C(n_297185385
		), .D(n_297085384), .Z(n_297685390));
	notech_ao4 i_146645038(.A(n_378664317), .B(\nbus_11290[8] ), .C(n_378764318
		), .D(nbus_11273[8]), .Z(n_297785391));
	notech_ao4 i_146545039(.A(n_378964320), .B(n_33253), .C(n_5269), .D(n_378864319
		), .Z(n_297885392));
	notech_ao4 i_146345041(.A(n_55975), .B(n_32067), .C(n_125926586), .D(n_33549
		), .Z(n_298085394));
	notech_and4 i_146945036(.A(n_298085394), .B(n_297885392), .C(n_297785391
		), .D(n_287185285), .Z(n_298285396));
	notech_ao4 i_144345061(.A(n_300822033), .B(n_25090), .C(n_262470619), .D
		(n_365428694), .Z(n_298385397));
	notech_ao4 i_144245062(.A(n_5243), .B(n_365328693), .C(n_365228692), .D(n_33206
		), .Z(n_298585399));
	notech_and3 i_144545059(.A(n_286885282), .B(n_298385397), .C(n_298585399
		), .Z(n_298685400));
	notech_ao4 i_143945065(.A(n_365628696), .B(n_60458), .C(n_365528695), .D
		(n_58983), .Z(n_298785401));
	notech_ao4 i_143845066(.A(n_31539), .B(n_61702), .C(n_56035), .D(n_32582
		), .Z(n_298985403));
	notech_ao4 i_140845088(.A(n_266870661), .B(n_24542), .C(n_266970662), .D
		(n_24541), .Z(n_299185405));
	notech_ao4 i_140745089(.A(n_267170664), .B(n_24539), .C(n_267470667), .D
		(n_381564346), .Z(n_299285406));
	notech_ao4 i_140545091(.A(n_61085), .B(n_30765), .C(n_300722032), .D(n_24716
		), .Z(n_299485408));
	notech_and4 i_141045086(.A(n_299485408), .B(n_299285406), .C(n_299185405
		), .D(n_285585269), .Z(n_299685410));
	notech_ao4 i_140245094(.A(n_381764348), .B(nbus_11273[8]), .C(n_381264343
		), .D(n_31481), .Z(n_299785411));
	notech_ao4 i_140145095(.A(n_5269), .B(n_381364344), .C(\nbus_11290[8] ),
		 .D(n_381664347), .Z(n_299885412));
	notech_ao4 i_139945097(.A(n_24527), .B(n_33548), .C(n_381464345), .D(n_33253
		), .Z(n_300085414));
	notech_and4 i_140445092(.A(n_300085414), .B(n_299885412), .C(n_299785411
		), .D(n_284885262), .Z(n_300285416));
	notech_ao4 i_110645353(.A(n_300822033), .B(n_388064411), .C(n_262470619)
		, .D(n_388164412), .Z(n_300385417));
	notech_ao4 i_110545354(.A(n_5243), .B(n_131626643), .C(n_131526642), .D(n_33206
		), .Z(n_300585419));
	notech_ao4 i_110245357(.A(n_387864409), .B(n_60458), .C(n_387964410), .D
		(n_58983), .Z(n_300785421));
	notech_and4 i_110445355(.A(n_300785421), .B(n_284085254), .C(n_30514), .D
		(n_283785251), .Z(n_301085424));
	notech_or2 i_41042880(.A(n_61816493), .B(n_4441), .Z(n_301185425));
	notech_or4 i_57442717(.A(n_28098), .B(n_26637), .C(n_61630), .D(n_59068)
		, .Z(n_301285426));
	notech_ao4 i_57642716(.A(n_324385655), .B(n_59068), .C(n_4440), .D(\nbus_11290[7] 
		), .Z(n_301385427));
	notech_or4 i_26643024(.A(n_28098), .B(n_340561033), .C(n_61621), .D(nbus_11271
		[1]), .Z(n_301985433));
	notech_or2 i_26143029(.A(n_60316478), .B(n_31482), .Z(n_302685440));
	notech_nand2 i_25243038(.A(add_src[9]), .B(n_30416), .Z(n_303585449));
	notech_or4 i_35242938(.A(n_28098), .B(n_340561033), .C(n_61611), .D(nbus_11271
		[6]), .Z(n_303685450));
	notech_or2 i_34742943(.A(n_60316478), .B(n_31487), .Z(n_304385457));
	notech_nand2 i_33842952(.A(add_src[14]), .B(n_30416), .Z(n_305285466));
	notech_or2 i_38342907(.A(n_60516480), .B(n_58357), .Z(n_305785471));
	notech_or4 i_38042910(.A(n_61890), .B(n_3964), .C(n_61711), .D(n_33160),
		 .Z(n_306085474));
	notech_nand2 i_39742893(.A(resb_shiftbox[17]), .B(n_30417), .Z(n_306585479
		));
	notech_nao3 i_39242898(.A(instrc[89]), .B(n_61702), .C(n_3964), .Z(n_307285486
		));
	notech_nand2 i_40942881(.A(resb_shiftbox[18]), .B(n_30417), .Z(n_307785491
		));
	notech_nao3 i_40442886(.A(instrc[90]), .B(n_61706), .C(n_3964), .Z(n_308485498
		));
	notech_or2 i_42042870(.A(n_60516480), .B(n_58384), .Z(n_309385507));
	notech_or4 i_41742873(.A(n_61890), .B(n_3964), .C(n_61717), .D(n_33138),
		 .Z(n_309685510));
	notech_or2 i_43242858(.A(n_60516480), .B(n_58393), .Z(n_310585519));
	notech_or4 i_42942861(.A(n_61890), .B(n_3964), .C(n_61711), .D(n_33163),
		 .Z(n_310885522));
	notech_or2 i_44442846(.A(n_60516480), .B(n_58402), .Z(n_311785531));
	notech_nao3 i_44142849(.A(instrc[93]), .B(n_61707), .C(n_3964), .Z(n_312085534
		));
	notech_or2 i_45642834(.A(n_60516480), .B(n_58411), .Z(n_312985543));
	notech_nao3 i_45342837(.A(instrc[94]), .B(n_61707), .C(n_3964), .Z(n_313285546
		));
	notech_or2 i_46842822(.A(n_60516480), .B(n_58420), .Z(n_314185555));
	notech_or4 i_46542825(.A(n_61878), .B(n_3964), .C(n_61711), .D(n_33141),
		 .Z(n_314485558));
	notech_or2 i_48042810(.A(n_60516480), .B(n_58429), .Z(n_315385567));
	notech_nao3 i_47742813(.A(instrc[96]), .B(n_61707), .C(n_3964), .Z(n_315785570
		));
	notech_or2 i_49242798(.A(n_60516480), .B(n_58438), .Z(n_316685579));
	notech_or4 i_48942801(.A(n_61878), .B(n_3964), .C(n_61711), .D(n_33159),
		 .Z(n_316985582));
	notech_or2 i_50442786(.A(n_60516480), .B(n_58447), .Z(n_317885591));
	notech_or4 i_50142789(.A(n_61880), .B(n_3964), .C(n_61717), .D(n_33178),
		 .Z(n_318185594));
	notech_or2 i_51642774(.A(n_60516480), .B(n_58456), .Z(n_319085603));
	notech_or4 i_51342777(.A(n_61878), .B(n_3964), .C(n_61717), .D(n_33139),
		 .Z(n_319385606));
	notech_or2 i_52842762(.A(n_56891), .B(n_58465), .Z(n_320385615));
	notech_or4 i_52542765(.A(n_61878), .B(n_3964), .C(n_61717), .D(n_33143),
		 .Z(n_320685618));
	notech_or2 i_55342738(.A(n_56891), .B(n_58483), .Z(n_321585627));
	notech_nao3 i_54942741(.A(instrc[102]), .B(n_61707), .C(n_3964), .Z(n_321885630
		));
	notech_or2 i_56642725(.A(n_56891), .B(n_60458), .Z(n_322785639));
	notech_or2 i_56342728(.A(n_61116486), .B(n_33142), .Z(n_323085642));
	notech_ao4 i_170941644(.A(n_61716492), .B(n_32256), .C(n_4438), .D(n_31539
		), .Z(n_323585647));
	notech_ao4 i_170841645(.A(n_323151206), .B(n_58983), .C(n_4436), .D(n_32345
		), .Z(n_323685648));
	notech_ao4 i_170641647(.A(n_60916484), .B(n_32240), .C(n_61016485), .D(n_60591
		), .Z(n_323885650));
	notech_and4 i_171141642(.A(n_323085642), .B(n_323885650), .C(n_323685648
		), .D(n_323585647), .Z(n_324085652));
	notech_ao4 i_170341650(.A(n_60216477), .B(n_5243), .C(n_60316478), .D(n_31507
		), .Z(n_324185653));
	notech_or4 i_171341641(.A(n_309960727), .B(n_339661024), .C(\opcode[0] )
		, .D(n_61824), .Z(n_324385655));
	notech_and2 i_72543300(.A(n_322951208), .B(n_301285426), .Z(n_324585657)
		);
	notech_and2 i_90343291(.A(n_324585657), .B(n_446968053), .Z(n_324685658)
		);
	notech_ao4 i_170141652(.A(n_4437), .B(n_32191), .C(n_59316468), .D(n_32734
		), .Z(n_324785659));
	notech_and4 i_170541648(.A(n_324685658), .B(n_324785659), .C(n_324185653
		), .D(n_322785639), .Z(n_324985661));
	notech_ao4 i_169841655(.A(n_61716492), .B(n_32298), .C(n_4438), .D(n_31538
		), .Z(n_325085662));
	notech_ao4 i_169741656(.A(n_323151206), .B(n_58992), .C(n_4436), .D(n_32344
		), .Z(n_325185663));
	notech_ao4 i_169541658(.A(n_60916484), .B(n_32239), .C(n_61016485), .D(n_60611
		), .Z(n_325385665));
	notech_and4 i_170041653(.A(n_321885630), .B(n_325385665), .C(n_325185663
		), .D(n_325085662), .Z(n_325585667));
	notech_ao4 i_169241661(.A(n_60216477), .B(n_5758), .C(n_60316478), .D(n_31506
		), .Z(n_325685668));
	notech_and2 i_191843271(.A(n_58016455), .B(n_324585657), .Z(n_325885670)
		);
	notech_ao4 i_169041663(.A(n_4437), .B(n_32190), .C(n_59316468), .D(n_32733
		), .Z(n_325985671));
	notech_and4 i_169441659(.A(n_325885670), .B(n_325985671), .C(n_325685668
		), .D(n_321585627), .Z(n_326185673));
	notech_ao4 i_167641677(.A(n_61716492), .B(n_32297), .C(n_4438), .D(n_31536
		), .Z(n_326285674));
	notech_ao4 i_167541678(.A(n_323151206), .B(n_58929), .C(n_4436), .D(n_32341
		), .Z(n_326385675));
	notech_ao4 i_167341680(.A(n_60916484), .B(n_32237), .C(n_61016485), .D(n_60564
		), .Z(n_326585677));
	notech_and4 i_167841675(.A(n_320685618), .B(n_326585677), .C(n_326385675
		), .D(n_326285674), .Z(n_326785679));
	notech_ao4 i_167041683(.A(n_60216477), .B(n_4427), .C(n_60316478), .D(n_31504
		), .Z(n_326885680));
	notech_ao4 i_166841685(.A(n_4437), .B(n_32187), .C(n_59316468), .D(n_32731
		), .Z(n_327085682));
	notech_and4 i_167241681(.A(n_324685658), .B(n_327085682), .C(n_326885680
		), .D(n_320385615), .Z(n_327285684));
	notech_ao4 i_166441688(.A(n_61716492), .B(n_32296), .C(n_4438), .D(n_31535
		), .Z(n_327385685));
	notech_ao4 i_166341689(.A(n_323151206), .B(n_58938), .C(n_4436), .D(n_32340
		), .Z(n_327485686));
	notech_ao4 i_166141691(.A(n_60916484), .B(n_32236), .C(n_61016485), .D(n_60573
		), .Z(n_327685688));
	notech_and4 i_166741686(.A(n_319385606), .B(n_327685688), .C(n_327485686
		), .D(n_327385685), .Z(n_327885690));
	notech_ao4 i_165841694(.A(n_60216477), .B(n_5711), .C(n_60316478), .D(n_31503
		), .Z(n_327985691));
	notech_ao4 i_165641696(.A(n_4437), .B(n_32185), .C(n_59316468), .D(n_32730
		), .Z(n_328185693));
	notech_and4 i_166041692(.A(n_324685658), .B(n_328185693), .C(n_327985691
		), .D(n_319085603), .Z(n_328385695));
	notech_ao4 i_165341699(.A(n_61716492), .B(n_32295), .C(n_4438), .D(n_31534
		), .Z(n_328485696));
	notech_ao4 i_165241700(.A(n_323151206), .B(n_58911), .C(n_4436), .D(n_32339
		), .Z(n_328585697));
	notech_ao4 i_165041702(.A(n_60916484), .B(n_32234), .C(n_61016485), .D(n_60582
		), .Z(n_328785699));
	notech_and4 i_165541697(.A(n_318185594), .B(n_328785699), .C(n_328585697
		), .D(n_328485696), .Z(n_328985701));
	notech_ao4 i_164741705(.A(n_60216477), .B(n_5720), .C(n_60316478), .D(n_31502
		), .Z(n_329085702));
	notech_ao4 i_164541707(.A(n_4437), .B(n_32183), .C(n_59316468), .D(n_32729
		), .Z(n_329285704));
	notech_and4 i_164941703(.A(n_325885670), .B(n_329285704), .C(n_329085702
		), .D(n_317885591), .Z(n_329485706));
	notech_ao4 i_164141710(.A(n_61716492), .B(n_32294), .C(n_4438), .D(n_31533
		), .Z(n_329585707));
	notech_ao4 i_164041711(.A(n_323151206), .B(n_58920), .C(n_4436), .D(n_32338
		), .Z(n_329685708));
	notech_ao4 i_163841713(.A(n_60916484), .B(n_32233), .C(n_61016485), .D(n_60510
		), .Z(n_329885710));
	notech_and4 i_164441708(.A(n_316985582), .B(n_329885710), .C(n_329685708
		), .D(n_329585707), .Z(n_330085712));
	notech_ao4 i_163541716(.A(n_101026337), .B(n_60216477), .C(n_60316478), 
		.D(n_31501), .Z(n_330185713));
	notech_ao4 i_163341718(.A(n_4437), .B(n_32182), .C(n_59316468), .D(n_32728
		), .Z(n_330385715));
	notech_and4 i_163741714(.A(n_325885670), .B(n_330385715), .C(n_330185713
		), .D(n_316685579), .Z(n_330585717));
	notech_ao4 i_163041721(.A(n_61716492), .B(n_32293), .C(n_4438), .D(n_31532
		), .Z(n_330685718));
	notech_ao4 i_162941722(.A(n_323151206), .B(n_58893), .C(n_4436), .D(n_32337
		), .Z(n_330785719));
	notech_ao4 i_162741724(.A(n_60916484), .B(n_32232), .C(n_61016485), .D(n_60519
		), .Z(n_330985721));
	notech_and4 i_163241719(.A(n_315785570), .B(n_330985721), .C(n_330785719
		), .D(n_330685718), .Z(n_331185723));
	notech_ao4 i_162441727(.A(n_60216477), .B(n_106826395), .C(n_60316478), 
		.D(n_31500), .Z(n_331285724));
	notech_ao4 i_162241729(.A(n_4437), .B(n_32180), .C(n_59316468), .D(n_32727
		), .Z(n_331685726));
	notech_and4 i_162641725(.A(n_324685658), .B(n_331685726), .C(n_331285724
		), .D(n_315385567), .Z(n_331885728));
	notech_ao4 i_161941732(.A(n_61716492), .B(n_32291), .C(n_56841), .D(n_31531
		), .Z(n_331985729));
	notech_ao4 i_161841733(.A(n_323151206), .B(n_58902), .C(n_4436), .D(n_32336
		), .Z(n_332085730));
	notech_ao4 i_161541735(.A(n_60916484), .B(n_32231), .C(n_61016485), .D(n_60528
		), .Z(n_332285732));
	notech_and4 i_162141730(.A(n_314485558), .B(n_332285732), .C(n_332085730
		), .D(n_331985729), .Z(n_332485734));
	notech_ao4 i_161141738(.A(n_109226419), .B(n_60216477), .C(n_56914), .D(n_31499
		), .Z(n_332585735));
	notech_ao4 i_160941740(.A(n_4437), .B(n_32179), .C(n_56871), .D(n_32726)
		, .Z(n_332785737));
	notech_and4 i_161341736(.A(n_324685658), .B(n_332785737), .C(n_332585735
		), .D(n_314185555), .Z(n_332985739));
	notech_ao4 i_160641743(.A(n_56823), .B(n_32289), .C(n_56841), .D(n_31530
		), .Z(n_333085740));
	notech_ao4 i_160541744(.A(n_323151206), .B(n_58875), .C(n_4436), .D(n_32333
		), .Z(n_333185741));
	notech_ao4 i_160341746(.A(n_60916484), .B(n_32230), .C(n_61016485), .D(n_60537
		), .Z(n_333385743));
	notech_and4 i_160841741(.A(n_313285546), .B(n_333385743), .C(n_333185741
		), .D(n_333085740), .Z(n_333585745));
	notech_ao4 i_159841749(.A(n_59464), .B(n_60216477), .C(n_56914), .D(n_31496
		), .Z(n_333685746));
	notech_ao4 i_159641751(.A(n_56904), .B(n_32178), .C(n_56871), .D(n_32725
		), .Z(n_333885748));
	notech_and4 i_160241747(.A(n_333885748), .B(n_333685746), .C(n_325885670
		), .D(n_312985543), .Z(n_334085750));
	notech_ao4 i_159341754(.A(n_56823), .B(n_32287), .C(n_56841), .D(n_31529
		), .Z(n_334185751));
	notech_ao4 i_159241755(.A(n_323151206), .B(n_58884), .C(n_4436), .D(n_32332
		), .Z(n_334285752));
	notech_ao4 i_159041757(.A(n_56861), .B(n_32229), .C(n_61016485), .D(n_60546
		), .Z(n_334485754));
	notech_and4 i_159541752(.A(n_312085534), .B(n_334485754), .C(n_334285752
		), .D(n_334185751), .Z(n_334685756));
	notech_ao4 i_158741760(.A(n_59465), .B(n_60216477), .C(n_56914), .D(n_31494
		), .Z(n_334885757));
	notech_ao4 i_158541762(.A(n_56904), .B(n_32177), .C(n_56871), .D(n_32724
		), .Z(n_335085759));
	notech_and4 i_158941758(.A(n_325885670), .B(n_335085759), .C(n_334885757
		), .D(n_311785531), .Z(n_335285761));
	notech_ao4 i_158241765(.A(n_56823), .B(n_32286), .C(n_56841), .D(n_31528
		), .Z(n_335385762));
	notech_ao4 i_158141766(.A(n_323151206), .B(n_58857), .C(n_56832), .D(n_32331
		), .Z(n_335485763));
	notech_ao4 i_157941768(.A(n_56861), .B(n_32228), .C(n_56850), .D(n_60555
		), .Z(n_335685765));
	notech_and4 i_158441763(.A(n_310885522), .B(n_335685765), .C(n_335485763
		), .D(n_335385762), .Z(n_335885767));
	notech_ao4 i_157641771(.A(n_59466), .B(n_56880), .C(n_56914), .D(n_31493
		), .Z(n_335985768));
	notech_ao4 i_157441773(.A(n_56904), .B(n_32175), .C(n_56871), .D(n_32723
		), .Z(n_336185770));
	notech_and4 i_157841769(.A(n_324685658), .B(n_336185770), .C(n_335985768
		), .D(n_310585519), .Z(n_336385772));
	notech_ao4 i_157141776(.A(n_56823), .B(n_32285), .C(n_56841), .D(n_31527
		), .Z(n_336485773));
	notech_ao4 i_157041777(.A(n_323151206), .B(n_58866), .C(n_56832), .D(n_32330
		), .Z(n_336585774));
	notech_ao4 i_156841779(.A(n_56861), .B(n_32226), .C(n_56850), .D(n_60483
		), .Z(n_336785776));
	notech_and4 i_157341774(.A(n_309685510), .B(n_336785776), .C(n_336585774
		), .D(n_336485773), .Z(n_336985778));
	notech_ao4 i_156541782(.A(n_56880), .B(n_5356), .C(n_56914), .D(n_31492)
		, .Z(n_337085779));
	notech_ao4 i_156341784(.A(n_56904), .B(n_32174), .C(n_56871), .D(n_32722
		), .Z(n_337285781));
	notech_and4 i_156741780(.A(n_337285781), .B(n_337085779), .C(n_324685658
		), .D(n_309385507), .Z(n_337485783));
	notech_ao4 i_156041787(.A(n_56823), .B(n_32284), .C(n_56841), .D(n_31526
		), .Z(n_337585784));
	notech_ao4 i_155941788(.A(n_323151206), .B(n_59077), .C(n_56832), .D(n_32329
		), .Z(n_337685785));
	notech_ao4 i_155741790(.A(n_56861), .B(n_32225), .C(n_56850), .D(n_60492
		), .Z(n_337885787));
	notech_and4 i_156241785(.A(n_308485498), .B(n_337885787), .C(n_337685785
		), .D(n_337585784), .Z(n_338085789));
	notech_ao4 i_155441793(.A(n_56880), .B(n_5436), .C(n_56914), .D(n_31491)
		, .Z(n_338185790));
	notech_ao4 i_155341794(.A(n_56871), .B(n_32720), .C(n_56891), .D(n_58375
		), .Z(n_338285791));
	notech_and4 i_155241795(.A(n_301185425), .B(n_324585657), .C(n_4435), .D
		(n_307785491), .Z(n_338685795));
	notech_ao4 i_154841799(.A(n_56823), .B(n_32283), .C(n_56841), .D(n_31525
		), .Z(n_338885797));
	notech_ao4 i_154741800(.A(n_323151206), .B(n_59086), .C(n_56832), .D(n_32328
		), .Z(n_338985798));
	notech_ao4 i_154541802(.A(n_56861), .B(n_32222), .C(n_56850), .D(n_60501
		), .Z(n_339185800));
	notech_and4 i_155041797(.A(n_307285486), .B(n_339185800), .C(n_338985798
		), .D(n_338885797), .Z(n_339385802));
	notech_ao4 i_154241805(.A(n_56880), .B(n_5397), .C(n_31490), .D(n_56914)
		, .Z(n_339485803));
	notech_ao4 i_154141806(.A(n_56871), .B(n_32719), .C(n_56891), .D(n_58366
		), .Z(n_339585804));
	notech_and4 i_154041807(.A(n_324585657), .B(n_301185425), .C(n_306585479
		), .D(n_4435), .Z(n_339885807));
	notech_ao4 i_153641811(.A(n_56823), .B(n_32282), .C(n_56841), .D(n_31524
		), .Z(n_340085809));
	notech_ao4 i_153541812(.A(n_323151206), .B(n_59059), .C(n_56832), .D(n_32327
		), .Z(n_340185810));
	notech_ao4 i_153341814(.A(n_56861), .B(n_32221), .C(n_56850), .D(n_60474
		), .Z(n_340385812));
	notech_and4 i_153841809(.A(n_306085474), .B(n_340385812), .C(n_340185810
		), .D(n_340085809), .Z(n_340585814));
	notech_ao4 i_153041817(.A(n_56880), .B(n_5444), .C(n_56914), .D(n_31489)
		, .Z(n_340685815));
	notech_ao4 i_152841819(.A(n_56904), .B(n_32173), .C(n_59316468), .D(n_32718
		), .Z(n_340885817));
	notech_and4 i_153241815(.A(n_340885817), .B(n_324685658), .C(n_340685815
		), .D(n_305785471), .Z(n_341085819));
	notech_ao4 i_150041845(.A(n_56823), .B(n_32277), .C(n_56841), .D(n_31522
		), .Z(n_341185820));
	notech_ao4 i_149941846(.A(n_40616281), .B(n_32281), .C(n_443982453), .D(n_59041
		), .Z(n_341385822));
	notech_and3 i_150241843(.A(n_341185820), .B(n_341385822), .C(n_305285466
		), .Z(n_341485823));
	notech_ao4 i_149741848(.A(n_40116276), .B(n_32879), .C(n_40216277), .D(n_31506
		), .Z(n_341585824));
	notech_ao4 i_149641849(.A(n_56850), .B(nbus_11271[14]), .C(n_40316278), 
		.D(n_32717), .Z(n_341685825));
	notech_ao4 i_149241853(.A(n_61116486), .B(n_33148), .C(n_56861), .D(n_32214
		), .Z(n_341985828));
	notech_ao4 i_149141854(.A(n_56891), .B(n_58339), .C(n_56880), .D(n_97342414
		), .Z(n_342185830));
	notech_ao4 i_148941856(.A(n_56929), .B(n_58992), .C(n_56904), .D(n_32171
		), .Z(n_342385832));
	notech_and4 i_149041855(.A(n_382982260), .B(n_58016455), .C(n_342385832)
		, .D(n_303685450), .Z(n_342585834));
	notech_and4 i_149541850(.A(n_304385457), .B(n_341985828), .C(n_342185830
		), .D(n_342585834), .Z(n_342685835));
	notech_ao4 i_142041925(.A(n_56823), .B(n_32280), .C(n_56841), .D(n_31517
		), .Z(n_342785836));
	notech_ao4 i_141941926(.A(n_40616281), .B(n_32279), .C(n_443982453), .D(n_59032
		), .Z(n_342985838));
	notech_and3 i_142241923(.A(n_342785836), .B(n_342985838), .C(n_303585449
		), .Z(n_343085839));
	notech_ao4 i_141741928(.A(n_40116276), .B(n_32874), .C(n_40216277), .D(n_31501
		), .Z(n_343185840));
	notech_ao4 i_141641929(.A(n_56850), .B(nbus_11271[9]), .C(n_40316278), .D
		(n_32712), .Z(n_343285841));
	notech_ao4 i_141241933(.A(n_61116486), .B(n_33150), .C(n_56861), .D(n_32206
		), .Z(n_343585844));
	notech_ao4 i_141141934(.A(n_56891), .B(n_58294), .C(n_56880), .D(n_99942440
		), .Z(n_343785846));
	notech_ao4 i_140741936(.A(n_56929), .B(n_58920), .C(n_56904), .D(n_32166
		), .Z(n_343985848));
	notech_and4 i_140841935(.A(n_382982260), .B(n_58016455), .C(n_343985848)
		, .D(n_301985433), .Z(n_344185850));
	notech_and4 i_141541930(.A(n_343585844), .B(n_343785846), .C(n_344185850
		), .D(n_302685440), .Z(n_344285851));
	notech_ao3 i_5461(.A(n_61611), .B(n_56965), .C(n_19707), .Z(n_344385852)
		);
	notech_nao3 i_73637521(.A(n_61917), .B(n_61903), .C(n_301960648), .Z(n_344485853
		));
	notech_ao4 i_18937337(.A(n_347185880), .B(n_58784), .C(n_351885926), .D(n_348485892
		), .Z(n_344685855));
	notech_ao4 i_130537741(.A(n_345285861), .B(n_59100), .C(n_25682), .D(n_349285900
		), .Z(n_344785856));
	notech_and2 i_183937742(.A(n_349185899), .B(n_349085898), .Z(n_344885857
		));
	notech_nor2 i_62737736(.A(n_4424), .B(n_345385862), .Z(n_345285861));
	notech_and3 i_47837083(.A(n_19707), .B(n_349385901), .C(n_30712), .Z(n_345385862
		));
	notech_ao4 i_3437740(.A(n_58707), .B(n_2820), .C(n_32217), .D(n_30491), 
		.Z(n_345585864));
	notech_nand2 i_119237735(.A(n_58716), .B(n_340361031), .Z(n_345785866)
		);
	notech_nao3 i_25437285(.A(n_4592), .B(n_25665), .C(n_27924), .Z(n_346085869
		));
	notech_nao3 i_25137288(.A(n_4594), .B(n_61707), .C(n_4452), .Z(n_346385872
		));
	notech_nand2 i_24837291(.A(add_src[4]), .B(n_30492), .Z(n_346685875));
	notech_nao3 i_24437294(.A(nbus_143[4]), .B(n_27843), .C(n_4351), .Z(n_346985878
		));
	notech_or2 i_37305(.A(n_349285900), .B(n_2127), .Z(n_347085879));
	notech_or4 i_37289(.A(n_59114), .B(n_56965), .C(n_56956), .D(n_58802), .Z
		(n_347185880));
	notech_nao3 i_37277(.A(n_57112), .B(n_30360), .C(n_4425), .Z(n_348285890
		));
	notech_and3 i_167737588(.A(n_19707), .B(n_19698), .C(n_56965), .Z(n_348385891
		));
	notech_nao3 i_178737587(.A(n_56965), .B(n_56956), .C(n_344485853), .Z(n_348485892
		));
	notech_ao4 i_107736571(.A(n_345585864), .B(n_32300), .C(n_50409), .D(n_57097
		), .Z(n_348585893));
	notech_mux2 i_128937586(.S(opd[0]), .A(n_59114), .B(n_344485853), .Z(n_348685894
		));
	notech_mux2 i_107636572(.S(opd[1]), .A(n_59115), .B(n_344485853), .Z(n_348785895
		));
	notech_and2 i_153237585(.A(n_348785895), .B(n_348685894), .Z(n_348885896
		));
	notech_mux2 i_107536573(.S(opd[2]), .A(n_59114), .B(n_344485853), .Z(n_348985897
		));
	notech_and2 i_167037584(.A(n_348985897), .B(n_348885896), .Z(n_349085898
		));
	notech_mux2 i_107436574(.S(opd[3]), .A(n_59114), .B(n_344485853), .Z(n_349185899
		));
	notech_nand2 i_197937452(.A(n_19707), .B(n_30712), .Z(n_349285900));
	notech_and3 i_17580(.A(n_19672), .B(n_61611), .C(n_30636), .Z(n_349385901
		));
	notech_or4 i_188737589(.A(n_19707), .B(n_61707), .C(n_56965), .D(n_56956
		), .Z(n_349485902));
	notech_ao4 i_72736874(.A(n_347085879), .B(n_31512), .C(n_344685855), .D(opd
		[4]), .Z(n_349585903));
	notech_ao4 i_72536876(.A(n_33553), .B(n_345285861), .C(n_2129), .D(n_32885
		), .Z(n_349785905));
	notech_and4 i_73036872(.A(n_349785905), .B(n_349585903), .C(n_346685875)
		, .D(n_346985878), .Z(n_349985907));
	notech_ao4 i_72036879(.A(n_4353), .B(nbus_11271[4]), .C(n_56974), .D(n_344885857
		), .Z(n_350085908));
	notech_ao4 i_71536881(.A(n_4352), .B(nbus_11273[4]), .C(n_4350), .D(n_33552
		), .Z(n_350285910));
	notech_and4 i_72336877(.A(n_350285910), .B(n_350085908), .C(n_346385872)
		, .D(n_346085869), .Z(n_350485912));
	notech_and4 i_194771994(.A(n_128983745), .B(n_114683602), .C(n_113883594
		), .D(n_113583591), .Z(n_350585913101150));
	notech_and4 i_194871993(.A(n_129483750), .B(n_114683602), .C(n_129283748
		), .D(n_114283598), .Z(n_350685914101151));
	notech_and4 i_194671992(.A(n_129883754), .B(n_114683602), .C(n_129683752
		), .D(n_114783603), .Z(n_350785915101152));
	notech_nao3 i_193871991(.A(n_114983605), .B(n_114883604), .C(n_348285890
		), .Z(n_350885916));
	notech_or2 i_183071990(.A(n_115083606), .B(n_348285890), .Z(n_350985917)
		);
	notech_or2 i_183171989(.A(n_115183607), .B(n_348285890), .Z(n_351085918)
		);
	notech_or2 i_20771988(.A(n_115283608), .B(n_57024), .Z(n_351185919));
	notech_or2 i_12471984(.A(n_115483610), .B(n_57024), .Z(n_351285920));
	notech_or2 i_19271983(.A(n_115583611), .B(n_57024), .Z(n_351385921));
	notech_or2 i_19771982(.A(n_115683612), .B(n_57024), .Z(n_351485922));
	notech_or2 i_20071981(.A(n_115783613), .B(n_57024), .Z(n_351585923));
	notech_nor2 i_61471963(.A(n_4424), .B(n_349385901), .Z(n_351685924));
	notech_ao4 i_121471961(.A(n_19672), .B(n_61707), .C(n_351685924), .D(n_59095
		), .Z(n_351785925));
	notech_or4 i_37198(.A(n_61878), .B(n_27930), .C(n_61717), .D(n_30521), .Z
		(n_2128));
	notech_or4 i_37196(.A(n_61878), .B(n_27930), .C(n_61717), .D(n_27843), .Z
		(n_2129));
	notech_nand3 i_37201(.A(n_19672), .B(n_61611), .C(n_19645), .Z(n_2127)
		);
	notech_xor2 i_140943358(.A(n_31604), .B(opz[1]), .Z(n_57104));
	notech_and4 i_2520855(.A(n_151283968), .B(n_152483980), .C(n_443068014),
		 .D(n_152383979), .Z(n_19364));
	notech_or4 i_1521005(.A(n_30558), .B(n_150483960), .C(n_153083986), .D(n_30456
		), .Z(n_18608));
	notech_nand2 i_3121341(.A(n_154383999), .B(n_153883994), .Z(n_16054));
	notech_and4 i_1521325(.A(n_154984005), .B(n_154884004), .C(n_148583941),
		 .D(n_155284008), .Z(n_15958));
	notech_and4 i_221312(.A(n_156284018), .B(n_156184017), .C(n_156084016), 
		.D(n_156684022), .Z(n_15880));
	notech_nand2 i_1521773(.A(n_157584031), .B(n_158084036), .Z(n_15254));
	notech_nand2 i_221760(.A(n_159484050), .B(n_158784043), .Z(n_15176));
	notech_and4 i_2517591(.A(n_143783893), .B(n_159584051), .C(n_159784053),
		 .D(n_160284058), .Z(n_11710));
	notech_and3 i_48760680(.A(n_2742), .B(n_2745), .C(n_272363654), .Z(n_377364304
		));
	notech_or4 i_3120765(.A(n_170584161), .B(n_168284138), .C(n_170084156), 
		.D(n_30457), .Z(n_19748));
	notech_or4 i_3120861(.A(n_170584161), .B(n_167484130), .C(n_171584167), 
		.D(n_30459), .Z(n_19400));
	notech_or4 i_3120989(.A(n_170584161), .B(n_166684122), .C(n_172284174), 
		.D(n_30460), .Z(n_19052));
	notech_nand3 i_3121021(.A(n_173384183), .B(n_173284182), .C(n_173184181)
		, .Z(n_18704));
	notech_nand2 i_220992(.A(n_175484194), .B(n_174984189), .Z(n_18530));
	notech_or4 i_3121181(.A(n_170584161), .B(n_163984095), .C(n_175884198), 
		.D(n_30461), .Z(n_13520));
	notech_and4 i_121311(.A(n_163084086), .B(n_177984209), .C(n_177884208), 
		.D(n_178284212), .Z(n_15874));
	notech_and4 i_3117597(.A(n_178484214), .B(n_178684216), .C(n_162584081),
		 .D(n_179184221), .Z(n_11746));
	notech_nand2 i_27877(.A(n_63790), .B(opc_10[14]), .Z(n_377264303));
	notech_nand2 i_27858(.A(n_63788), .B(opc[14]), .Z(n_377164302));
	notech_or2 i_46560692(.A(n_385364384), .B(n_57553), .Z(n_377064301));
	notech_or2 i_86863394(.A(n_379364324), .B(n_379164322), .Z(n_376964300)
		);
	notech_and2 i_42960773(.A(n_382264353), .B(n_180884236), .Z(n_58051));
	notech_and4 i_112260764(.A(n_384864379), .B(n_384964380), .C(n_258463528
		), .D(n_116542606), .Z(n_57383));
	notech_and3 i_125260756(.A(n_385464385), .B(n_257363519), .C(n_180784235
		), .Z(n_57260));
	notech_nao3 i_87663393(.A(n_32259), .B(n_30658), .C(n_379164322), .Z(n_376864299
		));
	notech_nao3 i_13363226(.A(n_57696), .B(n_286063762), .C(n_94542386), .Z(n_376764298
		));
	notech_nao3 i_12863231(.A(n_57696), .B(n_286063762), .C(n_379164322), .Z
		(n_376664297));
	notech_nand2 i_201369259(.A(n_57407), .B(n_30662), .Z(n_287744312));
	notech_nand2 i_521827(.A(n_189184318), .B(n_188684313), .Z(n_12668));
	notech_nand2 i_3121917(.A(n_190084327), .B(n_189684323), .Z(n_12472));
	notech_and4 i_1521901(.A(n_190484331), .B(n_190684333), .C(n_191184338),
		 .D(n_185584282), .Z(n_12376));
	notech_and4 i_521891(.A(n_192084347), .B(n_191984346), .C(n_191884345), 
		.D(n_192484351), .Z(n_12316));
	notech_nand2 i_221888(.A(n_193784364), .B(n_193284359), .Z(n_12298));
	notech_nand2 i_121887(.A(n_194784374), .B(n_194384370), .Z(n_12292));
	notech_nand3 i_110660667(.A(n_258463528), .B(n_116542606), .C(n_384864379
		), .Z(n_244036119));
	notech_or2 i_163469276(.A(n_303744471), .B(n_332363895), .Z(n_28742));
	notech_nao3 i_159269277(.A(n_290663806), .B(n_33173), .C(n_3290), .Z(n_28741
		));
	notech_and4 i_46218(.A(n_4465), .B(n_364350916), .C(n_330281779), .D(n_214884568
		), .Z(n_7415));
	notech_nao3 i_156769281(.A(n_290663806), .B(n_33173), .C(n_303744471), .Z
		(n_28743));
	notech_or4 i_2920763(.A(n_216384583), .B(n_213584555), .C(n_215884578), 
		.D(n_30464), .Z(n_19736));
	notech_or4 i_2820762(.A(n_217484594), .B(n_212084543), .C(n_216984589), 
		.D(n_30465), .Z(n_19730));
	notech_or4 i_2720761(.A(n_30574), .B(n_211284535), .C(n_218084600), .D(n_30466
		), .Z(n_19724));
	notech_or4 i_2920859(.A(n_216384583), .B(n_210284527), .C(n_218784607), 
		.D(n_30467), .Z(n_19388));
	notech_or4 i_2820858(.A(n_217484594), .B(n_209484519), .C(n_219484614), 
		.D(n_30469), .Z(n_19382));
	notech_or4 i_2720857(.A(n_30574), .B(n_208684511), .C(n_220184621), .D(n_30470
		), .Z(n_19376));
	notech_or4 i_2920987(.A(n_216384583), .B(n_207884503), .C(n_220884628), 
		.D(n_30471), .Z(n_19040));
	notech_nand3 i_2921019(.A(n_221784637), .B(n_221684636), .C(n_221584635)
		, .Z(n_18692));
	notech_nand3 i_2721017(.A(n_222484644), .B(n_222384643), .C(n_222284642)
		, .Z(n_18680));
	notech_and4 i_120991(.A(n_205484479), .B(n_223084650), .C(n_327860906), 
		.D(n_222984649), .Z(n_18524));
	notech_or4 i_2921179(.A(n_216384583), .B(n_204684471), .C(n_223684656), 
		.D(n_30472), .Z(n_13508));
	notech_nand2 i_2921339(.A(n_224984669), .B(n_224484664), .Z(n_16042));
	notech_nand2 i_2821338(.A(n_225984679), .B(n_225484674), .Z(n_16036));
	notech_nand2 i_2721337(.A(n_226984689), .B(n_226484684), .Z(n_16030));
	notech_and4 i_2921915(.A(n_200284429), .B(n_227484694), .C(n_227684696),
		 .D(n_227384693), .Z(n_12460));
	notech_nand2 i_2821914(.A(n_228684706), .B(n_228284702), .Z(n_12454));
	notech_and4 i_2721913(.A(n_198484411), .B(n_229184711), .C(n_229384713),
		 .D(n_229084710), .Z(n_12448));
	notech_and4 i_2917595(.A(n_198084407), .B(n_229584715), .C(n_229784717),
		 .D(n_230284722), .Z(n_11734));
	notech_and4 i_2817594(.A(n_197184398), .B(n_230384723), .C(n_230584725),
		 .D(n_231084730), .Z(n_11728));
	notech_and4 i_2717593(.A(n_196284389), .B(n_231184731), .C(n_231384733),
		 .D(n_231884738), .Z(n_11722));
	notech_nand2 i_9155835(.A(read_data[27]), .B(n_61611), .Z(n_274331424)
		);
	notech_and3 i_182569288(.A(n_60152), .B(n_162462656), .C(n_287744312), .Z
		(n_288144316));
	notech_and3 i_105569293(.A(n_57544), .B(n_164562677), .C(n_165062682), .Z
		(n_288444319));
	notech_or2 i_95769295(.A(n_376564296), .B(n_32259), .Z(n_29681));
	notech_or2 i_95269296(.A(n_94542386), .B(n_32259), .Z(n_29680));
	notech_or2 i_95069297(.A(n_94542386), .B(n_57489), .Z(n_29678));
	notech_or2 i_13063229(.A(n_29891), .B(n_94542386), .Z(n_376564296));
	notech_or2 i_94169301(.A(n_376564296), .B(n_57489), .Z(n_29677));
	notech_or4 i_2020754(.A(n_261285029), .B(n_259285009), .C(n_260785024), 
		.D(n_30475), .Z(n_19682));
	notech_or4 i_1920753(.A(n_262385040), .B(n_258084997), .C(n_261885035), 
		.D(n_30476), .Z(n_19676));
	notech_or4 i_1820752(.A(n_263485051), .B(n_256884985), .C(n_262985046), 
		.D(n_30477), .Z(n_19670));
	notech_or4 i_1720751(.A(n_264585062), .B(n_255684973), .C(n_264085057), 
		.D(n_30478), .Z(n_19664));
	notech_or4 i_2020850(.A(n_261285029), .B(n_254884965), .C(n_265185068), 
		.D(n_30479), .Z(n_19334));
	notech_or4 i_1920849(.A(n_262385040), .B(n_254084957), .C(n_265985076), 
		.D(n_30480), .Z(n_19328));
	notech_or4 i_1820848(.A(n_263485051), .B(n_253284949), .C(n_266785084), 
		.D(n_30481), .Z(n_19322));
	notech_or4 i_1720847(.A(n_264585062), .B(n_252484941), .C(n_267585092), 
		.D(n_30482), .Z(n_19316));
	notech_nand2 i_420994(.A(n_269085107), .B(n_268485101), .Z(n_18542));
	notech_nand2 i_421058(.A(n_270285119), .B(n_269685113), .Z(n_16241));
	notech_nand2 i_2021330(.A(n_271385129), .B(n_270785124), .Z(n_15988));
	notech_nand2 i_1921329(.A(n_272585139), .B(n_271985134), .Z(n_15982));
	notech_nand2 i_1821328(.A(n_273585149), .B(n_273085144), .Z(n_15976));
	notech_nand2 i_1721327(.A(n_274585159), .B(n_274085154), .Z(n_15970));
	notech_nand2 i_421826(.A(n_275685170), .B(n_275185165), .Z(n_12662));
	notech_and4 i_2021906(.A(n_243084849), .B(n_276185175), .C(n_276385177),
		 .D(n_276085174), .Z(n_12406));
	notech_nand2 i_1921905(.A(n_277385187), .B(n_276985183), .Z(n_12400));
	notech_and4 i_1821904(.A(n_241184831), .B(n_277885192), .C(n_278085194),
		 .D(n_277785191), .Z(n_12394));
	notech_nand2 i_1721903(.A(n_279085204), .B(n_278685200), .Z(n_12388));
	notech_and4 i_421890(.A(n_279985213), .B(n_279885212), .C(n_279785211), 
		.D(n_280385217), .Z(n_12310));
	notech_and4 i_2017586(.A(n_280585219), .B(n_280785221), .C(n_238484804),
		 .D(n_281285226), .Z(n_11680));
	notech_and4 i_1917585(.A(n_281385227), .B(n_281585229), .C(n_237584795),
		 .D(n_282085234), .Z(n_11674));
	notech_or4 i_1817584(.A(n_282885242), .B(n_236684786), .C(n_30485), .D(n_30486
		), .Z(n_11668));
	notech_and4 i_1717583(.A(n_282985243), .B(n_283185245), .C(n_235784777),
		 .D(n_283685250), .Z(n_11662));
	notech_nand2 i_3249697(.A(read_data[16]), .B(n_61611), .Z(n_314525222)
		);
	notech_nand2 i_3449695(.A(read_data[18]), .B(n_61611), .Z(n_314325220)
		);
	notech_ao4 i_26769308(.A(n_30723), .B(n_32208), .C(n_57562), .D(n_57657)
		, .Z(n_26949));
	notech_or4 i_32736(.A(instrc[93]), .B(n_321960847), .C(instrc[95]), .D(n_30551
		), .Z(n_26662));
	notech_or4 i_32735(.A(instrc[89]), .B(instrc[91]), .C(n_30551), .D(n_30334
		), .Z(n_26663));
	notech_or2 i_147446504(.A(n_370464235), .B(n_3290), .Z(n_28855));
	notech_nao3 i_146746505(.A(n_32247), .B(n_30674), .C(n_3290), .Z(n_28860
		));
	notech_or2 i_10713(.A(n_288144316), .B(n_3131), .Z(n_301744451));
	notech_or4 i_10711(.A(n_32275), .B(n_2382), .C(n_3131), .D(n_162262654),
		 .Z(n_301844452));
	notech_or4 i_3220766(.A(n_293885352), .B(n_291885332), .C(n_293385347), 
		.D(n_30488), .Z(n_19754));
	notech_or4 i_3220862(.A(n_293885352), .B(n_291085324), .C(n_294485358), 
		.D(n_30489), .Z(n_19406));
	notech_nand2 i_3221342(.A(n_295785371), .B(n_295285366), .Z(n_16060));
	notech_nand2 i_921319(.A(n_296985383), .B(n_296385377), .Z(n_15922));
	notech_nand2 i_921767(.A(n_298285396), .B(n_297685390), .Z(n_15218));
	notech_and4 i_3221918(.A(n_286385277), .B(n_298785401), .C(n_298985403),
		 .D(n_298685400), .Z(n_12478));
	notech_nand2 i_916999(.A(n_300285416), .B(n_299685410), .Z(n_11983));
	notech_and4 i_3217598(.A(n_284585259), .B(n_300385417), .C(n_300585419),
		 .D(n_301085424), .Z(n_11752));
	notech_or4 i_149869324(.A(n_32275), .B(n_56792), .C(n_26949), .D(n_162262654
		), .Z(n_26942));
	notech_nand2 i_3216222(.A(n_324985661), .B(n_324085652), .Z(n_13803));
	notech_nand2 i_3116221(.A(n_326185673), .B(n_325585667), .Z(n_13797));
	notech_nand2 i_2916219(.A(n_327285684), .B(n_326785679), .Z(n_13785));
	notech_nand2 i_2816218(.A(n_328385695), .B(n_327885690), .Z(n_13779));
	notech_nand2 i_2716217(.A(n_329485706), .B(n_328985701), .Z(n_13773));
	notech_nand2 i_2616216(.A(n_330585717), .B(n_330085712), .Z(n_13767));
	notech_nand2 i_2516215(.A(n_331885728), .B(n_331185723), .Z(n_13761));
	notech_nand2 i_2416214(.A(n_332985739), .B(n_332485734), .Z(n_13755));
	notech_nand2 i_2316213(.A(n_334085750), .B(n_333585745), .Z(n_13749));
	notech_nand2 i_2216212(.A(n_335285761), .B(n_334685756), .Z(n_13743));
	notech_nand2 i_2116211(.A(n_336385772), .B(n_335885767), .Z(n_13737));
	notech_nand2 i_2016210(.A(n_337485783), .B(n_336985778), .Z(n_13731));
	notech_and4 i_1916209(.A(n_338285791), .B(n_338185790), .C(n_338685795),
		 .D(n_338085789), .Z(n_13725));
	notech_and4 i_1816208(.A(n_339585804), .B(n_339485803), .C(n_339885807),
		 .D(n_339385802), .Z(n_13719));
	notech_nand2 i_1716207(.A(n_341085819), .B(n_340585814), .Z(n_13713));
	notech_and4 i_1516205(.A(n_341685825), .B(n_341585824), .C(n_342685835),
		 .D(n_341485823), .Z(n_13701));
	notech_and4 i_1016200(.A(n_343285841), .B(n_343185840), .C(n_344285851),
		 .D(n_343085839), .Z(n_13671));
	notech_ao4 i_71043302(.A(n_25705), .B(n_25680), .C(n_29534), .D(n_28098)
		, .Z(n_323151206));
	notech_or4 i_9415(.A(n_61917), .B(n_61903), .C(n_61878), .D(n_301385427)
		, .Z(n_322951208));
	notech_or2 i_130069327(.A(n_288144316), .B(n_164562677), .Z(n_302744461)
		);
	notech_nand2 i_194037743(.A(n_348585893), .B(n_30494), .Z(\nbus_11309[4] 
		));
	notech_nand2 i_512899(.A(n_350485912), .B(n_349985907), .Z(n_21327));
	notech_or4 i_129769328(.A(n_32275), .B(n_56792), .C(n_164562677), .D(n_162262654
		), .Z(n_302844462));
	notech_nand2 i_35173(.A(n_58802), .B(n_58784), .Z(n_351885926));
	notech_and2 i_127369329(.A(n_233663333), .B(n_165262684), .Z(n_302944463
		));
	notech_and2 i_127269330(.A(n_3293), .B(n_233563332), .Z(n_303044464));
	notech_and3 i_111469337(.A(n_190662933), .B(n_3314), .C(n_116342604), .Z
		(n_303744471));
	notech_nand2 i_44669355(.A(n_28854), .B(n_164962681), .Z(n_305044484));
	notech_and2 i_43069360(.A(n_305644490), .B(n_164762679), .Z(n_305544489)
		);
	notech_or4 i_39669361(.A(n_61824), .B(n_30309), .C(n_57633), .D(n_57091)
		, .Z(n_305644490));
	notech_ao4 i_27769364(.A(n_57553), .B(n_32208), .C(n_57672), .D(n_57566)
		, .Z(n_26951));
	notech_ao3 i_11469369(.A(n_339961027), .B(instrc[116]), .C(instrc[119]),
		 .Z(n_26957));
	notech_ao4 i_81137606(.A(n_381864349), .B(n_26028), .C(n_372564256), .D(n_372864259
		), .Z(n_376464295));
	notech_and2 i_182360727(.A(n_273863669), .B(n_60152), .Z(n_376364294));
	notech_ao3 i_188260719(.A(instrc[120]), .B(n_30646), .C(n_32269), .Z(n_376264293
		));
	notech_and2 i_97158158(.A(n_60152), .B(n_286163763), .Z(n_376064291));
	notech_or2 i_29814(.A(instrc[102]), .B(n_30550), .Z(n_29584));
	notech_ao3 i_12260792(.A(n_273263663), .B(n_57696), .C(instrc[119]), .Z(n_26063
		));
	notech_nand3 i_30206(.A(n_33173), .B(n_286063762), .C(n_63780), .Z(n_375764288
		));
	notech_nand2 i_178137617(.A(n_33164), .B(instrc[104]), .Z(n_375664287)
		);
	notech_or4 i_29168(.A(n_371764248), .B(n_30618), .C(n_33157), .D(n_30343
		), .Z(n_375564286));
	notech_ao3 i_11358218(.A(n_30727), .B(n_33173), .C(instrc[118]), .Z(n_29214
		));
	notech_or4 i_29161(.A(instrc[93]), .B(n_321960847), .C(n_30551), .D(n_33141
		), .Z(n_375464285));
	notech_or4 i_29144(.A(instrc[89]), .B(n_30551), .C(n_30334), .D(n_33138)
		, .Z(n_375364284));
	notech_or4 i_196337453(.A(n_32484), .B(instrc[102]), .C(n_61707), .D(instrc
		[101]), .Z(n_375264283));
	notech_or4 i_201037448(.A(n_32484), .B(n_61707), .C(instrc[98]), .D(instrc
		[97]), .Z(n_375164282));
	notech_or4 i_6671898(.A(n_32484), .B(n_61707), .C(instrc[98]), .D(n_33159
		), .Z(n_29572));
	notech_and2 i_3171933(.A(instrc[125]), .B(n_33175), .Z(n_29582));
	notech_and4 i_92443367(.A(n_360964140), .B(n_360864139), .C(n_360464135)
		, .D(n_360764138), .Z(n_375064281));
	notech_nand2 i_1417996(.A(n_154662578), .B(n_154562577), .Z(write_data_26
		[13]));
	notech_nand2 i_1117993(.A(n_154462576), .B(n_154362575), .Z(write_data_26
		[10]));
	notech_nand2 i_518115(.A(n_153462566), .B(n_153362565), .Z(write_data_27
		[4]));
	notech_and4 i_86536761(.A(n_374364274), .B(n_374164272), .C(n_374064271)
		, .D(n_367464205), .Z(n_374564276));
	notech_ao4 i_86036766(.A(n_378664317), .B(\nbus_11290[13] ), .C(n_378764318
		), .D(nbus_11273[13]), .Z(n_374364274));
	notech_ao4 i_86236764(.A(n_378964320), .B(n_33213), .C(n_378864319), .D(n_375064281
		), .Z(n_374164272));
	notech_ao4 i_86336763(.A(n_378564316), .B(n_31475), .C(n_378464315), .D(n_31486
		), .Z(n_374064271));
	notech_and4 i_87236754(.A(n_373764268), .B(n_373664267), .C(n_373464265)
		, .D(n_373364264), .Z(n_373964270));
	notech_ao4 i_86636760(.A(n_55975), .B(n_32072), .C(n_55966), .D(n_33210)
		, .Z(n_373764268));
	notech_ao4 i_86736759(.A(n_331560943), .B(n_366164192), .C(n_55946), .D(n_31521
		), .Z(n_373664267));
	notech_ao4 i_86936757(.A(n_31498), .B(n_26397), .C(n_26396), .D(n_31495)
		, .Z(n_373464265));
	notech_ao4 i_87036756(.A(n_26394), .B(n_31497), .C(n_55955), .D(n_30993)
		, .Z(n_373364264));
	notech_ao4 i_124236424(.A(n_32249), .B(n_365964190), .C(n_60196), .D(n_30340
		), .Z(n_372964260));
	notech_or4 i_128236386(.A(n_389864429), .B(n_389764428), .C(opa[5]), .D(opa
		[2]), .Z(n_372864259));
	notech_or4 i_128636382(.A(opa[7]), .B(opa[6]), .C(n_27798), .D(n_372264253
		), .Z(n_372564256));
	notech_or4 i_128436384(.A(n_63716), .B(n_32573), .C(n_27835), .D(n_61938
		), .Z(n_372264253));
	notech_ao4 i_139236289(.A(n_111445606), .B(n_30363), .C(n_114845640), .D
		(n_57195), .Z(n_372064251));
	notech_ao4 i_139336288(.A(n_29917), .B(n_365864189), .C(n_370864239), .D
		(n_336063932), .Z(n_371864249));
	notech_nao3 i_140336278(.A(n_30829), .B(n_30869), .C(instrc[105]), .Z(n_371764248
		));
	notech_and4 i_140036281(.A(n_369764228), .B(n_371464245), .C(n_371064241
		), .D(n_370064231), .Z(n_371664247));
	notech_ao4 i_139636285(.A(n_375464285), .B(n_28572), .C(n_375364284), .D
		(n_28581), .Z(n_371464245));
	notech_ao4 i_139836283(.A(n_366964200), .B(n_366864199), .C(n_375264283)
		, .D(n_370664237), .Z(n_371064241));
	notech_and2 i_144837489(.A(n_116645658), .B(n_30798), .Z(n_370864239));
	notech_nao3 i_143436253(.A(n_33162), .B(n_63818), .C(n_370464235), .Z(n_370764238
		));
	notech_or4 i_143536252(.A(n_30618), .B(n_30343), .C(n_436667950), .D(n_33142
		), .Z(n_370664237));
	notech_and2 i_97046511(.A(n_346564003), .B(n_60152), .Z(n_370464235));
	notech_nand2 i_70936886(.A(n_57195), .B(n_57595), .Z(n_370364234));
	notech_nand3 i_70836887(.A(n_57595), .B(n_57195), .C(n_63782), .Z(n_370264233
		));
	notech_ao3 i_29825(.A(n_61609), .B(n_33178), .C(n_32484), .Z(n_370164232
		));
	notech_nao3 i_69736897(.A(n_290663806), .B(n_367064201), .C(n_57696), .Z
		(n_370064231));
	notech_or4 i_70136894(.A(instrc[98]), .B(instrc[97]), .C(n_4464), .D(n_30550
		), .Z(n_369764228));
	notech_or2 i_70436891(.A(n_375564286), .B(n_29232), .Z(n_369464225));
	notech_nao3 i_46337098(.A(n_57436), .B(n_30903), .C(n_26624), .Z(n_368764218
		));
	notech_or2 i_33001(.A(n_378564316), .B(n_30788), .Z(n_26397));
	notech_or2 i_33002(.A(n_338061008), .B(n_56003), .Z(n_26396));
	notech_or2 i_33004(.A(n_378564316), .B(n_56003), .Z(n_26394));
	notech_nand2 i_35637198(.A(sav_esp[13]), .B(n_61858), .Z(n_367464205));
	notech_nao3 i_8937409(.A(n_323060858), .B(n_370264233), .C(n_322960857),
		 .Z(n_367064201));
	notech_and4 i_9037408(.A(n_116645658), .B(n_30798), .C(n_339261020), .D(n_370364234
		), .Z(n_366964200));
	notech_ao4 i_8837410(.A(n_365864189), .B(n_370764238), .C(n_30363), .D(n_3298
		), .Z(n_366864199));
	notech_or4 i_48937072(.A(n_61824), .B(n_30309), .C(n_57657), .D(n_32342)
		, .Z(n_366264193));
	notech_and4 i_143646513(.A(n_346264000), .B(n_346163999), .C(n_345363995
		), .D(n_346063998), .Z(n_366164192));
	notech_ao4 i_124537500(.A(n_63770), .B(n_61959), .C(n_32397), .D(n_30340
		), .Z(n_365964190));
	notech_nao3 i_130437497(.A(n_33175), .B(instrc[127]), .C(instrc[125]), .Z
		(n_365864189));
	notech_ao4 i_24537550(.A(n_32342), .B(n_30721), .C(n_57562), .D(n_30698)
		, .Z(n_23759));
	notech_or2 i_150337763(.A(n_23760), .B(n_390364434), .Z(n_23747));
	notech_or4 i_149737765(.A(n_32275), .B(n_32250), .C(n_365964190), .D(n_23760
		), .Z(n_23750));
	notech_or4 i_29864(.A(n_61917), .B(n_61903), .C(n_61880), .D(n_340561033
		), .Z(n_29534));
	notech_and4 i_143141914(.A(n_353964071), .B(n_364864179), .C(n_365064181
		), .D(n_365464185), .Z(n_365564186));
	notech_and4 i_142641919(.A(n_382982260), .B(n_58016455), .C(n_365264183)
		, .D(n_353264064), .Z(n_365464185));
	notech_ao4 i_142541920(.A(n_56929), .B(n_58911), .C(n_56904), .D(n_32167
		), .Z(n_365264183));
	notech_ao4 i_142741918(.A(n_56891), .B(nbus_11273[10]), .C(n_353164063),
		 .D(n_56880), .Z(n_365064181));
	notech_ao4 i_142841917(.A(n_61116486), .B(n_33151), .C(n_56861), .D(n_32207
		), .Z(n_364864179));
	notech_ao4 i_143241913(.A(n_56850), .B(nbus_11271[10]), .C(n_40316278), 
		.D(n_32713), .Z(n_364564176));
	notech_ao4 i_143341912(.A(n_40116276), .B(n_32875), .C(n_40216277), .D(n_31502
		), .Z(n_364464175));
	notech_and3 i_143841907(.A(n_364064171), .B(n_364264173), .C(n_354864080
		), .Z(n_364364174));
	notech_ao4 i_143541910(.A(n_40616281), .B(n_32242), .C(n_443982453), .D(\nbus_11290[10] 
		), .Z(n_364264173));
	notech_ao4 i_143641909(.A(n_56823), .B(n_32245), .C(n_56841), .D(n_31518
		), .Z(n_364064171));
	notech_ao4 i_196741409(.A(n_58592), .B(n_32010), .C(n_58565), .D(n_31978
		), .Z(n_363764168));
	notech_ao4 i_196841408(.A(n_58570), .B(n_31422), .C(n_57524), .D(n_33207
		), .Z(n_363664167));
	notech_and2 i_197241404(.A(n_363464165), .B(n_363364164), .Z(n_363564166
		));
	notech_ao4 i_197041406(.A(n_57444), .B(n_31586), .C(n_57436), .D(n_31946
		), .Z(n_363464165));
	notech_ao4 i_197141405(.A(n_57412), .B(n_31913), .C(n_57407), .D(n_31881
		), .Z(n_363364164));
	notech_and4 i_198041396(.A(n_363064161), .B(n_362964160), .C(n_362764158
		), .D(n_362664157), .Z(n_363264163));
	notech_ao4 i_197441402(.A(n_57512), .B(n_31849), .C(n_58550), .D(n_31817
		), .Z(n_363064161));
	notech_ao4 i_197541401(.A(n_57500), .B(n_31785), .C(n_57489), .D(n_31753
		), .Z(n_362964160));
	notech_ao4 i_197741399(.A(n_57622), .B(n_33208), .C(n_30363), .D(n_31721
		), .Z(n_362764158));
	notech_ao4 i_197841398(.A(n_57467), .B(n_31689), .C(n_57456), .D(n_31657
		), .Z(n_362664157));
	notech_ao4 i_199541381(.A(n_58592), .B(n_32006), .C(n_58561), .D(n_31974
		), .Z(n_362364154));
	notech_ao4 i_199641380(.A(n_58570), .B(n_31418), .C(n_57524), .D(n_33108
		), .Z(n_362264153));
	notech_and2 i_200141376(.A(n_362064151), .B(n_361964150), .Z(n_362164152
		));
	notech_ao4 i_199941378(.A(n_57444), .B(n_31582), .C(n_57436), .D(n_31941
		), .Z(n_362064151));
	notech_ao4 i_200041377(.A(n_57412), .B(n_31909), .C(n_57407), .D(n_31877
		), .Z(n_361964150));
	notech_and4 i_200941368(.A(n_361664147), .B(n_361564146), .C(n_361364144
		), .D(n_361264143), .Z(n_361864149));
	notech_ao4 i_200341374(.A(n_57512), .B(n_31845), .C(n_58550), .D(n_31813
		), .Z(n_361664147));
	notech_ao4 i_200441373(.A(n_57500), .B(n_31781), .C(n_57489), .D(n_31749
		), .Z(n_361564146));
	notech_ao4 i_200641371(.A(n_57622), .B(n_33209), .C(n_30363), .D(n_31717
		), .Z(n_361364144));
	notech_ao4 i_200741370(.A(n_57467), .B(n_31685), .C(n_57456), .D(n_31653
		), .Z(n_361264143));
	notech_ao4 i_212841252(.A(n_58592), .B(n_32009), .C(n_58561), .D(n_31977
		), .Z(n_360964140));
	notech_ao4 i_212941251(.A(n_58570), .B(n_31421), .C(n_57524), .D(n_33212
		), .Z(n_360864139));
	notech_and2 i_213341247(.A(n_360664137), .B(n_360564136), .Z(n_360764138
		));
	notech_ao4 i_213141249(.A(n_57444), .B(n_31585), .C(n_57436), .D(n_31945
		), .Z(n_360664137));
	notech_ao4 i_213241248(.A(n_57412), .B(n_31912), .C(n_57406), .D(n_31880
		), .Z(n_360564136));
	notech_and4 i_214141239(.A(n_360264133), .B(n_360164132), .C(n_359964130
		), .D(n_359864129), .Z(n_360464135));
	notech_ao4 i_213541245(.A(n_57512), .B(n_31848), .C(n_58550), .D(n_31816
		), .Z(n_360264133));
	notech_ao4 i_213641244(.A(n_57500), .B(n_31784), .C(n_57489), .D(n_31752
		), .Z(n_360164132));
	notech_ao4 i_213841242(.A(n_57622), .B(n_33211), .C(n_57480), .D(n_31720
		), .Z(n_359964130));
	notech_ao4 i_213941241(.A(n_57467), .B(n_31688), .C(n_57456), .D(n_31656
		), .Z(n_359864129));
	notech_nand2 i_26943021(.A(add_src[10]), .B(n_30416), .Z(n_354864080));
	notech_or2 i_27843012(.A(n_56914), .B(n_31483), .Z(n_353964071));
	notech_or4 i_28343007(.A(n_28098), .B(n_340561033), .C(n_61609), .D(nbus_11271
		[2]), .Z(n_353264064));
	notech_and4 i_92143353(.A(n_362364154), .B(n_362264153), .C(n_361864149)
		, .D(n_362164152), .Z(n_353164063));
	notech_ao4 i_149945007(.A(n_302744461), .B(n_60458), .C(n_302844462), .D
		(n_58983), .Z(n_352864060));
	notech_nand3 i_150545002(.A(n_352464056), .B(n_352664058), .C(n_333163903
		), .Z(n_352764059));
	notech_ao4 i_150145005(.A(n_125426581), .B(n_5243), .C(n_125326580), .D(n_33206
		), .Z(n_352664058));
	notech_ao4 i_150345004(.A(n_387664407), .B(n_300822033), .C(n_387764408)
		, .D(n_262470619), .Z(n_352464056));
	notech_and4 i_181544698(.A(n_352164053), .B(n_351964051), .C(n_351864050
		), .D(n_333463906), .Z(n_352364055));
	notech_ao4 i_181044703(.A(n_57034), .B(n_33205), .C(n_310371085), .D(n_33204
		), .Z(n_352164053));
	notech_ao4 i_181244701(.A(n_310771089), .B(n_353164063), .C(n_61085), .D
		(n_30875), .Z(n_351964051));
	notech_ao4 i_181344700(.A(n_309871081), .B(n_3299), .C(n_30326), .D(n_30639
		), .Z(n_351864050));
	notech_and4 i_182144692(.A(n_351564047), .B(n_351364045), .C(n_351264044
		), .D(n_334163913), .Z(n_351764049));
	notech_ao4 i_181644697(.A(n_299422019), .B(n_336163933), .C(n_265570648)
		, .D(nbus_11273[10]), .Z(n_351564047));
	notech_ao4 i_181844695(.A(n_299222017), .B(\nbus_11290[10] ), .C(n_265370646
		), .D(n_336263934), .Z(n_351364045));
	notech_ao4 i_181944694(.A(n_265070645), .B(n_336363935), .C(n_264970644)
		, .D(n_336463936), .Z(n_351264044));
	notech_and4 i_185144662(.A(n_350964041), .B(n_350764039), .C(n_350664038
		), .D(n_334863920), .Z(n_351164043));
	notech_ao4 i_184644667(.A(n_57034), .B(n_33203), .C(n_310371085), .D(n_33213
		), .Z(n_350964041));
	notech_ao4 i_184844665(.A(n_310771089), .B(n_375064281), .C(n_61085), .D
		(n_30878), .Z(n_350764039));
	notech_ao4 i_184944664(.A(n_366164192), .B(n_309871081), .C(n_30326), .D
		(n_30638), .Z(n_350664038));
	notech_and4 i_185744656(.A(n_350364035), .B(n_350064033), .C(n_349964032
		), .D(n_335563927), .Z(n_350564037));
	notech_ao4 i_185244661(.A(n_31475), .B(n_299422019), .C(nbus_11273[13]),
		 .D(n_265570648), .Z(n_350364035));
	notech_ao4 i_185444659(.A(\nbus_11290[13] ), .B(n_299222017), .C(n_31495
		), .D(n_265370646), .Z(n_350064033));
	notech_ao4 i_185544658(.A(n_31497), .B(n_265070645), .C(n_31498), .D(n_264970644
		), .Z(n_349964032));
	notech_ao4 i_198444529(.A(n_57112), .B(n_31785), .C(n_57604), .D(n_33208
		), .Z(n_349464028));
	notech_ao4 i_198544528(.A(n_57130), .B(n_31753), .C(n_57147), .D(n_33207
		), .Z(n_349364027));
	notech_and2 i_198944524(.A(n_349164025), .B(n_349064024), .Z(n_349264026
		));
	notech_ao4 i_198744526(.A(n_57164), .B(n_31849), .C(n_57174), .D(n_32010
		), .Z(n_349164025));
	notech_ao4 i_198844525(.A(n_57195), .B(n_31721), .C(n_57199), .D(n_31946
		), .Z(n_349064024));
	notech_and4 i_199744516(.A(n_348764021), .B(n_348664020), .C(n_348364018
		), .D(n_348164017), .Z(n_348964023));
	notech_ao4 i_199144522(.A(n_57057), .B(n_31689), .C(n_57068), .D(n_31817
		), .Z(n_348764021));
	notech_ao4 i_199244521(.A(n_57091), .B(n_31881), .C(n_57097), .D(n_31586
		), .Z(n_348664020));
	notech_ao4 i_199444519(.A(n_58691), .B(n_31978), .C(n_59095), .D(n_31913
		), .Z(n_348364018));
	notech_ao4 i_199544518(.A(n_57211), .B(n_31422), .C(n_57230), .D(n_31657
		), .Z(n_348164017));
	notech_ao4 i_202144493(.A(n_57112), .B(n_31781), .C(n_57604), .D(n_33209
		), .Z(n_347764014));
	notech_ao4 i_202244492(.A(n_57130), .B(n_31749), .C(n_57152), .D(n_33108
		), .Z(n_347664013));
	notech_and2 i_202644488(.A(n_347464011), .B(n_347364010), .Z(n_347564012
		));
	notech_ao4 i_202444490(.A(n_57163), .B(n_31845), .C(n_57174), .D(n_32006
		), .Z(n_347464011));
	notech_ao4 i_202544489(.A(n_57195), .B(n_31717), .C(n_57199), .D(n_31941
		), .Z(n_347364010));
	notech_and4 i_203444480(.A(n_347064008), .B(n_346964007), .C(n_346764005
		), .D(n_346664004), .Z(n_347264009));
	notech_ao4 i_202844486(.A(n_57057), .B(n_31685), .C(n_57068), .D(n_31813
		), .Z(n_347064008));
	notech_ao4 i_202944485(.A(n_57091), .B(n_31877), .C(n_57097), .D(n_31582
		), .Z(n_346964007));
	notech_ao4 i_203144483(.A(n_58691), .B(n_31974), .C(n_59095), .D(n_31909
		), .Z(n_346764005));
	notech_ao4 i_203244482(.A(n_57211), .B(n_31418), .C(n_57230), .D(n_31653
		), .Z(n_346664004));
	notech_ao4 i_209544419(.A(n_60182), .B(n_332363895), .C(n_32247), .D(n_3298
		), .Z(n_346564003));
	notech_ao4 i_209644418(.A(n_57112), .B(n_31784), .C(n_57604), .D(n_33211
		), .Z(n_346264000));
	notech_ao4 i_209744417(.A(n_57130), .B(n_31752), .C(n_57152), .D(n_33212
		), .Z(n_346163999));
	notech_and2 i_210144413(.A(n_345963997), .B(n_345463996), .Z(n_346063998
		));
	notech_ao4 i_209944415(.A(n_57163), .B(n_31848), .C(n_57174), .D(n_32009
		), .Z(n_345963997));
	notech_ao4 i_210044414(.A(n_57195), .B(n_31720), .C(n_57199), .D(n_31945
		), .Z(n_345463996));
	notech_and4 i_210944405(.A(n_345063993), .B(n_344963992), .C(n_344663990
		), .D(n_344563989), .Z(n_345363995));
	notech_ao4 i_210344411(.A(n_57057), .B(n_31688), .C(n_57068), .D(n_31816
		), .Z(n_345063993));
	notech_ao4 i_210444410(.A(n_57091), .B(n_31880), .C(n_57097), .D(n_31585
		), .Z(n_344963992));
	notech_ao4 i_210644408(.A(n_58691), .B(n_31977), .C(n_59095), .D(n_31912
		), .Z(n_344663990));
	notech_ao4 i_210744407(.A(n_57211), .B(n_31421), .C(n_57225), .D(n_31656
		), .Z(n_344563989));
	notech_nao3 i_27900(.A(n_63794), .B(opa[13]), .C(n_63700), .Z(n_31498)
		);
	notech_nand2 i_27901(.A(n_63794), .B(opc[13]), .Z(n_31497));
	notech_nand2 i_27903(.A(n_63794), .B(opc_10[13]), .Z(n_31495));
	notech_nao3 i_27923(.A(n_61938), .B(opa[13]), .C(n_63712), .Z(n_31475)
		);
	notech_nao3 i_28032(.A(n_63770), .B(opa[10]), .C(n_63712), .Z(n_336463936
		));
	notech_nand2 i_28033(.A(n_63740), .B(opc[10]), .Z(n_336363935));
	notech_nand2 i_28035(.A(n_63740), .B(opc_10[10]), .Z(n_336263934));
	notech_nao3 i_28056(.A(n_61938), .B(opa[10]), .C(n_63712), .Z(n_336163933
		));
	notech_nand3 i_30530(.A(n_290663806), .B(n_57686), .C(n_63780), .Z(n_336063932
		));
	notech_nao3 i_30531(.A(n_332363895), .B(n_63780), .C(n_3292), .Z(n_28867
		));
	notech_or4 i_30546(.A(instrc[113]), .B(instrc[114]), .C(n_32217), .D(n_57256
		), .Z(n_28852));
	notech_or2 i_35784(.A(n_386364394), .B(n_30340), .Z(n_23614));
	notech_or2 i_35785(.A(n_386364394), .B(n_23763), .Z(n_23613));
	notech_or2 i_35787(.A(n_23760), .B(n_23763), .Z(n_23611));
	notech_nand2 i_81045629(.A(opd[13]), .B(n_300322028), .Z(n_335563927));
	notech_nao3 i_81745622(.A(n_19655), .B(read_data[13]), .C(n_60453), .Z(n_334863920
		));
	notech_nand2 i_76845671(.A(n_300322028), .B(opd[10]), .Z(n_334163913));
	notech_nao3 i_77545664(.A(n_19655), .B(read_data[10]), .C(n_60453), .Z(n_333463906
		));
	notech_nand3 i_45845972(.A(n_57392), .B(n_32208), .C(opd[31]), .Z(n_333163903
		));
	notech_nor2 i_46345967(.A(n_387564406), .B(n_60591), .Z(n_332463896));
	notech_and2 i_11546439(.A(n_290663806), .B(n_57686), .Z(n_332363895));
	notech_or4 i_105245406(.A(n_61824), .B(n_30309), .C(n_57657), .D(n_32216
		), .Z(n_3314));
	notech_nao3 i_105145407(.A(n_58561), .B(n_30635), .C(n_390464435), .Z(n_3312
		));
	notech_nand2 i_104945408(.A(n_115442595), .B(n_32342), .Z(n_3311));
	notech_or4 i_104245415(.A(n_61824), .B(n_30309), .C(n_30698), .D(n_32216
		), .Z(n_3310));
	notech_and4 i_88945565(.A(n_3290), .B(n_3310), .C(n_57544), .D(n_3291), 
		.Z(n_3300));
	notech_and4 i_143346446(.A(n_347764014), .B(n_347664013), .C(n_347264009
		), .D(n_347564012), .Z(n_3299));
	notech_and3 i_115249769(.A(n_301844452), .B(n_26942), .C(n_26940), .Z(n_125426581
		));
	notech_and3 i_115149770(.A(n_301744451), .B(n_3118), .C(n_26935), .Z(n_125326580
		));
	notech_nao3 i_136346412(.A(n_290663806), .B(n_57686), .C(n_3300), .Z(n_28869
		));
	notech_ao4 i_83446418(.A(n_63770), .B(n_61959), .C(n_332363895), .D(n_32397
		), .Z(n_3298));
	notech_ao4 i_24846426(.A(n_30721), .B(n_32216), .C(n_57562), .D(n_30698)
		, .Z(n_3297));
	notech_or4 i_39346434(.A(instrc[113]), .B(instrc[114]), .C(n_32217), .D(n_30316
		), .Z(n_28854));
	notech_nor2 i_12509(.A(n_370464235), .B(n_3297), .Z(n_3296));
	notech_or2 i_151146502(.A(n_370464235), .B(n_3291), .Z(n_3295));
	notech_nao3 i_12507(.A(n_32247), .B(n_30674), .C(n_3297), .Z(n_3294));
	notech_nao3 i_150246503(.A(n_32247), .B(n_30674), .C(n_3291), .Z(n_3293)
		);
	notech_nao3 i_129346435(.A(n_32247), .B(n_30674), .C(n_3292), .Z(n_28863
		));
	notech_ao4 i_25846506(.A(n_30316), .B(n_32216), .C(n_57562), .D(n_57633)
		, .Z(n_3292));
	notech_ao4 i_26846436(.A(n_30723), .B(n_32216), .C(n_57562), .D(n_57657)
		, .Z(n_3291));
	notech_ao4 i_27846437(.A(n_57553), .B(n_32216), .C(n_57672), .D(n_57562)
		, .Z(n_3290));
	notech_or2 i_130146438(.A(n_3292), .B(n_370464235), .Z(n_28874));
	notech_and4 i_147948314(.A(n_65022753), .B(n_3287), .C(n_3285), .D(n_3139
		), .Z(n_3289));
	notech_ao4 i_147548318(.A(n_33118), .B(n_3118), .C(n_26942), .D(n_338361011
		), .Z(n_3287));
	notech_ao4 i_147748316(.A(n_74522848), .B(n_3117), .C(n_185962886), .D(n_74622849
		), .Z(n_3285));
	notech_and4 i_148548308(.A(n_3281), .B(n_3278), .C(n_3277), .D(n_3142), 
		.Z(n_3284));
	notech_ao4 i_148048313(.A(n_75522858), .B(n_3115), .C(n_75622859), .D(n_3114
		), .Z(n_3281));
	notech_ao4 i_148248311(.A(n_75322856), .B(n_3113), .C(n_75222855), .D(n_3112
		), .Z(n_3278));
	notech_ao4 i_148348310(.A(n_74922852), .B(n_3111), .C(n_66222765), .D(n_57091
		), .Z(n_3277));
	notech_ao4 i_148748306(.A(n_302844462), .B(n_59059), .C(n_305644490), .D
		(n_31489), .Z(n_3274));
	notech_nand3 i_149248301(.A(n_3269), .B(n_3271), .C(n_3154), .Z(n_3273)
		);
	notech_ao4 i_148948304(.A(n_125326580), .B(n_33199), .C(n_125426581), .D
		(n_5444), .Z(n_3271));
	notech_ao4 i_149048303(.A(n_267385090), .B(n_57091), .C(n_387564406), .D
		(n_60474), .Z(n_3269));
	notech_ao4 i_149448299(.A(n_302844462), .B(n_59086), .C(n_305644490), .D
		(n_31490), .Z(n_3260));
	notech_nao3 i_149948294(.A(n_3251), .B(n_3257), .C(n_3163), .Z(n_3259)
		);
	notech_ao4 i_149648297(.A(n_125326580), .B(n_33200), .C(n_5397), .D(n_125426581
		), .Z(n_3257));
	notech_ao4 i_149748296(.A(n_57091), .B(n_266585082), .C(n_387564406), .D
		(n_60501), .Z(n_3251));
	notech_ao4 i_150148292(.A(n_302844462), .B(n_59077), .C(n_305644490), .D
		(n_31491), .Z(n_3248));
	notech_nao3 i_150648287(.A(n_3244), .B(n_3246), .C(n_3171), .Z(n_3247)
		);
	notech_ao4 i_150348290(.A(n_125326580), .B(n_33201), .C(n_125426581), .D
		(n_5436), .Z(n_3246));
	notech_ao4 i_150448289(.A(n_57091), .B(n_265785074), .C(n_387564406), .D
		(n_60492), .Z(n_3244));
	notech_ao4 i_150848285(.A(n_302844462), .B(n_58866), .C(n_305644490), .D
		(n_31492), .Z(n_3241));
	notech_nao3 i_151348280(.A(n_3235), .B(n_3238), .C(n_3180), .Z(n_3240)
		);
	notech_ao4 i_151048283(.A(n_125326580), .B(n_33202), .C(n_125426581), .D
		(n_5356), .Z(n_3238));
	notech_ao4 i_151148282(.A(n_57081), .B(n_305478064), .C(n_387564406), .D
		(n_60483), .Z(n_3235));
	notech_and4 i_166748126(.A(n_65022753), .B(n_3231), .C(n_3229), .D(n_3185
		), .Z(n_3233));
	notech_ao4 i_166348130(.A(n_33118), .B(n_3295), .C(n_338361011), .D(n_3293
		), .Z(n_3231));
	notech_ao4 i_166548128(.A(n_74522848), .B(n_3129), .C(n_177362801), .D(n_74622849
		), .Z(n_3229));
	notech_and4 i_167348120(.A(n_3223), .B(n_3221), .C(n_3218), .D(n_3188), 
		.Z(n_3226));
	notech_ao4 i_166848125(.A(n_75522858), .B(n_3126), .C(n_75622859), .D(n_3124
		), .Z(n_3223));
	notech_ao4 i_167048123(.A(n_75322856), .B(n_3123), .C(n_75222855), .D(n_3122
		), .Z(n_3221));
	notech_ao4 i_167148122(.A(n_74922852), .B(n_3119), .C(n_66222765), .D(n_57187
		), .Z(n_3218));
	notech_ao4 i_169648097(.A(n_28874), .B(n_58384), .C(n_28863), .D(n_58866
		), .Z(n_3214));
	notech_nand3 i_170148092(.A(n_3207), .B(n_3209), .C(n_3200), .Z(n_3210)
		);
	notech_ao4 i_169848095(.A(n_388264413), .B(n_5356), .C(n_388364414), .D(n_33202
		), .Z(n_3209));
	notech_ao4 i_169948094(.A(n_319725273), .B(n_28852), .C(n_28869), .D(n_232870324
		), .Z(n_3207));
	notech_nand2 i_35657(.A(n_63770), .B(n_30340), .Z(n_23741));
	notech_nao3 i_59649156(.A(n_57378), .B(opd[19]), .C(n_57187), .Z(n_3200)
		);
	notech_nor2 i_60149151(.A(n_28867), .B(n_60483), .Z(n_3193));
	notech_or4 i_56449188(.A(n_60188), .B(n_332363895), .C(n_177362801), .D(n_58256
		), .Z(n_3188));
	notech_or2 i_56749185(.A(n_178762815), .B(n_58784), .Z(n_3185));
	notech_ao3 i_36349380(.A(opc_10[19]), .B(n_63780), .C(n_387764408), .Z(n_3180
		));
	notech_nor2 i_36849375(.A(n_302744461), .B(n_58384), .Z(n_3172));
	notech_ao3 i_35049388(.A(opc_10[18]), .B(n_63780), .C(n_387764408), .Z(n_3171
		));
	notech_nor2 i_35949383(.A(n_302744461), .B(n_58375), .Z(n_3164));
	notech_ao3 i_33949396(.A(opc_10[17]), .B(n_63782), .C(n_387764408), .Z(n_3163
		));
	notech_nor2 i_34749391(.A(n_302744461), .B(n_58366), .Z(n_3155));
	notech_nao3 i_33049404(.A(opc_10[16]), .B(n_63778), .C(n_387764408), .Z(n_3154
		));
	notech_nor2 i_33549399(.A(n_302744461), .B(n_58357), .Z(n_3147));
	notech_or4 i_32249412(.A(n_60182), .B(n_26957), .C(n_185962886), .D(n_58256
		), .Z(n_3142));
	notech_nand2 i_32549409(.A(n_30665), .B(opd[3]), .Z(n_3139));
	notech_nao3 i_119648585(.A(n_63790), .B(n_30340), .C(n_391064441), .Z(n_3133
		));
	notech_and4 i_118748594(.A(n_366264193), .B(n_116342604), .C(n_23760), .D
		(n_23759), .Z(n_3132));
	notech_ao4 i_24769309(.A(n_30721), .B(n_32208), .C(n_57562), .D(n_30698)
		, .Z(n_3131));
	notech_and4 i_118148596(.A(n_165062682), .B(n_57544), .C(n_26949), .D(n_26951
		), .Z(n_3130));
	notech_nao3 i_153769284(.A(n_290663806), .B(n_57686), .C(n_3291), .Z(n_3129
		));
	notech_nor2 i_128769289(.A(n_332363895), .B(n_177362801), .Z(n_3127));
	notech_or4 i_169569269(.A(instrc[121]), .B(n_2577), .C(instrc[122]), .D(n_30707
		), .Z(n_3126));
	notech_or4 i_167669272(.A(instrc[121]), .B(n_2577), .C(n_177362801), .D(instrc
		[122]), .Z(n_3124));
	notech_or2 i_167269274(.A(n_177362801), .B(n_32247), .Z(n_3123));
	notech_nand2 i_172769266(.A(n_57476), .B(n_3127), .Z(n_3122));
	notech_nao3 i_156269282(.A(n_290663806), .B(n_57686), .C(n_177362801), .Z
		(n_3119));
	notech_or2 i_150969323(.A(n_288144316), .B(n_26949), .Z(n_3118));
	notech_nao3 i_154269283(.A(instrc[116]), .B(n_188662913), .C(n_26949), .Z
		(n_3117));
	notech_or2 i_128369290(.A(n_26957), .B(n_185962886), .Z(n_3116));
	notech_or4 i_174269263(.A(instrc[123]), .B(instrc[121]), .C(n_56792), .D
		(n_3116), .Z(n_3115));
	notech_or4 i_172369268(.A(instrc[123]), .B(instrc[121]), .C(n_56792), .D
		(n_185962886), .Z(n_3114));
	notech_or2 i_172669267(.A(n_185962886), .B(n_32272), .Z(n_3113));
	notech_or2 i_172869265(.A(n_3116), .B(n_32272), .Z(n_3112));
	notech_nao3 i_158669279(.A(instrc[116]), .B(n_188662913), .C(n_185962886
		), .Z(n_3111));
	notech_and4 i_212950965(.A(n_3106), .B(n_3105), .C(n_3103), .D(n_3040), 
		.Z(n_3108));
	notech_ao4 i_212650968(.A(n_131526642), .B(n_33288), .C(n_59465), .D(n_131626643
		), .Z(n_3106));
	notech_ao4 i_212550969(.A(n_387964410), .B(n_58884), .C(n_387864409), .D
		(n_58402), .Z(n_3105));
	notech_ao4 i_212450970(.A(n_131426641), .B(n_60546), .C(n_56035), .D(n_32549
		), .Z(n_3103));
	notech_and4 i_192951164(.A(n_3095), .B(n_3027), .C(n_3098), .D(n_3030), 
		.Z(n_3101));
	notech_and3 i_192551168(.A(n_375575066), .B(n_3096), .C(n_3026), .Z(n_3098
		));
	notech_ao4 i_192351170(.A(n_382264353), .B(n_31493), .C(n_56035), .D(n_32570
		), .Z(n_3096));
	notech_ao4 i_192751166(.A(n_59466), .B(n_365328693), .C(n_365528695), .D
		(n_58857), .Z(n_3095));
	notech_nand3 i_148551605(.A(n_3090), .B(n_3089), .C(n_3088), .Z(n_3092)
		);
	notech_ao4 i_148251608(.A(n_101026337), .B(n_125426581), .C(n_302844462)
		, .D(n_58920), .Z(n_3090));
	notech_ao4 i_148151609(.A(n_302744461), .B(n_58438), .C(n_387564406), .D
		(n_60510), .Z(n_3089));
	notech_ao4 i_148351607(.A(n_31501), .B(n_305644490), .C(n_125326580), .D
		(n_33172), .Z(n_3088));
	notech_and4 i_108751998(.A(n_3083), .B(n_3082), .C(n_3081), .D(n_74526072
		), .Z(n_3086));
	notech_ao4 i_108352002(.A(n_59466), .B(n_388264413), .C(n_28863), .D(n_58857
		), .Z(n_3083));
	notech_ao4 i_108252003(.A(n_28874), .B(n_58393), .C(n_28867), .D(n_60555
		), .Z(n_3082));
	notech_ao4 i_108452001(.A(n_28854), .B(n_31493), .C(n_388364414), .D(n_33292
		), .Z(n_3081));
	notech_nand3 i_107052015(.A(n_307663892), .B(n_3075), .C(n_3074), .Z(n_3078
		));
	notech_ao4 i_106752018(.A(n_59465), .B(n_388264413), .C(n_28863), .D(n_58884
		), .Z(n_307663892));
	notech_ao4 i_106652019(.A(n_28874), .B(n_58402), .C(n_28867), .D(n_60546
		), .Z(n_3075));
	notech_ao4 i_106852017(.A(n_28854), .B(n_31494), .C(n_388364414), .D(n_33288
		), .Z(n_3074));
	notech_and4 i_105552030(.A(n_3069), .B(n_3068), .C(n_3067), .D(n_354467708
		), .Z(n_3072));
	notech_ao4 i_105152034(.A(n_59464), .B(n_388264413), .C(n_28863), .D(n_58875
		), .Z(n_3069));
	notech_ao4 i_105052035(.A(n_28874), .B(n_58411), .C(n_28867), .D(n_60537
		), .Z(n_3068));
	notech_ao4 i_105252033(.A(n_28854), .B(n_31496), .C(n_388364414), .D(n_33284
		), .Z(n_3067));
	notech_nand3 i_103852047(.A(n_3062), .B(n_3061), .C(n_3060), .Z(n_3064)
		);
	notech_ao4 i_103552050(.A(n_109226419), .B(n_388264413), .C(n_28863), .D
		(n_58902), .Z(n_3062));
	notech_ao4 i_103452051(.A(n_28874), .B(n_58420), .C(n_28867), .D(n_60528
		), .Z(n_3061));
	notech_ao4 i_103652049(.A(n_28854), .B(n_31499), .C(n_388364414), .D(n_33170
		), .Z(n_3060));
	notech_nand2 i_102252063(.A(n_3056), .B(n_3055), .Z(n_3057));
	notech_ao4 i_102052065(.A(n_388364414), .B(n_33171), .C(n_106826395), .D
		(n_388264413), .Z(n_3056));
	notech_ao4 i_101952066(.A(n_28863), .B(n_58893), .C(n_28874), .D(n_58429
		), .Z(n_3055));
	notech_nao3 i_102152064(.A(n_443068014), .B(n_297063868), .C(n_297563873
		), .Z(n_3054));
	notech_nand3 i_100652079(.A(n_3048), .B(n_3047), .C(n_3046), .Z(n_3050)
		);
	notech_ao4 i_100352082(.A(n_101026337), .B(n_388264413), .C(n_28863), .D
		(n_58920), .Z(n_3048));
	notech_ao4 i_100252083(.A(n_28874), .B(n_58438), .C(n_28867), .D(n_60510
		), .Z(n_3047));
	notech_ao4 i_100452081(.A(n_31501), .B(n_28854), .C(n_388364414), .D(n_33172
		), .Z(n_3046));
	notech_or4 i_2217588(.A(n_75626083), .B(n_3041), .C(n_3033), .D(n_30708)
		, .Z(n_3042));
	notech_ao3 i_212350971(.A(opc_10[21]), .B(n_63782), .C(n_388164412), .Z(n_3041
		));
	notech_nao3 i_212150973(.A(n_57382), .B(opd[21]), .C(n_58691), .Z(n_3040
		));
	notech_nor2 i_212250972(.A(n_3466), .B(n_388064411), .Z(n_3033));
	notech_nand3 i_2121907(.A(n_3031), .B(n_3101), .C(n_3023), .Z(n_3032));
	notech_nao3 i_192051173(.A(opc_10[20]), .B(n_63778), .C(n_365428694), .Z
		(n_3031));
	notech_or2 i_191951174(.A(n_365228692), .B(n_33292), .Z(n_3030));
	notech_or2 i_191651177(.A(n_365628696), .B(n_58393), .Z(n_3027));
	notech_or2 i_192151172(.A(n_25110), .B(n_60555), .Z(n_3026));
	notech_or4 i_192251171(.A(n_58716), .B(n_58707), .C(n_57256), .D(n_346771358
		), .Z(n_3023));
	notech_or4 i_2621624(.A(n_353367697), .B(n_3092), .C(n_3021), .D(n_3014)
		, .Z(n_3022));
	notech_ao3 i_148051610(.A(n_63790), .B(opc_10[25]), .C(n_387764408), .Z(n_3021
		));
	notech_nor2 i_147951611(.A(n_363350926), .B(n_387664407), .Z(n_3014));
	notech_nand3 i_2121171(.A(n_3086), .B(n_3012), .C(n_3005), .Z(n_3013));
	notech_nao3 i_108152004(.A(opc_10[20]), .B(n_63756), .C(n_28869), .Z(n_3012
		));
	notech_or4 i_108052005(.A(n_340361031), .B(n_32217), .C(n_57256), .D(n_346771358
		), .Z(n_3005));
	notech_or4 i_2221172(.A(n_75626083), .B(n_3078), .C(n_3003), .D(n_2996),
		 .Z(n_3004));
	notech_ao3 i_106552020(.A(opc_10[21]), .B(n_63756), .C(n_28869), .Z(n_3003
		));
	notech_nor2 i_106452021(.A(n_3466), .B(n_28852), .Z(n_2996));
	notech_nand3 i_2321173(.A(n_3072), .B(n_2994), .C(n_298763885), .Z(n_2995
		));
	notech_nao3 i_104952036(.A(opc_10[22]), .B(n_63756), .C(n_28869), .Z(n_2994
		));
	notech_or4 i_104852037(.A(n_340361031), .B(n_32217), .C(n_57256), .D(n_3464
		), .Z(n_298763885));
	notech_or4 i_2421174(.A(n_77826105), .B(n_3064), .C(n_298563883), .D(n_297863876
		), .Z(n_298663884));
	notech_ao3 i_103352052(.A(n_63768), .B(opc_10[23]), .C(n_28869), .Z(n_298563883
		));
	notech_nor2 i_103252053(.A(n_363450925), .B(n_28852), .Z(n_297863876));
	notech_or4 i_2521175(.A(n_3057), .B(n_3054), .C(n_297663874), .D(n_296963867
		), .Z(n_297763875));
	notech_ao3 i_101752068(.A(n_63786), .B(opc_10[24]), .C(n_28869), .Z(n_297663874
		));
	notech_ao3 i_101552070(.A(n_57382), .B(opd[24]), .C(n_57187), .Z(n_297563873
		));
	notech_or2 i_101052075(.A(n_28867), .B(n_60519), .Z(n_297063868));
	notech_nor2 i_101652069(.A(n_364628688), .B(n_28852), .Z(n_296963867));
	notech_or4 i_2621176(.A(n_353367697), .B(n_3050), .C(n_296763865), .D(n_296063858
		), .Z(n_296863866));
	notech_ao3 i_100152084(.A(n_63786), .B(opc_10[25]), .C(n_28869), .Z(n_296763865
		));
	notech_nor2 i_100052085(.A(n_363350926), .B(n_28852), .Z(n_296063858));
	notech_and2 i_8753085(.A(n_63752), .B(n_25121), .Z(n_295963857));
	notech_ao4 i_120854782(.A(n_302744461), .B(n_58447), .C(n_302844462), .D
		(n_58911), .Z(n_295663854));
	notech_nand3 i_121354777(.A(n_295263850), .B(n_295463852), .C(n_287663777
		), .Z(n_295563853));
	notech_ao4 i_121054780(.A(n_125426581), .B(n_5720), .C(n_125326580), .D(n_33198
		), .Z(n_295463852));
	notech_ao4 i_121154779(.A(n_284231523), .B(n_387664407), .C(n_175169787)
		, .D(n_387764408), .Z(n_295263850));
	notech_ao4 i_121554775(.A(n_302744461), .B(n_58456), .C(n_302844462), .D
		(n_58938), .Z(n_294963847));
	notech_nand3 i_122054770(.A(n_294563843), .B(n_294763845), .C(n_288463785
		), .Z(n_294863846));
	notech_ao4 i_121754773(.A(n_125426581), .B(n_5711), .C(n_125326580), .D(n_33195
		), .Z(n_294763845));
	notech_ao4 i_121854772(.A(n_387664407), .B(n_284131522), .C(n_387764408)
		, .D(n_172669762), .Z(n_294563843));
	notech_ao4 i_122254768(.A(n_302744461), .B(n_58465), .C(n_302844462), .D
		(\nbus_11290[28] ), .Z(n_294263840));
	notech_nand3 i_122754763(.A(n_293863836), .B(n_294063838), .C(n_289263793
		), .Z(n_294163839));
	notech_ao4 i_122454766(.A(n_125426581), .B(n_4427), .C(n_125326580), .D(n_33196
		), .Z(n_294063838));
	notech_ao4 i_122554765(.A(n_387664407), .B(n_440082450), .C(n_387764408)
		, .D(n_7636), .Z(n_293863836));
	notech_ao4 i_122954761(.A(n_302744461), .B(n_58474), .C(n_302844462), .D
		(\nbus_11290[29] ), .Z(n_293563833));
	notech_and3 i_123454756(.A(n_293163829), .B(n_293363831), .C(n_290063800
		), .Z(n_293463832));
	notech_ao4 i_123154759(.A(n_125426581), .B(n_4428), .C(n_125326580), .D(n_33197
		), .Z(n_293363831));
	notech_ao4 i_123254758(.A(n_387664407), .B(n_4387), .C(n_387764408), .D(n_94229643
		), .Z(n_293163829));
	notech_ao3 i_51855921(.A(n_292863826), .B(n_293063828), .C(n_290463804),
		 .Z(n_65029351));
	notech_ao4 i_163154362(.A(n_30695), .B(n_58447), .C(n_31534), .D(n_61706
		), .Z(n_293063828));
	notech_ao4 i_163254361(.A(n_30689), .B(n_5720), .C(n_30697), .D(n_33198)
		, .Z(n_292863826));
	notech_or4 i_183354164(.A(opa[28]), .B(opa[29]), .C(opa[26]), .D(opa[27]
		), .Z(n_292663824));
	notech_or4 i_183654161(.A(opa[16]), .B(opa[17]), .C(opa[18]), .D(opa[19]
		), .Z(n_292363821));
	notech_or4 i_184054157(.A(opa[20]), .B(opa[21]), .C(opa[22]), .D(opa[23]
		), .Z(n_291963817));
	notech_or4 i_184354154(.A(opa[24]), .B(opa[25]), .C(opa[31]), .D(opa[30]
		), .Z(n_291663814));
	notech_nand2 i_184654151(.A(n_58312), .B(nbus_11273[10]), .Z(n_291163809
		));
	notech_or4 i_185054147(.A(opa[15]), .B(opa[12]), .C(opa[13]), .D(opa[14]
		), .Z(n_2910));
	notech_ao4 i_188154116(.A(n_286263764), .B(n_32244), .C(n_60182), .D(n_29557
		), .Z(n_290763807));
	notech_ao3 i_29840(.A(instrc[119]), .B(n_33152), .C(instrc[118]), .Z(n_290663806
		));
	notech_nand3 i_30064(.A(n_290663806), .B(n_57696), .C(n_30283), .Z(n_29334
		));
	notech_nao3 i_30065(.A(n_57696), .B(n_290663806), .C(n_378364314), .Z(n_29333
		));
	notech_nor2 i_78355184(.A(n_30693), .B(n_58911), .Z(n_290463804));
	notech_nand3 i_36455591(.A(n_57382), .B(n_32208), .C(opd[29]), .Z(n_290063800
		));
	notech_or2 i_36955586(.A(n_387564406), .B(n_60620), .Z(n_289363794));
	notech_nand3 i_35655599(.A(n_57382), .B(n_32208), .C(opd[28]), .Z(n_289263793
		));
	notech_nor2 i_36155594(.A(n_387564406), .B(n_60564), .Z(n_288563786));
	notech_nao3 i_34855607(.A(n_57382), .B(opd[27]), .C(n_57081), .Z(n_288463785
		));
	notech_nor2 i_35355602(.A(n_387564406), .B(n_60573), .Z(n_287763778));
	notech_nao3 i_34055615(.A(n_57382), .B(opd[26]), .C(n_57081), .Z(n_287663777
		));
	notech_nor2 i_34555610(.A(n_387564406), .B(n_60582), .Z(n_286963771));
	notech_or4 i_99854986(.A(n_61824), .B(n_30309), .C(n_30698), .D(n_32211)
		, .Z(n_286763769));
	notech_nand2 i_99154992(.A(n_32211), .B(n_115942600), .Z(n_286363765));
	notech_ao4 i_83655915(.A(n_63786), .B(n_61959), .C(n_32397), .D(n_29557)
		, .Z(n_286263764));
	notech_or4 i_53555917(.A(n_2910), .B(opa[8]), .C(opa[9]), .D(n_291163809
		), .Z(n_27835));
	notech_ao4 i_142556769(.A(n_32252), .B(n_285763759), .C(n_60182), .D(n_29214
		), .Z(n_286163763));
	notech_ao3 i_29506(.A(n_57714), .B(instrc[116]), .C(instrc[118]), .Z(n_286063762
		));
	notech_ao4 i_83558125(.A(n_63796), .B(n_61959), .C(n_32397), .D(n_29214)
		, .Z(n_285763759));
	notech_ao3 i_85259853(.A(n_259163535), .B(n_256363510), .C(n_335060978),
		 .Z(n_285563757));
	notech_ao4 i_85359852(.A(n_336463936), .B(n_23614), .C(n_336363935), .D(n_23613
		), .Z(n_285263754));
	notech_ao4 i_85459851(.A(n_336263934), .B(n_23611), .C(n_386364394), .D(n_336163933
		), .Z(n_285163753));
	notech_and4 i_86259843(.A(n_284863750), .B(n_284663748), .C(n_284563747)
		, .D(n_259863541), .Z(n_285063752));
	notech_ao4 i_85759848(.A(n_33204), .B(n_23747), .C(n_353164063), .D(n_23750
		), .Z(n_284863750));
	notech_ao4 i_85959846(.A(n_386164392), .B(\nbus_11290[10] ), .C(n_386064391
		), .D(nbus_11273[10]), .Z(n_284663748));
	notech_ao4 i_86059845(.A(n_56035), .B(n_32539), .C(n_58691), .D(n_256263509
		), .Z(n_284563747));
	notech_and3 i_108959626(.A(n_55802), .B(n_260363546), .C(n_256363510), .Z
		(n_284363745));
	notech_ao4 i_109059625(.A(n_336463936), .B(n_4533), .C(n_441768001), .D(nbus_11273
		[10]), .Z(n_284063742));
	notech_and4 i_109859617(.A(n_283763739), .B(n_283563737), .C(n_283463736
		), .D(n_2609), .Z(n_283963741));
	notech_ao4 i_109359622(.A(n_441668000), .B(\nbus_11290[10] ), .C(n_56035
		), .D(n_32562), .Z(n_283763739));
	notech_ao4 i_109559620(.A(n_57174), .B(n_256263509), .C(n_385464385), .D
		(n_336263934), .Z(n_283563737));
	notech_ao4 i_109659619(.A(n_33204), .B(n_385664387), .C(n_353164063), .D
		(n_385864389), .Z(n_283463736));
	notech_and3 i_112459594(.A(n_55802), .B(n_261463556), .C(n_30468), .Z(n_283263734
		));
	notech_ao4 i_112559593(.A(n_31498), .B(n_4533), .C(n_441768001), .D(nbus_11273
		[13]), .Z(n_282963731));
	notech_and4 i_113459585(.A(n_282663728), .B(n_282463726), .C(n_282363725
		), .D(n_262063562), .Z(n_282863730));
	notech_ao4 i_112959590(.A(\nbus_11290[13] ), .B(n_441668000), .C(n_56035
		), .D(n_32565), .Z(n_282663728));
	notech_ao4 i_113159588(.A(n_57174), .B(n_30474), .C(n_385464385), .D(n_31495
		), .Z(n_282463726));
	notech_ao4 i_113259587(.A(n_385664387), .B(n_33213), .C(n_375064281), .D
		(n_385864389), .Z(n_282363725));
	notech_nao3 i_125859475(.A(n_55802), .B(n_256363510), .C(n_262563566), .Z
		(n_282163723));
	notech_ao4 i_125959474(.A(n_336263934), .B(n_333978345), .C(n_336163933)
		, .D(n_57393), .Z(n_281863720));
	notech_and4 i_126859467(.A(n_281563717), .B(n_281363715), .C(n_263163572
		), .D(n_263463575), .Z(n_281763719));
	notech_ao4 i_126359471(.A(n_33204), .B(n_323978248), .C(n_353164063), .D
		(n_323778246), .Z(n_281563717));
	notech_ao4 i_126559469(.A(nbus_11273[10]), .B(n_57243), .C(n_57068), .D(n_256263509
		), .Z(n_281363715));
	notech_and4 i_134559395(.A(n_187576933), .B(n_281063712), .C(n_280863710
		), .D(n_263963580), .Z(n_281263714));
	notech_ao4 i_134159399(.A(n_3112), .B(n_31075), .C(n_3117), .D(n_31068),
		 .Z(n_281063712));
	notech_ao4 i_134359397(.A(n_3114), .B(n_31072), .C(n_3115), .D(n_31074),
		 .Z(n_280863710));
	notech_and4 i_135159389(.A(n_280563707), .B(n_280363705), .C(n_280263704
		), .D(n_264263583), .Z(n_280763709));
	notech_ao4 i_134659394(.A(n_31048), .B(n_3116), .C(n_185962886), .D(n_31047
		), .Z(n_280563707));
	notech_ao4 i_134859392(.A(n_56974), .B(n_305544489), .C(n_3118), .D(n_33104
		), .Z(n_280363705));
	notech_ao4 i_134959391(.A(n_26942), .B(n_334660974), .C(n_57081), .D(n_187176929
		), .Z(n_280263704));
	notech_and4 i_143859309(.A(n_187576933), .B(n_279963702), .C(n_279763700
		), .D(n_265163592), .Z(n_280163703));
	notech_ao4 i_143459313(.A(n_3122), .B(n_31075), .C(n_3129), .D(n_31068),
		 .Z(n_279963702));
	notech_ao4 i_143659311(.A(n_3124), .B(n_31072), .C(n_3126), .D(n_31074),
		 .Z(n_279763700));
	notech_and4 i_144459303(.A(n_2794), .B(n_279263696), .C(n_279163695), .D
		(n_265463595), .Z(n_279663699));
	notech_ao4 i_143959308(.A(n_31048), .B(n_30707), .C(n_177362801), .D(n_31047
		), .Z(n_2794));
	notech_ao4 i_144159306(.A(n_178762815), .B(n_56974), .C(n_3295), .D(n_33104
		), .Z(n_279263696));
	notech_ao4 i_144259305(.A(n_3293), .B(n_334660974), .C(n_57187), .D(n_187176929
		), .Z(n_279163695));
	notech_nand2 i_144759300(.A(n_278763691), .B(n_266463603), .Z(n_278863692
		));
	notech_ao4 i_144659301(.A(n_28741), .B(n_336263934), .C(n_336163933), .D
		(n_303744471), .Z(n_278763691));
	notech_and4 i_145359294(.A(n_278463688), .B(n_278263686), .C(n_266963606
		), .D(n_267263609), .Z(n_278663690));
	notech_ao4 i_144959298(.A(n_28855), .B(n_33204), .C(n_353164063), .D(n_28860
		), .Z(n_278463688));
	notech_ao4 i_145159296(.A(nbus_11273[10]), .B(n_302944463), .C(n_57187),
		 .D(n_256263509), .Z(n_278263686));
	notech_and4 i_147459276(.A(n_187576933), .B(n_277963683), .C(n_277763681
		), .D(n_277663680), .Z(n_278163685));
	notech_ao4 i_146759281(.A(n_31075), .B(n_29341), .C(n_29334), .D(n_31068
		), .Z(n_277963683));
	notech_ao4 i_147159279(.A(n_29333), .B(n_31067), .C(n_31072), .D(n_29338
		), .Z(n_277763681));
	notech_ao4 i_147259278(.A(n_29340), .B(n_31074), .C(n_31071), .D(n_29337
		), .Z(n_277663680));
	notech_and4 i_148259270(.A(n_277363677), .B(n_277163675), .C(n_277063674
		), .D(n_268163618), .Z(n_277563679));
	notech_ao4 i_147559275(.A(n_378364314), .B(n_31047), .C(n_386464395), .D
		(n_56974), .Z(n_277363677));
	notech_ao4 i_147959273(.A(n_29550), .B(n_33104), .C(n_29540), .D(n_334660974
		), .Z(n_277163675));
	notech_ao4 i_148059272(.A(n_29533), .B(\nbus_11290[4] ), .C(n_57057), .D
		(n_187176929), .Z(n_277063674));
	notech_nand2 i_148559267(.A(n_2766), .B(n_268963626), .Z(n_2767));
	notech_ao4 i_148459268(.A(n_336263934), .B(n_29416), .C(n_336163933), .D
		(n_445168035), .Z(n_2766));
	notech_and4 i_149259261(.A(n_2763), .B(n_2761), .C(n_269263629), .D(n_269563632
		), .Z(n_2765));
	notech_ao4 i_148759265(.A(n_33204), .B(n_57612), .C(n_353164063), .D(n_57611
		), .Z(n_2763));
	notech_ao4 i_148959263(.A(nbus_11273[10]), .B(n_445068034), .C(n_57057),
		 .D(n_256263509), .Z(n_2761));
	notech_nand2 i_152159236(.A(n_2757), .B(n_269963636), .Z(n_2758));
	notech_ao4 i_152059237(.A(n_336263934), .B(n_30078), .C(n_336163933), .D
		(n_72542166), .Z(n_2757));
	notech_and4 i_152759230(.A(n_2754), .B(n_2752), .C(n_270263639), .D(n_2706
		), .Z(n_2756));
	notech_ao4 i_152359234(.A(n_304744481), .B(n_33204), .C(n_353164063), .D
		(n_304644480), .Z(n_2754));
	notech_ao4 i_152559232(.A(n_72742168), .B(nbus_11273[10]), .C(n_57112), 
		.D(n_256263509), .Z(n_2752));
	notech_ao4 i_155959200(.A(n_353164063), .B(n_30503), .C(n_30496), .D(\nbus_11290[10] 
		), .Z(n_2751));
	notech_ao4 i_156059199(.A(n_30499), .B(nbus_11273[10]), .C(n_30501), .D(n_33204
		), .Z(n_2749));
	notech_ao4 i_156959191(.A(n_375064281), .B(n_30503), .C(n_30496), .D(\nbus_11290[13] 
		), .Z(n_2748));
	notech_ao4 i_157059190(.A(nbus_11273[13]), .B(n_30499), .C(n_30501), .D(n_33213
		), .Z(n_2746));
	notech_ao4 i_157259188(.A(n_97342414), .B(n_30503), .C(n_30496), .D(n_59041
		), .Z(n_2745));
	notech_ao4 i_157359187(.A(n_30499), .B(n_58339), .C(n_30501), .D(n_33215
		), .Z(n_2742));
	notech_ao4 i_159259168(.A(n_32263), .B(n_256563512), .C(n_60188), .D(n_26063
		), .Z(n_273863669));
	notech_ao4 i_159859162(.A(n_32241), .B(n_256763514), .C(n_60188), .D(n_30314
		), .Z(n_273763668));
	notech_or4 i_160159159(.A(n_61880), .B(n_57672), .C(n_61711), .D(n_61858
		), .Z(n_273463665));
	notech_or4 i_160259158(.A(n_61880), .B(n_61711), .C(n_61858), .D(n_1850)
		, .Z(n_273363664));
	notech_nor2 i_160659154(.A(n_57705), .B(n_33152), .Z(n_273263663));
	notech_ao4 i_162559135(.A(n_60163), .B(n_58601), .C(n_258963533), .D(n_25121
		), .Z(n_273063661));
	notech_nand2 i_6260578(.A(n_256863515), .B(n_57696), .Z(n_272763658));
	notech_nand3 i_38432(.A(n_290663806), .B(n_57696), .C(n_56002), .Z(n_20897
		));
	notech_nao3 i_77059935(.A(n_58574), .B(n_30647), .C(n_380864339), .Z(n_272463655
		));
	notech_or2 i_34856(.A(n_381564346), .B(n_30314), .Z(n_24542));
	notech_or2 i_34857(.A(n_381564346), .B(n_24736), .Z(n_24541));
	notech_or2 i_34859(.A(n_24733), .B(n_24736), .Z(n_24539));
	notech_or4 i_34870(.A(n_61859), .B(n_61706), .C(n_30524), .D(n_32451), .Z
		(n_24528));
	notech_or4 i_34871(.A(n_61859), .B(n_61706), .C(n_30524), .D(n_61286), .Z
		(n_24527));
	notech_nand2 i_75559950(.A(n_61609), .B(read_data[14]), .Z(n_272363654)
		);
	notech_nand2 i_75059955(.A(n_61609), .B(read_data[13]), .Z(n_271663649)
		);
	notech_nand2 i_73559970(.A(n_61609), .B(read_data[10]), .Z(n_271163644)
		);
	notech_or2 i_68560020(.A(n_4924), .B(\nbus_11290[10] ), .Z(n_2706));
	notech_or2 i_68860017(.A(n_4922), .B(n_31483), .Z(n_270263639));
	notech_nao3 i_69160014(.A(n_63796), .B(opc[10]), .C(n_30075), .Z(n_269963636
		));
	notech_ao3 i_69260013(.A(opa[10]), .B(n_30076), .C(n_60188), .Z(n_269663633
		));
	notech_or2 i_64960054(.A(n_444968033), .B(\nbus_11290[10] ), .Z(n_269563632
		));
	notech_or2 i_65260051(.A(n_445268036), .B(n_31483), .Z(n_269263629));
	notech_nao3 i_65560048(.A(n_63796), .B(opc[10]), .C(n_29418), .Z(n_268963626
		));
	notech_ao3 i_65660047(.A(opa[10]), .B(n_29417), .C(n_60188), .Z(n_268663623
		));
	notech_or4 i_64060063(.A(n_63706), .B(n_29342), .C(n_61938), .D(nbus_11273
		[4]), .Z(n_268163618));
	notech_nand2 i_61360090(.A(opb[10]), .B(n_30631), .Z(n_267263609));
	notech_nand2 i_61660087(.A(n_305044484), .B(opd[10]), .Z(n_266963606));
	notech_nao3 i_61960084(.A(n_63752), .B(opc[10]), .C(n_28743), .Z(n_266463603
		));
	notech_nor2 i_62060083(.A(n_28742), .B(n_336463936), .Z(n_266163600));
	notech_or4 i_60560098(.A(n_177362801), .B(n_60163), .C(n_32247), .D(nbus_11273
		[4]), .Z(n_265463595));
	notech_nao3 i_60860095(.A(n_63796), .B(opc[4]), .C(n_3119), .Z(n_265163592
		));
	notech_or2 i_52160179(.A(n_3113), .B(n_31071), .Z(n_264263583));
	notech_nao3 i_52460176(.A(n_63752), .B(opc[4]), .C(n_3111), .Z(n_263963580
		));
	notech_or2 i_50660193(.A(n_57244), .B(\nbus_11290[10] ), .Z(n_263463575)
		);
	notech_or2 i_51060190(.A(n_58030), .B(n_31483), .Z(n_263163572));
	notech_or4 i_17349(.A(n_301560644), .B(n_316160789), .C(n_2091), .D(n_33242
		), .Z(n_115087077));
	notech_and3 i_7571889(.A(n_57340), .B(n_57799), .C(n_56663), .Z(n_115187078
		));
	notech_nand2 i_7971885(.A(n_115387080), .B(n_62441), .Z(n_115287079));
	notech_or2 i_7671888(.A(n_30722), .B(n_124545737), .Z(n_115387080));
	notech_nand2 i_46872(.A(n_129187218), .B(n_115287079), .Z(n_8484));
	notech_ao4 i_47155(.A(n_348689368), .B(n_2178), .C(n_1835), .D(n_348889370
		), .Z(\nbus_11287[0] ));
	notech_or4 i_9371871(.A(n_61859), .B(n_61609), .C(n_33496), .D(n_364150918
		), .Z(n_115787084));
	notech_nand2 i_46754(.A(n_129287219), .B(n_115787084), .Z(\nbus_11280[0] 
		));
	notech_or4 i_34871632(.A(n_116587092), .B(n_61859), .C(n_61706), .D(n_30538
		), .Z(n_116187088));
	notech_or4 i_35171629(.A(n_61880), .B(n_48030), .C(n_61711), .D(n_61859)
		, .Z(n_116487091));
	notech_and4 i_54647(.A(n_119787124), .B(n_116487091), .C(n_129687223), .D
		(n_129587222), .Z(\nbus_11352[9] ));
	notech_ao4 i_2371941(.A(n_347971365), .B(n_186266289), .C(n_30524), .D(n_30936
		), .Z(n_116587092));
	notech_nand2 i_54648(.A(n_116187088), .B(n_30520), .Z(\nbus_11352[10] )
		);
	notech_nand2 i_54646(.A(n_119787124), .B(n_30950), .Z(\nbus_11352[8] )
		);
	notech_nand3 i_54645(.A(n_116187088), .B(n_129487221), .C(n_129987226), 
		.Z(\nbus_11352[6] ));
	notech_and3 i_36371617(.A(n_57657), .B(n_30698), .C(n_27843), .Z(n_116887095
		));
	notech_nand3 i_54644(.A(n_116187088), .B(n_129487221), .C(n_130087227), 
		.Z(\nbus_11352[2] ));
	notech_ao3 i_36871612(.A(n_30650), .B(n_30382), .C(n_186266289), .Z(n_117187098
		));
	notech_or4 i_54643(.A(n_117187098), .B(n_30722), .C(n_179566227), .D(n_251347005
		), .Z(\nbus_11352[1] ));
	notech_nao3 i_54642(.A(n_129487221), .B(n_116187088), .C(n_30670), .Z(\nbus_11352[0] 
		));
	notech_ao4 i_40971571(.A(n_130487231), .B(n_130387230), .C(n_30649), .D(n_348071366
		), .Z(n_117587102));
	notech_ao4 i_48504(.A(n_130587232), .B(n_33242), .C(n_61846), .D(n_117587102
		), .Z(\nbus_11301[0] ));
	notech_ao4 i_46567(.A(n_348689368), .B(n_4402), .C(n_239446886), .D(n_33496
		), .Z(\nbus_11277[0] ));
	notech_and4 i_43671544(.A(n_2112), .B(n_2111), .C(n_4452), .D(n_4467), .Z
		(n_117987106));
	notech_ao4 i_47694(.A(n_239346885), .B(n_130687233), .C(n_117987106), .D
		(n_348689368), .Z(\nbus_11289[16] ));
	notech_and4 i_44271538(.A(n_4330), .B(n_4345), .C(n_4458), .D(n_4452), .Z
		(n_118387110));
	notech_ao4 i_47692(.A(n_118387110), .B(n_348689368), .C(n_4468), .D(n_33496
		), .Z(\nbus_11289[5] ));
	notech_and3 i_47071510(.A(n_59515), .B(n_349171376), .C(n_118587112), .Z
		(n_118487111));
	notech_or4 i_5371911(.A(tss_esp0), .B(\opcode[0] ), .C(n_30321), .D(n_329571252
		), .Z(n_118587112));
	notech_nor2 i_47571505(.A(n_56867), .B(n_30672), .Z(n_118887115));
	notech_ao4 i_54918(.A(n_118887115), .B(n_33496), .C(n_348689368), .D(n_57099
		), .Z(\nbus_11354[0] ));
	notech_or4 i_54796(.A(n_2019), .B(n_30540), .C(n_131187238), .D(n_30539)
		, .Z(\nbus_11353[0] ));
	notech_nor2 i_48871492(.A(sema_rw), .B(n_57688), .Z(n_119387120));
	notech_or4 i_53091(.A(n_61859), .B(n_2019), .C(n_119387120), .D(n_30541)
		, .Z(n_18351));
	notech_and2 i_50171479(.A(write_ack), .B(n_30529), .Z(n_119487121));
	notech_ao4 i_49971481(.A(n_311371095), .B(n_30307), .C(n_331271269), .D(n_2081
		), .Z(n_119587122));
	notech_nand2 i_50071480(.A(n_83245324), .B(n_30672), .Z(n_119687123));
	notech_or4 i_47327(.A(n_336789252), .B(n_61859), .C(n_131787244), .D(n_119487121
		), .Z(n_9187));
	notech_or4 i_6071904(.A(n_49651676), .B(n_2152), .C(n_63818), .D(n_61824
		), .Z(n_119787124));
	notech_or4 i_50671474(.A(n_61880), .B(n_61711), .C(n_61859), .D(n_349571380
		), .Z(n_119887125));
	notech_nand3 i_47076(.A(n_119787124), .B(n_119887125), .C(n_3456), .Z(n_8737
		));
	notech_and2 i_56571415(.A(imm[16]), .B(n_32203), .Z(n_119987126));
	notech_and2 i_56771413(.A(imm[17]), .B(n_32203), .Z(n_120087127));
	notech_and2 i_56971411(.A(imm[18]), .B(n_32203), .Z(n_120187128));
	notech_and2 i_57171409(.A(imm[19]), .B(n_32203), .Z(n_120287129));
	notech_and2 i_57371407(.A(imm[20]), .B(n_32203), .Z(n_120387130));
	notech_and2 i_57571405(.A(imm[21]), .B(n_32203), .Z(n_120487131));
	notech_and2 i_57771403(.A(imm[25]), .B(n_32203), .Z(n_120587132));
	notech_and2 i_57971401(.A(imm[27]), .B(n_32203), .Z(n_120687133));
	notech_ao4 i_1915633(.A(n_249536174), .B(n_31526), .C(n_194891308), .D(n_31950
		), .Z(n_14427));
	notech_nand2 i_86271121(.A(divr_1[50]), .B(n_61614), .Z(n_120987136));
	notech_nand2 i_5127390(.A(n_132087247), .B(n_120987136), .Z(n_16752));
	notech_ao4 i_91171072(.A(n_4424), .B(n_384582276), .C(n_4347), .D(n_120687133
		), .Z(n_121287139));
	notech_nand2 i_2812922(.A(n_132787254), .B(n_30530), .Z(n_21442));
	notech_ao4 i_92871055(.A(n_4424), .B(n_384582276), .C(n_4347), .D(n_120587132
		), .Z(n_122187148));
	notech_nand2 i_2612920(.A(n_133487261), .B(n_30531), .Z(n_21432));
	notech_ao4 i_94571038(.A(n_4424), .B(n_384582276), .C(n_4347), .D(n_120487131
		), .Z(n_123087157));
	notech_nand2 i_2212916(.A(n_134187268), .B(n_30532), .Z(n_21412));
	notech_ao4 i_96271021(.A(n_4424), .B(n_384582276), .C(n_4347), .D(n_120387130
		), .Z(n_123987166));
	notech_nand2 i_2112915(.A(n_134887275), .B(n_30533), .Z(n_21407));
	notech_ao4 i_97971004(.A(n_56321), .B(n_384582276), .C(n_4347), .D(n_120287129
		), .Z(n_124887175));
	notech_nand2 i_2012914(.A(n_135587282), .B(n_30534), .Z(n_21402));
	notech_ao4 i_99670987(.A(n_56321), .B(n_384582276), .C(n_4347), .D(n_120187128
		), .Z(n_125787184));
	notech_or2 i_181771977(.A(n_120187128), .B(n_4347), .Z(\nbus_11309[18] )
		);
	notech_nand2 i_1912913(.A(n_136287289), .B(n_30535), .Z(n_21397));
	notech_ao4 i_101370970(.A(n_56321), .B(n_384582276), .C(n_4347), .D(n_120087127
		), .Z(n_126687193));
	notech_nand2 i_1812912(.A(n_136987296), .B(n_30536), .Z(n_21392));
	notech_ao4 i_103070953(.A(n_56321), .B(n_384582276), .C(n_4347), .D(n_119987126
		), .Z(n_127587202));
	notech_nand2 i_1712911(.A(n_137687303), .B(n_30537), .Z(n_21387));
	notech_or4 i_136770618(.A(n_61917), .B(n_61903), .C(n_61880), .D(n_128787214
		), .Z(n_128687213));
	notech_and3 i_2471940(.A(n_30560), .B(n_316471137), .C(n_335489239), .Z(n_128787214
		));
	notech_ao4 i_222665(.A(n_348789369), .B(n_137987306), .C(n_61706), .D(n_19629
		), .Z(n_7469));
	notech_ao4 i_8071884(.A(n_348689368), .B(n_115187078), .C(n_1835), .D(n_348889370
		), .Z(n_129187218));
	notech_ao4 i_9471870(.A(n_348889370), .B(n_30618), .C(n_56583), .D(n_33496
		), .Z(n_129287219));
	notech_ao4 i_35071630(.A(n_61846), .B(n_242146913), .C(n_250947001), .D(n_30804
		), .Z(n_129487221));
	notech_and2 i_77671962(.A(n_116187088), .B(n_129487221), .Z(n_129587222)
		);
	notech_or4 i_6471900(.A(n_61711), .B(n_61880), .C(n_240546897), .D(n_61861
		), .Z(n_129687223));
	notech_mux2 i_36171619(.S(n_4450), .A(n_57041), .B(n_129687223), .Z(n_129987226
		));
	notech_ao4 i_36671614(.A(n_116887095), .B(n_57041), .C(n_57047), .D(n_129687223
		), .Z(n_130087227));
	notech_nao3 i_41271568(.A(n_63728), .B(n_63712), .C(n_61797), .Z(n_130387230
		));
	notech_nand2 i_41371567(.A(n_32646), .B(n_63800), .Z(n_130487231));
	notech_or4 i_41671564(.A(n_57006), .B(n_30304), .C(n_61880), .D(n_31069)
		, .Z(n_130587232));
	notech_nand3 i_43971541(.A(n_61085), .B(n_61611), .C(n_62441), .Z(n_130687233
		));
	notech_ao4 i_48371497(.A(n_30681), .B(n_339489279), .C(n_57016), .D(n_33242
		), .Z(n_130987236));
	notech_nand2 i_48271498(.A(n_2130), .B(n_57717), .Z(n_131187238));
	notech_ao4 i_49071490(.A(n_83245324), .B(n_57717), .C(n_57681), .D(n_33242
		), .Z(n_131387240));
	notech_nand2 i_50371477(.A(n_2130), .B(n_119687123), .Z(n_131787244));
	notech_ao4 i_86371120(.A(n_24216), .B(n_33554), .C(n_56411), .D(n_60492)
		, .Z(n_132087247));
	notech_ao4 i_91271071(.A(n_4349), .B(n_33555), .C(n_112042561), .D(n_32340
		), .Z(n_132187248));
	notech_ao4 i_91371070(.A(n_24142), .B(n_33557), .C(n_4350), .D(n_33556),
		 .Z(n_132287249));
	notech_ao4 i_91471069(.A(n_4353), .B(n_60573), .C(n_4351), .D(n_32908), 
		.Z(n_132487251));
	notech_ao4 i_91571068(.A(n_4348), .B(n_31535), .C(n_4352), .D(n_58456), 
		.Z(n_132587252));
	notech_and4 i_91871065(.A(n_132587252), .B(n_132487251), .C(n_132287249)
		, .D(n_132187248), .Z(n_132787254));
	notech_ao4 i_92971054(.A(n_4349), .B(n_33558), .C(n_112042561), .D(n_32338
		), .Z(n_132887255));
	notech_ao4 i_93071053(.A(n_24142), .B(n_33560), .C(n_4350), .D(n_33559),
		 .Z(n_132987256));
	notech_ao4 i_93171052(.A(n_4353), .B(n_60510), .C(n_4351), .D(n_32906), 
		.Z(n_133187258));
	notech_ao4 i_93271051(.A(n_4348), .B(n_31533), .C(n_4352), .D(n_58438), 
		.Z(n_133287259));
	notech_and4 i_93571048(.A(n_133287259), .B(n_133187258), .C(n_132987256)
		, .D(n_132887255), .Z(n_133487261));
	notech_ao4 i_94671037(.A(n_4349), .B(n_33561), .C(n_112042561), .D(n_32332
		), .Z(n_133587262));
	notech_ao4 i_94771036(.A(n_4350), .B(n_33562), .C(n_4353), .D(n_60546), 
		.Z(n_133687263));
	notech_ao4 i_94871035(.A(n_4351), .B(n_32902), .C(n_56718), .D(n_33563),
		 .Z(n_133887265));
	notech_ao4 i_94971034(.A(n_4348), .B(n_31529), .C(n_4352), .D(n_58402), 
		.Z(n_133987266));
	notech_and4 i_95271031(.A(n_133987266), .B(n_133887265), .C(n_133687263)
		, .D(n_133587262), .Z(n_134187268));
	notech_ao4 i_96371020(.A(n_4349), .B(n_33564), .C(n_112042561), .D(n_32331
		), .Z(n_134287269));
	notech_ao4 i_96471019(.A(n_56718), .B(n_33566), .C(n_56341), .D(n_33565)
		, .Z(n_134387270));
	notech_ao4 i_96571018(.A(n_56359), .B(n_60555), .C(n_4351), .D(n_32901),
		 .Z(n_134587272));
	notech_ao4 i_96671017(.A(n_4348), .B(n_31528), .C(n_56350), .D(n_58393),
		 .Z(n_134687273));
	notech_and4 i_96971014(.A(n_134687273), .B(n_134587272), .C(n_134387270)
		, .D(n_134287269), .Z(n_134887275));
	notech_ao4 i_98071003(.A(n_56330), .B(n_33567), .C(n_112042561), .D(n_32330
		), .Z(n_134987276));
	notech_ao4 i_98171002(.A(n_56718), .B(n_33569), .C(n_56341), .D(n_33568)
		, .Z(n_135087277));
	notech_ao4 i_98271001(.A(n_56359), .B(n_60483), .C(n_4351), .D(n_32900),
		 .Z(n_135287279));
	notech_ao4 i_98371000(.A(n_4348), .B(n_31527), .C(n_56350), .D(n_58384),
		 .Z(n_135387280));
	notech_and4 i_98670997(.A(n_135387280), .B(n_135287279), .C(n_135087277)
		, .D(n_134987276), .Z(n_135587282));
	notech_ao4 i_99770986(.A(n_56330), .B(n_33570), .C(n_112042561), .D(n_32329
		), .Z(n_135687283));
	notech_ao4 i_99870985(.A(n_56718), .B(n_33572), .C(n_56341), .D(n_33571)
		, .Z(n_135787284));
	notech_ao4 i_99970984(.A(n_56359), .B(n_60492), .C(n_4351), .D(n_32899),
		 .Z(n_135987286));
	notech_ao4 i_100070983(.A(n_4348), .B(n_31526), .C(n_56350), .D(n_58375)
		, .Z(n_136087287));
	notech_and4 i_100370980(.A(n_136087287), .B(n_135987286), .C(n_135787284
		), .D(n_135687283), .Z(n_136287289));
	notech_ao4 i_101470969(.A(n_56330), .B(n_33573), .C(n_112042561), .D(n_32328
		), .Z(n_136387290));
	notech_ao4 i_101570968(.A(n_56718), .B(n_33575), .C(n_56341), .D(n_33574
		), .Z(n_136487291));
	notech_ao4 i_101670967(.A(n_56359), .B(n_60501), .C(n_4351), .D(n_32898)
		, .Z(n_136687293));
	notech_ao4 i_101770966(.A(n_4348), .B(n_31525), .C(n_56350), .D(n_58366)
		, .Z(n_136787294));
	notech_and4 i_102070963(.A(n_136787294), .B(n_136687293), .C(n_136487291
		), .D(n_136387290), .Z(n_136987296));
	notech_ao4 i_103170952(.A(n_56330), .B(n_33576), .C(n_112042561), .D(n_32327
		), .Z(n_137087297));
	notech_ao4 i_103270951(.A(n_56718), .B(n_33578), .C(n_56341), .D(n_33577
		), .Z(n_137187298));
	notech_ao4 i_103370950(.A(n_56359), .B(n_60474), .C(n_4351), .D(n_32897)
		, .Z(n_137387300));
	notech_ao4 i_103470949(.A(n_4348), .B(n_31524), .C(n_56350), .D(n_58357)
		, .Z(n_137487301));
	notech_and4 i_103770946(.A(n_137487301), .B(n_137387300), .C(n_137187298
		), .D(n_137087297), .Z(n_137687303));
	notech_mux2 i_2171943(.S(n_61707), .A(n_19629), .B(n_30627), .Z(n_137787304
		));
	notech_nand2 i_137070615(.A(calc_sz[2]), .B(n_57657), .Z(n_137987306));
	notech_and2 i_14669119(.A(imm[22]), .B(n_32203), .Z(n_138087307));
	notech_and2 i_14869117(.A(imm[23]), .B(n_32203), .Z(n_138187308));
	notech_and2 i_15069115(.A(imm[24]), .B(n_32203), .Z(n_138287309));
	notech_and2 i_15269113(.A(imm[26]), .B(n_57236), .Z(n_138387310));
	notech_and2 i_15469111(.A(imm[28]), .B(n_57236), .Z(n_138487311));
	notech_nao3 i_161167739(.A(n_3516), .B(n_60607), .C(n_56428), .Z(n_138587312
		));
	notech_nand2 i_2927368(.A(n_144587372), .B(n_138587312), .Z(n_16642));
	notech_nao3 i_162167729(.A(n_3514), .B(n_60605), .C(n_56428), .Z(n_138887315
		));
	notech_nand2 i_2727366(.A(n_144687373), .B(n_138887315), .Z(n_16632));
	notech_nao3 i_163167719(.A(n_3512), .B(n_60605), .C(n_56428), .Z(n_139187318
		));
	notech_nand2 i_2527364(.A(n_144787374), .B(n_139187318), .Z(n_16622));
	notech_nao3 i_163767714(.A(n_3511), .B(n_60605), .C(n_56428), .Z(n_139487321
		));
	notech_nand2 i_2427363(.A(n_144887375), .B(n_139487321), .Z(n_16617));
	notech_nao3 i_164367709(.A(n_3510), .B(n_60605), .C(n_56428), .Z(n_139787324
		));
	notech_nand2 i_2327362(.A(n_144987376), .B(n_139787324), .Z(n_16612));
	notech_ao4 i_182767540(.A(n_56321), .B(n_384582276), .C(n_4347), .D(n_138487311
		), .Z(n_140087327));
	notech_or2 i_19669317(.A(n_138487311), .B(n_4347), .Z(\nbus_11309[28] )
		);
	notech_nand2 i_2912923(.A(n_145687383), .B(n_30542), .Z(n_21447));
	notech_ao4 i_184467523(.A(n_56321), .B(n_384582276), .C(n_4347), .D(n_138387310
		), .Z(n_140987336));
	notech_or2 i_20669318(.A(n_138387310), .B(n_57024), .Z(\nbus_11309[26] )
		);
	notech_nand2 i_2712921(.A(n_146387390), .B(n_30543), .Z(n_21437));
	notech_ao4 i_186267506(.A(n_56321), .B(n_384582276), .C(n_57020), .D(n_138287309
		), .Z(n_141887345));
	notech_or2 i_19569319(.A(n_138287309), .B(n_57020), .Z(\nbus_11309[24] )
		);
	notech_nand2 i_2512919(.A(n_147087397), .B(n_30544), .Z(n_21427));
	notech_ao4 i_187967489(.A(n_56321), .B(n_384582276), .C(n_57020), .D(n_138187308
		), .Z(n_142787354));
	notech_or2 i_14169320(.A(n_138187308), .B(n_57020), .Z(\nbus_11309[23] )
		);
	notech_nand2 i_2412918(.A(n_147787404), .B(n_30545), .Z(n_21422));
	notech_ao4 i_189667472(.A(n_56321), .B(n_384582276), .C(n_57020), .D(n_138087307
		), .Z(n_143687363));
	notech_or2 i_20169321(.A(n_138087307), .B(n_57020), .Z(\nbus_11309[22] )
		);
	notech_nand2 i_2312917(.A(n_148487411), .B(n_30546), .Z(n_21417));
	notech_ao4 i_161267738(.A(n_56411), .B(n_58465), .C(n_61707), .D(n_32622
		), .Z(n_144587372));
	notech_ao4 i_162267728(.A(n_56411), .B(n_58447), .C(n_61707), .D(n_32620
		), .Z(n_144687373));
	notech_ao4 i_163267718(.A(n_56411), .B(n_58429), .C(n_61706), .D(n_32617
		), .Z(n_144787374));
	notech_ao4 i_163867713(.A(n_56411), .B(n_58420), .C(n_61707), .D(n_32616
		), .Z(n_144887375));
	notech_ao4 i_164467708(.A(n_56407), .B(n_58411), .C(n_61702), .D(n_32615
		), .Z(n_144987376));
	notech_ao4 i_182867539(.A(n_4348), .B(n_31536), .C(n_112042561), .D(n_32341
		), .Z(n_145087377));
	notech_ao4 i_182967538(.A(n_56359), .B(n_60564), .C(n_56330), .D(n_33579
		), .Z(n_145187378));
	notech_ao4 i_183067537(.A(n_56718), .B(n_33581), .C(n_56341), .D(n_33580
		), .Z(n_145387380));
	notech_ao4 i_183167536(.A(n_56350), .B(n_58465), .C(n_4351), .D(n_32909)
		, .Z(n_145487381));
	notech_and4 i_183467533(.A(n_145487381), .B(n_145387380), .C(n_145187378
		), .D(n_145087377), .Z(n_145687383));
	notech_ao4 i_184567522(.A(n_4348), .B(n_31534), .C(n_112042561), .D(n_32339
		), .Z(n_145787384));
	notech_ao4 i_184667521(.A(n_56359), .B(n_60582), .C(n_56330), .D(n_33582
		), .Z(n_145887385));
	notech_ao4 i_184767520(.A(n_56718), .B(n_33584), .C(n_56341), .D(n_33583
		), .Z(n_146087387));
	notech_ao4 i_184867519(.A(n_56350), .B(n_58447), .C(n_4351), .D(n_32907)
		, .Z(n_146187388));
	notech_and4 i_185267516(.A(n_146187388), .B(n_146087387), .C(n_145887385
		), .D(n_145787384), .Z(n_146387390));
	notech_ao4 i_186367505(.A(n_4348), .B(n_31532), .C(n_112042561), .D(n_32337
		), .Z(n_146487391));
	notech_ao4 i_186467504(.A(n_56359), .B(n_60519), .C(n_56330), .D(n_33585
		), .Z(n_146587392));
	notech_ao4 i_186567503(.A(n_56718), .B(n_33587), .C(n_56341), .D(n_33586
		), .Z(n_146787394));
	notech_ao4 i_186667502(.A(n_56350), .B(n_58429), .C(n_4351), .D(n_32905)
		, .Z(n_146887395));
	notech_and4 i_186967499(.A(n_146887395), .B(n_146787394), .C(n_146587392
		), .D(n_146487391), .Z(n_147087397));
	notech_ao4 i_188067488(.A(n_4348), .B(n_31531), .C(n_112042561), .D(n_32336
		), .Z(n_147187398));
	notech_ao4 i_188167487(.A(n_56359), .B(n_60528), .C(n_56330), .D(n_33588
		), .Z(n_147287399));
	notech_ao4 i_188267486(.A(n_56718), .B(n_33590), .C(n_56341), .D(n_33589
		), .Z(n_147487401));
	notech_ao4 i_188367485(.A(n_56350), .B(n_58420), .C(n_4351), .D(n_32904)
		, .Z(n_147587402));
	notech_and4 i_188667482(.A(n_147587402), .B(n_147487401), .C(n_147287399
		), .D(n_147187398), .Z(n_147787404));
	notech_ao4 i_189767471(.A(n_4348), .B(n_31530), .C(n_112042561), .D(n_32333
		), .Z(n_147887405));
	notech_ao4 i_189867470(.A(n_56359), .B(n_60537), .C(n_56330), .D(n_33591
		), .Z(n_147987406));
	notech_ao4 i_189967469(.A(n_56718), .B(n_33593), .C(n_56341), .D(n_33592
		), .Z(n_148187408));
	notech_ao4 i_190067468(.A(n_56350), .B(n_58411), .C(n_4351), .D(n_32903)
		, .Z(n_148287409));
	notech_and4 i_190367465(.A(n_148287409), .B(n_148187408), .C(n_147987406
		), .D(n_147887405), .Z(n_148487411));
	notech_ao3 i_4566111(.A(n_150687433), .B(n_323060858), .C(n_322960857), 
		.Z(n_148687413));
	notech_nao3 i_4666110(.A(n_150587432), .B(n_150987436), .C(n_150487431),
		 .Z(n_148787414));
	notech_ao4 i_066152(.A(n_163196017), .B(n_57456), .C(n_322460852), .D(n_151387440
		), .Z(n_148887415));
	notech_and4 i_4766109(.A(n_322760855), .B(n_322860856), .C(n_151487441),
		 .D(n_150187428), .Z(n_148987416));
	notech_nao3 i_101965149(.A(n_33157), .B(n_1464), .C(n_30835), .Z(n_149287419
		));
	notech_or4 i_101865150(.A(n_2383), .B(n_111445606), .C(instrc[120]), .D(n_32161
		), .Z(n_149587422));
	notech_nand2 i_101365155(.A(n_30869), .B(n_148787414), .Z(n_150087427)
		);
	notech_nand2 i_102565143(.A(n_57595), .B(n_57225), .Z(n_150187428));
	notech_and4 i_102165147(.A(instrc[101]), .B(instrc[102]), .C(n_33142), .D
		(n_29906), .Z(n_150487431));
	notech_nao3 i_102265146(.A(instrc[98]), .B(instrc[97]), .C(n_26978), .Z(n_150587432
		));
	notech_nand3 i_102065148(.A(n_57225), .B(n_63794), .C(n_57595), .Z(n_150687433
		));
	notech_ao4 i_191064283(.A(n_152787454), .B(n_30815), .C(n_30822), .D(n_152887455
		), .Z(n_150987436));
	notech_ao4 i_190064293(.A(n_30549), .B(n_148687413), .C(n_61841), .D(n_163296016
		), .Z(n_151187438));
	notech_nand3 i_190764286(.A(n_33162), .B(n_63818), .C(n_30912), .Z(n_151387440
		));
	notech_ao4 i_1766139(.A(n_57633), .B(n_2810), .C(n_30798), .D(n_57236), 
		.Z(n_151487441));
	notech_nand2 i_190564288(.A(n_322760855), .B(n_322860856), .Z(n_151687443
		));
	notech_ao4 i_189964294(.A(n_151487441), .B(n_27371), .C(n_148987416), .D
		(n_148887415), .Z(n_151787444));
	notech_ao4 i_189664297(.A(n_57225), .B(n_114845640), .C(n_26987), .D(n_37407
		), .Z(n_151987446));
	notech_and4 i_189864295(.A(n_151987446), .B(n_149287419), .C(n_149587422
		), .D(n_30519), .Z(n_152287449));
	notech_and3 i_5960581(.A(n_390564436), .B(n_387964410), .C(n_391164442),
		 .Z(n_152387450));
	notech_ao3 i_6060580(.A(n_387864409), .B(n_391264443), .C(n_390664437), 
		.Z(n_152487451));
	notech_nao3 i_31278(.A(n_32353), .B(n_32481), .C(n_1465), .Z(n_152787454
		));
	notech_nao3 i_31274(.A(n_32353), .B(n_32481), .C(n_1466), .Z(n_152887455
		));
	notech_and3 i_2560615(.A(n_339161019), .B(n_339861026), .C(n_30798), .Z(n_152987456
		));
	notech_or4 i_15360489(.A(n_63706), .B(n_386364394), .C(n_63794), .D(nbus_11273
		[13]), .Z(n_153487461));
	notech_or2 i_15060492(.A(n_386264393), .B(n_31486), .Z(n_153787464));
	notech_or2 i_16560477(.A(n_58664), .B(nbus_11271[14]), .Z(n_154287469)
		);
	notech_or4 i_16460478(.A(n_23760), .B(n_61924), .C(n_31625), .D(n_23763)
		, .Z(n_154587472));
	notech_or2 i_16160481(.A(n_23747), .B(n_33215), .Z(n_154887475));
	notech_or2 i_15860484(.A(n_377064301), .B(n_58696), .Z(n_155187478));
	notech_nao3 i_66760037(.A(n_63796), .B(opc[4]), .C(n_376764298), .Z(n_155687483
		));
	notech_or2 i_66460040(.A(n_31071), .B(n_29680), .Z(n_155987486));
	notech_nao3 i_68060025(.A(n_63788), .B(opc[4]), .C(n_29994), .Z(n_156887495
		));
	notech_or2 i_67760028(.A(n_30001), .B(n_31071), .Z(n_157187498));
	notech_nao3 i_70260003(.A(n_63728), .B(opc[4]), .C(n_30391), .Z(n_158087507
		));
	notech_or4 i_69960006(.A(n_303944473), .B(n_60169), .C(n_32266), .D(nbus_11273
		[4]), .Z(n_158387510));
	notech_ao3 i_81659889(.A(instrc[97]), .B(n_370164232), .C(n_26978), .Z(n_158887515
		));
	notech_ao3 i_81559890(.A(n_29229), .B(n_30869), .C(n_152887455), .Z(n_159187518
		));
	notech_ao3 i_81259893(.A(n_1464), .B(n_33157), .C(n_29232), .Z(n_159487521
		));
	notech_or4 i_80759898(.A(n_29584), .B(instrc[103]), .C(n_33161), .D(n_30554
		), .Z(n_159587522));
	notech_or4 i_80859897(.A(instrc[123]), .B(n_318060808), .C(n_111445606),
		 .D(instrc[120]), .Z(n_159687523));
	notech_ao4 i_80959896(.A(n_151687443), .B(n_30555), .C(n_295963857), .D(n_160287529
		), .Z(n_159787524));
	notech_and4 i_81759888(.A(n_436567949), .B(n_382964360), .C(n_33153), .D
		(n_29582), .Z(n_159987526));
	notech_or2 i_162359137(.A(n_159987526), .B(n_91234596), .Z(n_160287529)
		);
	notech_ao4 i_162159139(.A(n_57633), .B(n_2810), .C(n_152987456), .D(n_32219
		), .Z(n_160487531));
	notech_nao3 i_161859142(.A(n_159687523), .B(n_159587522), .C(n_159787524
		), .Z(n_160887535));
	notech_ao4 i_161559145(.A(n_57174), .B(n_114845640), .C(n_30553), .D(n_323060858
		), .Z(n_160987536));
	notech_ao4 i_161259148(.A(n_28572), .B(n_152787454), .C(n_26987), .D(n_30552
		), .Z(n_161287539));
	notech_or4 i_161459146(.A(n_159187518), .B(n_158887515), .C(n_4463), .D(n_30557
		), .Z(n_161587542));
	notech_ao4 i_153859221(.A(n_334660974), .B(n_323860866), .C(n_57163), .D
		(n_187176929), .Z(n_161687543));
	notech_ao4 i_153759222(.A(n_56974), .B(n_305344487), .C(n_323960867), .D
		(n_33104), .Z(n_161787544));
	notech_ao4 i_153459224(.A(n_31048), .B(n_30578), .C(n_31047), .D(n_303944473
		), .Z(n_161987546));
	notech_and4 i_154059219(.A(n_161987546), .B(n_161787544), .C(n_161687543
		), .D(n_158387510), .Z(n_162187548));
	notech_ao4 i_153159227(.A(n_30390), .B(n_31072), .C(n_30387), .D(n_31074
		), .Z(n_162287549));
	notech_ao4 i_152859229(.A(n_30394), .B(n_31075), .C(n_30393), .D(n_31068
		), .Z(n_162487551));
	notech_and4 i_153359225(.A(n_187576933), .B(n_162487551), .C(n_162287549
		), .D(n_158087507), .Z(n_162687553));
	notech_ao4 i_151659241(.A(n_30196), .B(n_334660974), .C(n_57112), .D(n_187176929
		), .Z(n_162787554));
	notech_ao4 i_151559242(.A(n_305244486), .B(n_56974), .C(n_30191), .D(n_33104
		), .Z(n_162887555));
	notech_ao4 i_151359244(.A(n_31048), .B(n_30576), .C(n_1532), .D(n_31047)
		, .Z(n_163087557));
	notech_and4 i_151859239(.A(n_163087557), .B(n_162887555), .C(n_162787554
		), .D(n_157187498), .Z(n_163287559));
	notech_ao4 i_150959247(.A(n_30002), .B(n_31072), .C(n_29998), .D(n_31074
		), .Z(n_163387560));
	notech_ao4 i_150759249(.A(n_29997), .B(n_31075), .C(n_29993), .D(n_31068
		), .Z(n_163587562));
	notech_and4 i_151259245(.A(n_187576933), .B(n_163587562), .C(n_163387560
		), .D(n_156887495), .Z(n_163787564));
	notech_ao4 i_150359252(.A(n_334660974), .B(n_376864299), .C(n_187176929)
		, .D(n_57130), .Z(n_163887565));
	notech_ao4 i_150259253(.A(n_54741988), .B(n_56974), .C(n_376964300), .D(n_33104
		), .Z(n_163987566));
	notech_ao4 i_149959255(.A(n_31048), .B(n_376564296), .C(n_31047), .D(n_94542386
		), .Z(n_164187568));
	notech_and4 i_150659250(.A(n_164187568), .B(n_163987566), .C(n_163887565
		), .D(n_155987486), .Z(n_164387570));
	notech_ao4 i_149559258(.A(n_31072), .B(n_29678), .C(n_31074), .D(n_29677
		), .Z(n_164487571));
	notech_ao4 i_149359260(.A(n_31075), .B(n_29681), .C(n_31068), .D(n_376664297
		), .Z(n_164687573));
	notech_and4 i_149859256(.A(n_187576933), .B(n_164687573), .C(n_164487571
		), .D(n_155687483), .Z(n_164887575));
	notech_ao4 i_90259803(.A(nbus_11273[14]), .B(n_152487451), .C(n_59041), 
		.D(n_152387450), .Z(n_165187578));
	notech_ao4 i_90059805(.A(n_97342414), .B(n_23750), .C(n_56035), .D(n_32543
		), .Z(n_165387580));
	notech_and4 i_90459801(.A(n_165387580), .B(n_155187478), .C(n_165187578)
		, .D(n_154887475), .Z(n_165587582));
	notech_ao4 i_89759808(.A(n_377164302), .B(n_23613), .C(n_386264393), .D(n_31487
		), .Z(n_165687583));
	notech_and4 i_89959806(.A(n_154587472), .B(n_165687583), .C(n_377364304)
		, .D(n_154287469), .Z(n_165987586));
	notech_ao4 i_89359812(.A(n_56035), .B(n_32542), .C(n_58696), .D(n_30474)
		, .Z(n_166087587));
	notech_ao4 i_89259813(.A(n_386164392), .B(\nbus_11290[13] ), .C(n_386064391
		), .D(nbus_11273[13]), .Z(n_166187588));
	notech_ao4 i_89059815(.A(n_23747), .B(n_33213), .C(n_375064281), .D(n_23750
		), .Z(n_166387590));
	notech_and4 i_89559810(.A(n_166387590), .B(n_166187588), .C(n_166087587)
		, .D(n_153787464), .Z(n_166587592));
	notech_ao4 i_88759818(.A(n_31498), .B(n_23614), .C(n_31497), .D(n_23613)
		, .Z(n_166687593));
	notech_ao4 i_88559820(.A(n_25094), .B(nbus_11271[13]), .C(n_31495), .D(n_23611
		), .Z(n_166887595));
	notech_and4 i_88959816(.A(n_166887595), .B(n_166687593), .C(n_153487461)
		, .D(n_30468), .Z(n_167087597));
	notech_or4 i_8658035(.A(n_60169), .B(n_315460782), .C(n_30652), .D(n_30649
		), .Z(n_167187598));
	notech_ao4 i_67258128(.A(n_61611), .B(n_56794), .C(n_213333664), .D(n_30649
		), .Z(n_167287599));
	notech_nand2 i_48757666(.A(n_335489239), .B(n_167487601), .Z(n_167387600
		));
	notech_or2 i_3858083(.A(n_57283), .B(n_30649), .Z(n_167487601));
	notech_or4 i_49157662(.A(n_19612), .B(n_19629), .C(n_61697), .D(n_19645)
		, .Z(n_167887605));
	notech_ao3 i_7358048(.A(Daddrs_8[0]), .B(n_61697), .C(n_391464445), .Z(n_168387610
		));
	notech_and2 i_7058051(.A(regs_4_2[0]), .B(n_212433655), .Z(n_168687613)
		);
	notech_ao3 i_6758054(.A(Daddrs_3[0]), .B(n_30680), .C(n_207687990), .Z(n_168987616
		));
	notech_nand3 i_6258059(.A(n_210633637), .B(opd[0]), .C(n_61693), .Z(n_169087617
		));
	notech_or4 i_6358058(.A(n_61711), .B(n_61878), .C(n_56794), .D(n_58956),
		 .Z(n_169187618));
	notech_nand2 i_6458057(.A(Daddrs_1[0]), .B(n_30683), .Z(n_169287619));
	notech_nao3 i_9958022(.A(Daddrs_8[2]), .B(n_61693), .C(n_391464445), .Z(n_169587622
		));
	notech_or4 i_9658025(.A(n_28007), .B(n_61614), .C(n_60152), .D(n_56965),
		 .Z(n_169887625));
	notech_or2 i_9358028(.A(n_209388005), .B(nbus_11271[2]), .Z(n_170187628)
		);
	notech_nao3 i_11258009(.A(Daddrs_8[3]), .B(n_61693), .C(n_391464445), .Z
		(n_170887635));
	notech_or4 i_10958012(.A(n_28007), .B(n_61614), .C(n_60152), .D(n_56956)
		, .Z(n_171187638));
	notech_or2 i_10658015(.A(n_209388005), .B(nbus_11271[3]), .Z(n_171487641
		));
	notech_nao3 i_12757996(.A(Daddrs_8[4]), .B(n_61697), .C(n_391464445), .Z
		(n_172187648));
	notech_or4 i_12457999(.A(n_28007), .B(n_61614), .C(n_60152), .D(n_58802)
		, .Z(n_172487651));
	notech_or2 i_12158002(.A(n_209388005), .B(nbus_11271[4]), .Z(n_172787654
		));
	notech_nao3 i_14057983(.A(Daddrs_8[5]), .B(n_61697), .C(n_391464445), .Z
		(n_173487661));
	notech_or4 i_13757986(.A(n_28007), .B(n_61611), .C(n_60152), .D(n_58784)
		, .Z(n_173787664));
	notech_or2 i_13457989(.A(n_209388005), .B(nbus_11271[5]), .Z(n_174087667
		));
	notech_nao3 i_15357970(.A(Daddrs_8[6]), .B(n_61697), .C(n_391464445), .Z
		(n_174787674));
	notech_or4 i_15057973(.A(n_28007), .B(n_61611), .C(n_60152), .D(n_56974)
		, .Z(n_175087677));
	notech_or2 i_14757976(.A(n_209388005), .B(nbus_11271[6]), .Z(n_175387680
		));
	notech_nao3 i_16657957(.A(Daddrs_8[7]), .B(n_61697), .C(n_391464445), .Z
		(n_176087687));
	notech_or4 i_16357960(.A(n_28007), .B(n_61611), .C(n_60152), .D(n_56983)
		, .Z(n_176387690));
	notech_or2 i_16057963(.A(n_209388005), .B(nbus_11271[7]), .Z(n_176687693
		));
	notech_nao3 i_17957944(.A(Daddrs_8[8]), .B(n_61697), .C(n_391464445), .Z
		(n_177387700));
	notech_or4 i_17657947(.A(n_60152), .B(n_61611), .C(n_28007), .D(n_31479)
		, .Z(n_177687703));
	notech_or2 i_17357950(.A(n_209388005), .B(nbus_11271[8]), .Z(n_177987706
		));
	notech_nao3 i_19257931(.A(Daddrs_8[9]), .B(n_61693), .C(n_391464445), .Z
		(n_178687713));
	notech_or4 i_18957934(.A(n_60152), .B(n_28007), .C(n_61611), .D(n_31480)
		, .Z(n_178987716));
	notech_or2 i_18657937(.A(n_209388005), .B(nbus_11271[9]), .Z(n_179287719
		));
	notech_nao3 i_20457919(.A(Daddrs_8[10]), .B(n_61693), .C(n_391464445), .Z
		(n_180087726));
	notech_or2 i_20157922(.A(n_30682), .B(n_32069), .Z(n_180387729));
	notech_nao3 i_19857925(.A(Daddrs_3[10]), .B(n_30680), .C(n_207687990), .Z
		(n_180687732));
	notech_nand2 i_19557928(.A(Daddrs_1[10]), .B(n_30683), .Z(n_180987735)
		);
	notech_nao3 i_22557907(.A(Daddrs_8[11]), .B(n_61693), .C(n_391464445), .Z
		(n_181287738));
	notech_or2 i_21857910(.A(n_30682), .B(n_32070), .Z(n_181587741));
	notech_nao3 i_21057913(.A(Daddrs_3[11]), .B(n_30680), .C(n_207687990), .Z
		(n_181887744));
	notech_nand2 i_20757916(.A(Daddrs_1[11]), .B(n_30683), .Z(n_182187747)
		);
	notech_nao3 i_23757895(.A(Daddrs_8[12]), .B(n_61693), .C(n_391464445), .Z
		(n_182487750));
	notech_or2 i_23457898(.A(n_30682), .B(n_32071), .Z(n_182787753));
	notech_nao3 i_23157901(.A(Daddrs_3[12]), .B(n_30680), .C(n_207687990), .Z
		(n_183287756));
	notech_nand2 i_22857904(.A(Daddrs_1[12]), .B(n_30683), .Z(n_183687759)
		);
	notech_nao3 i_25157883(.A(Daddrs_8[13]), .B(n_61693), .C(n_391464445), .Z
		(n_183987762));
	notech_or2 i_24857886(.A(n_30682), .B(n_32072), .Z(n_184487765));
	notech_nao3 i_24557889(.A(Daddrs_3[13]), .B(n_30680), .C(n_207687990), .Z
		(n_184787768));
	notech_nand2 i_24157892(.A(Daddrs_1[13]), .B(n_30683), .Z(n_185287771)
		);
	notech_nao3 i_26557871(.A(Daddrs_8[14]), .B(n_61693), .C(n_391464445), .Z
		(n_185587774));
	notech_or2 i_26157874(.A(n_30682), .B(n_32073), .Z(n_185887777));
	notech_nao3 i_25857877(.A(Daddrs_3[14]), .B(n_30680), .C(n_207687990), .Z
		(n_186187780));
	notech_nand2 i_25557880(.A(Daddrs_1[14]), .B(n_30683), .Z(n_186487783)
		);
	notech_nao3 i_27857859(.A(Daddrs_8[15]), .B(n_61693), .C(n_391464445), .Z
		(n_186787786));
	notech_or2 i_27557862(.A(n_30682), .B(n_32074), .Z(n_187087789));
	notech_nao3 i_27157865(.A(Daddrs_3[15]), .B(n_30680), .C(n_207687990), .Z
		(n_187387792));
	notech_nand2 i_26857868(.A(Daddrs_1[15]), .B(n_30683), .Z(n_187687795)
		);
	notech_nao3 i_29157847(.A(Daddrs_8[16]), .B(n_61693), .C(n_58848), .Z(n_187987798
		));
	notech_or2 i_28857850(.A(n_30682), .B(n_32075), .Z(n_188287801));
	notech_nao3 i_28557853(.A(Daddrs_3[16]), .B(n_30680), .C(n_207687990), .Z
		(n_188587804));
	notech_nand2 i_28157856(.A(Daddrs_1[16]), .B(n_30683), .Z(n_188887807)
		);
	notech_nao3 i_30757835(.A(Daddrs_8[17]), .B(n_61693), .C(n_58848), .Z(n_189187810
		));
	notech_or2 i_30057838(.A(n_30682), .B(n_32076), .Z(n_189487813));
	notech_nao3 i_29757841(.A(Daddrs_3[17]), .B(n_30680), .C(n_207687990), .Z
		(n_189787816));
	notech_nand2 i_29457844(.A(Daddrs_1[17]), .B(n_30683), .Z(n_190087819)
		);
	notech_nao3 i_32057823(.A(Daddrs_8[18]), .B(n_61693), .C(n_58848), .Z(n_190387822
		));
	notech_or2 i_31757826(.A(n_30682), .B(n_32077), .Z(n_190687825));
	notech_nao3 i_31457829(.A(Daddrs_3[18]), .B(n_30680), .C(n_207687990), .Z
		(n_190987828));
	notech_nand2 i_31157832(.A(Daddrs_1[18]), .B(n_30683), .Z(n_191287831)
		);
	notech_nao3 i_33257811(.A(Daddrs_8[19]), .B(n_61697), .C(n_58848), .Z(n_191587834
		));
	notech_or2 i_32957814(.A(n_30682), .B(n_32078), .Z(n_191887837));
	notech_nao3 i_32657817(.A(Daddrs_3[19]), .B(n_30680), .C(n_207687990), .Z
		(n_192187840));
	notech_nand2 i_32357820(.A(Daddrs_1[19]), .B(n_30683), .Z(n_192487843)
		);
	notech_nao3 i_34457799(.A(Daddrs_8[20]), .B(n_61698), .C(n_58848), .Z(n_192787846
		));
	notech_or2 i_34157802(.A(n_30682), .B(n_32079), .Z(n_193087849));
	notech_nao3 i_33857805(.A(Daddrs_3[20]), .B(n_30680), .C(n_207687990), .Z
		(n_193387852));
	notech_nand2 i_33557808(.A(Daddrs_1[20]), .B(n_30683), .Z(n_193687855)
		);
	notech_nao3 i_35657787(.A(Daddrs_8[21]), .B(n_61698), .C(n_58848), .Z(n_193987858
		));
	notech_or2 i_35357790(.A(n_30682), .B(n_32080), .Z(n_194287861));
	notech_nao3 i_35057793(.A(Daddrs_3[21]), .B(n_58628), .C(n_207687990), .Z
		(n_194587864));
	notech_nand2 i_34757796(.A(Daddrs_1[21]), .B(n_56188), .Z(n_194887867)
		);
	notech_nao3 i_36857775(.A(Daddrs_8[22]), .B(n_61698), .C(n_58848), .Z(n_195187870
		));
	notech_or2 i_36557778(.A(n_30682), .B(n_32081), .Z(n_195487873));
	notech_nao3 i_36257781(.A(Daddrs_3[22]), .B(n_58628), .C(n_207687990), .Z
		(n_195787876));
	notech_nand2 i_35957784(.A(Daddrs_1[22]), .B(n_56188), .Z(n_196087879)
		);
	notech_nao3 i_38057763(.A(Daddrs_8[23]), .B(n_61698), .C(n_58848), .Z(n_196387882
		));
	notech_or2 i_37757766(.A(n_30682), .B(n_32082), .Z(n_196687885));
	notech_nao3 i_37457769(.A(Daddrs_3[23]), .B(n_58628), .C(n_56226), .Z(n_196987888
		));
	notech_nand2 i_37157772(.A(Daddrs_1[23]), .B(n_56188), .Z(n_197287891)
		);
	notech_nao3 i_39357751(.A(Daddrs_8[24]), .B(n_61698), .C(n_58848), .Z(n_197587894
		));
	notech_or2 i_38957754(.A(n_30682), .B(n_32083), .Z(n_197887897));
	notech_nao3 i_38657757(.A(Daddrs_3[24]), .B(n_58628), .C(n_56226), .Z(n_198187900
		));
	notech_nand2 i_38357760(.A(Daddrs_1[24]), .B(n_56188), .Z(n_198487903)
		);
	notech_nao3 i_40657739(.A(Daddrs_8[25]), .B(n_61698), .C(n_58848), .Z(n_198787906
		));
	notech_or2 i_40257742(.A(n_30682), .B(n_32084), .Z(n_199187909));
	notech_nao3 i_39957745(.A(Daddrs_3[25]), .B(n_58628), .C(n_56226), .Z(n_199487912
		));
	notech_nand2 i_39657748(.A(Daddrs_1[25]), .B(n_56188), .Z(n_199787915)
		);
	notech_nao3 i_42057727(.A(Daddrs_8[26]), .B(n_61698), .C(n_58848), .Z(n_200087918
		));
	notech_or2 i_41557730(.A(n_56246), .B(n_32085), .Z(n_200487921));
	notech_nao3 i_41257733(.A(Daddrs_3[26]), .B(n_58628), .C(n_56226), .Z(n_200787924
		));
	notech_nand2 i_40957736(.A(Daddrs_1[26]), .B(n_56188), .Z(n_201087927)
		);
	notech_nao3 i_43457715(.A(Daddrs_8[27]), .B(n_61698), .C(n_58848), .Z(n_201387930
		));
	notech_or2 i_43157718(.A(n_56246), .B(n_32086), .Z(n_201687933));
	notech_nao3 i_42857721(.A(Daddrs_3[27]), .B(n_58628), .C(n_56226), .Z(n_202087936
		));
	notech_nand2 i_42457724(.A(Daddrs_1[27]), .B(n_56188), .Z(n_202387939)
		);
	notech_nao3 i_44757703(.A(Daddrs_8[28]), .B(n_61698), .C(n_58848), .Z(n_202687942
		));
	notech_or2 i_44457706(.A(n_56246), .B(n_32087), .Z(n_202987945));
	notech_nao3 i_44157709(.A(Daddrs_3[28]), .B(n_58628), .C(n_56226), .Z(n_203387948
		));
	notech_nand2 i_43857712(.A(Daddrs_1[28]), .B(n_56188), .Z(n_203687951)
		);
	notech_nao3 i_45957691(.A(Daddrs_8[29]), .B(n_61698), .C(n_58848), .Z(n_203987954
		));
	notech_or2 i_45657694(.A(n_56246), .B(n_32088), .Z(n_204287957));
	notech_nao3 i_45357697(.A(Daddrs_3[29]), .B(n_58628), .C(n_56226), .Z(n_204587960
		));
	notech_nand2 i_45057700(.A(Daddrs_1[29]), .B(n_56188), .Z(n_204887963)
		);
	notech_nao3 i_47457679(.A(Daddrs_8[30]), .B(n_61697), .C(n_58848), .Z(n_205187966
		));
	notech_or2 i_47157682(.A(n_56246), .B(n_32089), .Z(n_205487969));
	notech_nao3 i_46757685(.A(Daddrs_3[30]), .B(n_30680), .C(n_56226), .Z(n_205787972
		));
	notech_nand2 i_46457688(.A(Daddrs_1[30]), .B(n_56188), .Z(n_206087975)
		);
	notech_nao3 i_48657667(.A(Daddrs_8[31]), .B(n_61697), .C(n_58848), .Z(n_206487978
		));
	notech_or2 i_48357670(.A(n_56246), .B(n_32090), .Z(n_206787981));
	notech_nao3 i_48057673(.A(Daddrs_3[31]), .B(n_58628), .C(n_56226), .Z(n_207087984
		));
	notech_nand2 i_47757676(.A(Daddrs_1[31]), .B(n_56188), .Z(n_207387987)
		);
	notech_nand2 i_201758115(.A(n_32521), .B(n_61611), .Z(n_207687990));
	notech_nand2 i_113557044(.A(n_347671363), .B(n_347271361), .Z(n_207787991
		));
	notech_nand2 i_67358127(.A(n_167387600), .B(n_61697), .Z(n_207887992));
	notech_ao4 i_112857051(.A(n_167287599), .B(n_58983), .C(n_207887992), .D
		(n_31507), .Z(n_208187994));
	notech_or2 i_64058133(.A(n_207687990), .B(n_347271361), .Z(n_208387996)
		);
	notech_or4 i_65058131(.A(n_316160789), .B(n_56226), .C(n_315560783), .D(n_58628
		), .Z(n_208587998));
	notech_or4 i_64258132(.A(n_61917), .B(n_61903), .C(n_61877), .D(n_57915)
		, .Z(n_208687999));
	notech_ao4 i_112657053(.A(n_208687999), .B(n_33686), .C(n_208587998), .D
		(n_33685), .Z(n_208788000));
	notech_and4 i_113057049(.A(n_208788000), .B(n_208187994), .C(n_207387987
		), .D(n_207087984), .Z(n_208988002));
	notech_ao3 i_113157048(.A(n_317460802), .B(n_316260790), .C(n_301760646)
		, .Z(n_209188003));
	notech_or4 i_63058134(.A(n_60169), .B(n_32383), .C(n_32394), .D(n_61611)
		, .Z(n_209388005));
	notech_ao4 i_112357056(.A(n_31963), .B(n_212333654), .C(n_209388005), .D
		(n_60591), .Z(n_209588007));
	notech_ao4 i_112157058(.A(n_348989371), .B(n_31359), .C(n_1840), .D(n_33684
		), .Z(n_209788009));
	notech_and4 i_112557054(.A(n_209788009), .B(n_209588007), .C(n_206787981
		), .D(n_206487978), .Z(n_209988011));
	notech_ao4 i_111857061(.A(n_167287599), .B(\nbus_11290[30] ), .C(n_207887992
		), .D(n_31506), .Z(n_210088012));
	notech_ao4 i_111557063(.A(n_208687999), .B(n_33683), .C(n_208587998), .D
		(n_33682), .Z(n_210288014));
	notech_and4 i_112057059(.A(n_210288014), .B(n_210088012), .C(n_206087975
		), .D(n_205787972), .Z(n_210488016));
	notech_ao4 i_111257066(.A(n_31962), .B(n_212333654), .C(n_209388005), .D
		(n_60611), .Z(n_210588017));
	notech_ao4 i_111057068(.A(n_348989371), .B(n_31358), .C(n_1840), .D(n_33681
		), .Z(n_210788019));
	notech_and4 i_111457064(.A(n_210788019), .B(n_210588017), .C(n_205487969
		), .D(n_205187966), .Z(n_210988021));
	notech_ao4 i_110757071(.A(n_167287599), .B(n_58947), .C(n_207887992), .D
		(n_31505), .Z(n_211088022));
	notech_ao4 i_110557073(.A(n_208687999), .B(n_33680), .C(n_208587998), .D
		(n_33679), .Z(n_211288024));
	notech_and4 i_110957069(.A(n_211288024), .B(n_211088022), .C(n_204887963
		), .D(n_204587960), .Z(n_211488026));
	notech_ao4 i_110257076(.A(n_212333654), .B(n_31961), .C(n_209388005), .D
		(n_60620), .Z(n_211588027));
	notech_ao4 i_110057078(.A(n_348989371), .B(n_31357), .C(n_1840), .D(n_33678
		), .Z(n_211788029));
	notech_and4 i_110457074(.A(n_211788029), .B(n_211588027), .C(n_204287957
		), .D(n_203987954), .Z(n_211988031));
	notech_ao4 i_109757081(.A(n_167287599), .B(n_58929), .C(n_207887992), .D
		(n_31504), .Z(n_212088032));
	notech_ao4 i_109557083(.A(n_208687999), .B(n_33677), .C(n_208587998), .D
		(n_33676), .Z(n_212288034));
	notech_and4 i_109957079(.A(n_212288034), .B(n_212088032), .C(n_203687951
		), .D(n_203387948), .Z(n_212488036));
	notech_ao4 i_109257086(.A(n_31960), .B(n_212333654), .C(n_60564), .D(n_209388005
		), .Z(n_212588037));
	notech_ao4 i_109057088(.A(n_348989371), .B(n_31356), .C(n_1840), .D(n_33675
		), .Z(n_212788039));
	notech_and4 i_109457084(.A(n_212788039), .B(n_212588037), .C(n_202987945
		), .D(n_202687942), .Z(n_212988041));
	notech_ao4 i_108757091(.A(n_167287599), .B(n_58938), .C(n_207887992), .D
		(n_31503), .Z(n_213188042));
	notech_ao4 i_108557093(.A(n_208687999), .B(n_33674), .C(n_208587998), .D
		(n_33673), .Z(n_213388044));
	notech_and4 i_108957089(.A(n_213388044), .B(n_213188042), .C(n_202387939
		), .D(n_202087936), .Z(n_213588046));
	notech_ao4 i_108257096(.A(n_31959), .B(n_212333654), .C(n_60573), .D(n_209388005
		), .Z(n_213688047));
	notech_ao4 i_108057098(.A(n_348989371), .B(n_31355), .C(n_1840), .D(n_33672
		), .Z(n_213888049));
	notech_and4 i_108457094(.A(n_213888049), .B(n_213688047), .C(n_201687933
		), .D(n_201387930), .Z(n_214088051));
	notech_ao4 i_107557101(.A(n_167287599), .B(n_58911), .C(n_207887992), .D
		(n_31502), .Z(n_214188052));
	notech_ao4 i_107257103(.A(n_208687999), .B(n_33671), .C(n_208587998), .D
		(n_33670), .Z(n_214388054));
	notech_and4 i_107857099(.A(n_214388054), .B(n_214188052), .C(n_201087927
		), .D(n_200787924), .Z(n_214588056));
	notech_ao4 i_106957106(.A(n_31958), .B(n_212333654), .C(n_60582), .D(n_209388005
		), .Z(n_214688057));
	notech_ao4 i_106757108(.A(n_348989371), .B(n_31354), .C(n_1840), .D(n_33669
		), .Z(n_214888059));
	notech_and4 i_107157104(.A(n_214888059), .B(n_214688057), .C(n_200487921
		), .D(n_200087918), .Z(n_215088061));
	notech_ao4 i_106457111(.A(n_167287599), .B(\nbus_11290[25] ), .C(n_207887992
		), .D(n_31501), .Z(n_215188062));
	notech_ao4 i_106257113(.A(n_208687999), .B(n_33668), .C(n_208587998), .D
		(n_33667), .Z(n_215388064));
	notech_and4 i_106657109(.A(n_215388064), .B(n_215188062), .C(n_199787915
		), .D(n_199487912), .Z(n_215588066));
	notech_ao4 i_105857116(.A(n_31957), .B(n_212333654), .C(n_209388005), .D
		(n_60510), .Z(n_215688067));
	notech_ao4 i_105657118(.A(n_348989371), .B(n_31353), .C(n_1840), .D(n_33666
		), .Z(n_215888069));
	notech_and4 i_106057114(.A(n_215888069), .B(n_215688067), .C(n_199187909
		), .D(n_198787906), .Z(n_216088071));
	notech_ao4 i_105357121(.A(n_167287599), .B(n_58893), .C(n_207887992), .D
		(n_31500), .Z(n_216188072));
	notech_ao4 i_105157123(.A(n_208687999), .B(n_33665), .C(n_208587998), .D
		(n_33664), .Z(n_216388074));
	notech_and4 i_105557119(.A(n_216388074), .B(n_216188072), .C(n_198487903
		), .D(n_198187900), .Z(n_216588076));
	notech_ao4 i_104857126(.A(n_31956), .B(n_212333654), .C(n_60519), .D(n_209388005
		), .Z(n_216688077));
	notech_ao4 i_104657128(.A(n_348989371), .B(n_31352), .C(n_1840), .D(n_33663
		), .Z(n_216888079));
	notech_and4 i_105057124(.A(n_216888079), .B(n_216688077), .C(n_197887897
		), .D(n_197587894), .Z(n_217088081));
	notech_ao4 i_104357131(.A(n_167287599), .B(n_58902), .C(n_207887992), .D
		(n_31499), .Z(n_217188082));
	notech_ao4 i_104157133(.A(n_208687999), .B(n_33662), .C(n_208587998), .D
		(n_33661), .Z(n_217388084));
	notech_and4 i_104557129(.A(n_217388084), .B(n_217188082), .C(n_197287891
		), .D(n_196987888), .Z(n_217588086));
	notech_ao4 i_103857136(.A(n_212333654), .B(n_31955), .C(n_56257), .D(n_60528
		), .Z(n_217688087));
	notech_ao4 i_103557138(.A(n_348989371), .B(n_31351), .C(n_1840), .D(n_33660
		), .Z(n_217988089));
	notech_and4 i_104057134(.A(n_217988089), .B(n_217688087), .C(n_196687885
		), .D(n_196387882), .Z(n_218188091));
	notech_ao4 i_103257141(.A(n_167287599), .B(n_58875), .C(n_207887992), .D
		(n_31496), .Z(n_218288092));
	notech_ao4 i_103057143(.A(n_208687999), .B(n_33659), .C(n_208587998), .D
		(n_33658), .Z(n_218488094));
	notech_and4 i_103457139(.A(n_218488094), .B(n_218288092), .C(n_196087879
		), .D(n_195787876), .Z(n_218688096));
	notech_ao4 i_102757146(.A(n_31954), .B(n_212333654), .C(n_56257), .D(n_60537
		), .Z(n_218788097));
	notech_ao4 i_102557148(.A(n_348989371), .B(n_31350), .C(n_1840), .D(n_33657
		), .Z(n_218988099));
	notech_and4 i_102957144(.A(n_218988099), .B(n_218788097), .C(n_195487873
		), .D(n_195187870), .Z(n_219188101));
	notech_ao4 i_102257151(.A(n_167287599), .B(n_58884), .C(n_207887992), .D
		(n_31494), .Z(n_219288102));
	notech_ao4 i_102057153(.A(n_208687999), .B(n_33656), .C(n_208587998), .D
		(n_33655), .Z(n_219488104));
	notech_and4 i_102457149(.A(n_219488104), .B(n_219288102), .C(n_194887867
		), .D(n_194587864), .Z(n_219688106));
	notech_ao4 i_101757156(.A(n_212333654), .B(n_31953), .C(n_56257), .D(n_60546
		), .Z(n_219788107));
	notech_ao4 i_101557158(.A(n_348989371), .B(n_31349), .C(n_1840), .D(n_33654
		), .Z(n_219988109));
	notech_and4 i_101957154(.A(n_219988109), .B(n_219788107), .C(n_194287861
		), .D(n_193987858), .Z(n_220188111));
	notech_ao4 i_101257161(.A(n_167287599), .B(n_58857), .C(n_207887992), .D
		(n_31493), .Z(n_220288112));
	notech_ao4 i_100957163(.A(n_208687999), .B(n_33653), .C(n_208587998), .D
		(n_33652), .Z(n_220488114));
	notech_and4 i_101457159(.A(n_220488114), .B(n_220288112), .C(n_193687855
		), .D(n_193387852), .Z(n_220688116));
	notech_ao4 i_100657166(.A(n_31952), .B(n_212333654), .C(n_56257), .D(n_60555
		), .Z(n_220788117));
	notech_ao4 i_100457168(.A(n_348989371), .B(n_31348), .C(n_1840), .D(n_33651
		), .Z(n_220988119));
	notech_and4 i_100857164(.A(n_220988119), .B(n_220788117), .C(n_193087849
		), .D(n_192787846), .Z(n_221188121));
	notech_ao4 i_100157171(.A(n_167287599), .B(n_58866), .C(n_207887992), .D
		(n_31492), .Z(n_221288122));
	notech_ao4 i_99957173(.A(n_208687999), .B(n_33650), .C(n_208587998), .D(n_33649
		), .Z(n_221488124));
	notech_and4 i_100357169(.A(n_221488124), .B(n_221288122), .C(n_192487843
		), .D(n_192187840), .Z(n_221688126));
	notech_ao4 i_99657176(.A(n_31951), .B(n_212333654), .C(n_60483), .D(n_56257
		), .Z(n_221788127));
	notech_ao4 i_99457178(.A(n_348989371), .B(n_31347), .C(n_1840), .D(n_33648
		), .Z(n_221988129));
	notech_and4 i_99857174(.A(n_221988129), .B(n_221788127), .C(n_191887837)
		, .D(n_191587834), .Z(n_222188131));
	notech_ao4 i_99157181(.A(n_167287599), .B(n_59077), .C(n_207887992), .D(n_31491
		), .Z(n_222288132));
	notech_ao4 i_98957183(.A(n_208687999), .B(n_33647), .C(n_208587998), .D(n_33646
		), .Z(n_222488134));
	notech_and4 i_99357179(.A(n_222488134), .B(n_222288132), .C(n_191287831)
		, .D(n_190987828), .Z(n_222688136));
	notech_ao4 i_98657186(.A(n_31950), .B(n_212333654), .C(n_60492), .D(n_56257
		), .Z(n_222788137));
	notech_ao4 i_98457188(.A(n_348989371), .B(n_31346), .C(n_1840), .D(n_33645
		), .Z(n_222988139));
	notech_and4 i_98857184(.A(n_222988139), .B(n_222788137), .C(n_190687825)
		, .D(n_190387822), .Z(n_223188141));
	notech_ao4 i_98157191(.A(n_167287599), .B(n_59086), .C(n_207887992), .D(n_31490
		), .Z(n_223288142));
	notech_ao4 i_97957193(.A(n_208687999), .B(n_33644), .C(n_208587998), .D(n_33643
		), .Z(n_223488144));
	notech_and4 i_98357189(.A(n_223488144), .B(n_223288142), .C(n_190087819)
		, .D(n_189787816), .Z(n_223688146));
	notech_ao4 i_97657196(.A(n_31949), .B(n_212333654), .C(n_60501), .D(n_56257
		), .Z(n_223788147));
	notech_ao4 i_97457198(.A(n_348989371), .B(n_31345), .C(n_1840), .D(n_33642
		), .Z(n_223988149));
	notech_and4 i_97857194(.A(n_223988149), .B(n_223788147), .C(n_189487813)
		, .D(n_189187810), .Z(n_224188151));
	notech_ao4 i_97057201(.A(n_56206), .B(n_59059), .C(n_56197), .D(n_31489)
		, .Z(n_224288152));
	notech_ao4 i_96857203(.A(n_208687999), .B(n_33641), .C(n_208587998), .D(n_33640
		), .Z(n_224488154));
	notech_and4 i_97357199(.A(n_224488154), .B(n_224288152), .C(n_188887807)
		, .D(n_188587804), .Z(n_224688156));
	notech_ao4 i_96557206(.A(n_212333654), .B(n_31948), .C(n_56257), .D(n_60474
		), .Z(n_224788157));
	notech_ao4 i_96357208(.A(n_348989371), .B(n_31344), .C(n_58646), .D(n_33639
		), .Z(n_224988159));
	notech_and4 i_96757204(.A(n_224988159), .B(n_224788157), .C(n_188287801)
		, .D(n_187987798), .Z(n_225188161));
	notech_ao4 i_96057211(.A(n_56206), .B(\nbus_11290[15] ), .C(n_56197), .D
		(n_31488), .Z(n_225288162));
	notech_ao4 i_95857213(.A(n_56235), .B(n_33638), .C(n_56215), .D(n_33637)
		, .Z(n_225488164));
	notech_and4 i_96257209(.A(n_225488164), .B(n_225288162), .C(n_187687795)
		, .D(n_187387792), .Z(n_225688166));
	notech_ao4 i_95557216(.A(n_31947), .B(n_56268), .C(n_56257), .D(nbus_11271
		[15]), .Z(n_225788167));
	notech_ao4 i_95357218(.A(n_348989371), .B(n_31343), .C(n_58646), .D(n_33636
		), .Z(n_225988169));
	notech_and4 i_95757214(.A(n_225988169), .B(n_225788167), .C(n_187087789)
		, .D(n_186787786), .Z(n_226188171));
	notech_ao4 i_95057221(.A(n_56206), .B(n_59041), .C(n_56197), .D(n_31487)
		, .Z(n_226288172));
	notech_ao4 i_94857223(.A(n_56235), .B(n_33635), .C(n_56215), .D(n_33634)
		, .Z(n_226488174));
	notech_and4 i_95257219(.A(n_226488174), .B(n_226288172), .C(n_186487783)
		, .D(n_186187780), .Z(n_226688176));
	notech_ao4 i_94557226(.A(n_31946), .B(n_56268), .C(n_56257), .D(nbus_11271
		[14]), .Z(n_226788177));
	notech_ao4 i_94357228(.A(n_58619), .B(n_31342), .C(n_58646), .D(n_33633)
		, .Z(n_226988179));
	notech_and4 i_94757224(.A(n_226988179), .B(n_226788177), .C(n_185887777)
		, .D(n_185587774), .Z(n_227188181));
	notech_ao4 i_94057231(.A(n_56206), .B(\nbus_11290[13] ), .C(n_56197), .D
		(n_31486), .Z(n_227288182));
	notech_ao4 i_93857233(.A(n_56235), .B(n_33632), .C(n_56215), .D(n_33631)
		, .Z(n_227488184));
	notech_and4 i_94257229(.A(n_227488184), .B(n_227288182), .C(n_185287771)
		, .D(n_184787768), .Z(n_227688186));
	notech_ao4 i_93557236(.A(n_31945), .B(n_56268), .C(n_56257), .D(nbus_11271
		[13]), .Z(n_227788187));
	notech_ao4 i_93357238(.A(n_58619), .B(n_31341), .C(n_58646), .D(n_33630)
		, .Z(n_227988189));
	notech_and4 i_93757234(.A(n_227988189), .B(n_227788187), .C(n_184487765)
		, .D(n_183987762), .Z(n_228188191));
	notech_ao4 i_93057241(.A(n_56206), .B(n_59050), .C(n_56197), .D(n_31485)
		, .Z(n_228288192));
	notech_ao4 i_92857243(.A(n_56235), .B(n_33629), .C(n_56215), .D(n_33628)
		, .Z(n_228488194));
	notech_and4 i_93257239(.A(n_228488194), .B(n_228288192), .C(n_183687759)
		, .D(n_183287756), .Z(n_228688196));
	notech_ao4 i_92557246(.A(n_31944), .B(n_56268), .C(n_56257), .D(nbus_11271
		[12]), .Z(n_228788197));
	notech_ao4 i_92357248(.A(n_58619), .B(n_31340), .C(n_58646), .D(n_33627)
		, .Z(n_228988199));
	notech_and4 i_92757244(.A(n_228988199), .B(n_228788197), .C(n_182787753)
		, .D(n_182487750), .Z(n_229188201));
	notech_ao4 i_92057251(.A(n_56206), .B(n_58974), .C(n_56197), .D(n_31484)
		, .Z(n_229288202));
	notech_ao4 i_91857253(.A(n_56235), .B(n_33626), .C(n_56215), .D(n_33625)
		, .Z(n_229488204));
	notech_and4 i_92257249(.A(n_229488204), .B(n_229288202), .C(n_182187747)
		, .D(n_181887744), .Z(n_229688206));
	notech_ao4 i_91557256(.A(n_31943), .B(n_56268), .C(n_56257), .D(nbus_11271
		[11]), .Z(n_229788207));
	notech_ao4 i_91357258(.A(n_58619), .B(n_31339), .C(n_58646), .D(n_33624)
		, .Z(n_229988209));
	notech_and4 i_91757254(.A(n_229988209), .B(n_229788207), .C(n_181587741)
		, .D(n_181287738), .Z(n_230188211));
	notech_ao4 i_91057261(.A(n_56206), .B(\nbus_11290[10] ), .C(n_56197), .D
		(n_31483), .Z(n_230288212));
	notech_ao4 i_90857263(.A(n_56235), .B(n_33623), .C(n_56215), .D(n_33622)
		, .Z(n_230488214));
	notech_and4 i_91257259(.A(n_230488214), .B(n_230288212), .C(n_180987735)
		, .D(n_180687732), .Z(n_230688216));
	notech_ao4 i_90557266(.A(n_31941), .B(n_56268), .C(nbus_11271[10]), .D(n_56257
		), .Z(n_230788217));
	notech_ao4 i_90357268(.A(n_58619), .B(n_31338), .C(n_58646), .D(n_33621)
		, .Z(n_230988219));
	notech_and4 i_90757264(.A(n_230988219), .B(n_230788217), .C(n_180387729)
		, .D(n_180087726), .Z(n_231188221));
	notech_ao4 i_90057271(.A(n_56206), .B(n_59032), .C(n_56197), .D(n_31482)
		, .Z(n_231288222));
	notech_ao4 i_89957272(.A(n_56215), .B(n_33620), .C(n_211833649), .D(n_32664
		), .Z(n_231388223));
	notech_ao4 i_89757274(.A(n_208387996), .B(n_32655), .C(n_56235), .D(n_33619
		), .Z(n_231588225));
	notech_and4 i_90257269(.A(n_231588225), .B(n_231388223), .C(n_231288222)
		, .D(n_179287719), .Z(n_231788227));
	notech_ao4 i_89457277(.A(n_56246), .B(n_32068), .C(n_31940), .D(n_56268)
		, .Z(n_231888228));
	notech_ao4 i_89257279(.A(n_58619), .B(n_31337), .C(n_58646), .D(n_33618)
		, .Z(n_232088230));
	notech_and4 i_89657275(.A(n_232088230), .B(n_231888228), .C(n_178987716)
		, .D(n_178687713), .Z(n_232288232));
	notech_ao4 i_88757282(.A(n_56206), .B(\nbus_11290[8] ), .C(n_31481), .D(n_56197
		), .Z(n_232388233));
	notech_ao4 i_88657283(.A(n_56215), .B(n_33617), .C(n_211833649), .D(n_32662
		), .Z(n_232488234));
	notech_ao4 i_88457285(.A(n_208387996), .B(n_32654), .C(n_56235), .D(n_33616
		), .Z(n_232688236));
	notech_and4 i_89157280(.A(n_232688236), .B(n_232488234), .C(n_232388233)
		, .D(n_177987706), .Z(n_232888238));
	notech_ao4 i_88157288(.A(n_56246), .B(n_32067), .C(n_31939), .D(n_56268)
		, .Z(n_232988239));
	notech_ao4 i_87957290(.A(n_58619), .B(n_31336), .C(n_58646), .D(n_33615)
		, .Z(n_233188241));
	notech_and4 i_88357286(.A(n_233188241), .B(n_177687703), .C(n_232988239)
		, .D(n_177387700), .Z(n_233388243));
	notech_ao4 i_87657293(.A(n_56206), .B(\nbus_11290[7] ), .C(n_56197), .D(n_31480
		), .Z(n_233488244));
	notech_ao4 i_87557294(.A(n_56215), .B(n_33614), .C(n_211833649), .D(n_32661
		), .Z(n_233588245));
	notech_ao4 i_87357296(.A(n_208387996), .B(n_32653), .C(n_56235), .D(n_33613
		), .Z(n_233788247));
	notech_and4 i_87857291(.A(n_233788247), .B(n_233588245), .C(n_233488244)
		, .D(n_176687693), .Z(n_233988249));
	notech_ao4 i_87057299(.A(n_56246), .B(n_32066), .C(n_56268), .D(n_31938)
		, .Z(n_234088250));
	notech_ao4 i_86857301(.A(n_58619), .B(n_31335), .C(n_58646), .D(n_33612)
		, .Z(n_234288252));
	notech_and4 i_87257297(.A(n_234288252), .B(n_176387690), .C(n_234088250)
		, .D(n_176087687), .Z(n_234488254));
	notech_ao4 i_86557304(.A(n_56206), .B(\nbus_11290[6] ), .C(n_56197), .D(n_31479
		), .Z(n_234588255));
	notech_ao4 i_86457305(.A(n_56215), .B(n_33611), .C(n_211833649), .D(n_32660
		), .Z(n_234688256));
	notech_ao4 i_86257307(.A(n_208387996), .B(n_32652), .C(n_56235), .D(n_33610
		), .Z(n_234888258));
	notech_and4 i_86757302(.A(n_234888258), .B(n_234688256), .C(n_234588255)
		, .D(n_175387680), .Z(n_235088260));
	notech_ao4 i_85957310(.A(n_56246), .B(n_32065), .C(n_31937), .D(n_56268)
		, .Z(n_235188261));
	notech_ao4 i_85757312(.A(n_58619), .B(n_31334), .C(n_58646), .D(n_33609)
		, .Z(n_235388263));
	notech_and4 i_86157308(.A(n_235388263), .B(n_175087677), .C(n_235188261)
		, .D(n_174787674), .Z(n_235588265));
	notech_ao4 i_85457315(.A(n_56206), .B(\nbus_11290[5] ), .C(n_56197), .D(n_56983
		), .Z(n_235688266));
	notech_ao4 i_85357316(.A(n_56215), .B(n_33608), .C(n_211833649), .D(n_32659
		), .Z(n_235788267));
	notech_ao4 i_85157318(.A(n_208387996), .B(n_32651), .C(n_56235), .D(n_33607
		), .Z(n_235988269));
	notech_and4 i_85657313(.A(n_235988269), .B(n_235788267), .C(n_235688266)
		, .D(n_174087667), .Z(n_236188271));
	notech_ao4 i_84857321(.A(n_56246), .B(n_32064), .C(n_31936), .D(n_56268)
		, .Z(n_236288272));
	notech_ao4 i_84657323(.A(n_58619), .B(n_31333), .C(n_1840), .D(n_33606),
		 .Z(n_236488274));
	notech_and4 i_85057319(.A(n_236488274), .B(n_173787664), .C(n_236288272)
		, .D(n_173487661), .Z(n_236688276));
	notech_ao4 i_84357326(.A(n_56206), .B(\nbus_11290[4] ), .C(n_56197), .D(n_56974
		), .Z(n_236788277));
	notech_ao4 i_84257327(.A(n_56215), .B(n_33605), .C(n_211833649), .D(n_32658
		), .Z(n_236888278));
	notech_ao4 i_83957329(.A(n_208387996), .B(n_32649), .C(n_56235), .D(n_33604
		), .Z(n_237088280));
	notech_and4 i_84557324(.A(n_237088280), .B(n_236888278), .C(n_236788277)
		, .D(n_172787654), .Z(n_237288282));
	notech_ao4 i_83657332(.A(n_56246), .B(n_32063), .C(n_31935), .D(n_56268)
		, .Z(n_237388283));
	notech_ao4 i_83357334(.A(n_348989371), .B(n_31332), .C(n_58646), .D(n_33603
		), .Z(n_237588285));
	notech_and4 i_83857330(.A(n_237588285), .B(n_172487651), .C(n_237388283)
		, .D(n_172187648), .Z(n_237788287));
	notech_ao4 i_83057337(.A(n_56206), .B(\nbus_11290[3] ), .C(n_56197), .D(n_58784
		), .Z(n_237888288));
	notech_ao4 i_82957338(.A(n_56215), .B(n_33602), .C(n_211833649), .D(n_32657
		), .Z(n_237988289));
	notech_ao4 i_82757340(.A(n_208387996), .B(n_32648), .C(n_56235), .D(n_33601
		), .Z(n_238188291));
	notech_and4 i_83257335(.A(n_238188291), .B(n_237988289), .C(n_237888288)
		, .D(n_171487641), .Z(n_238388293));
	notech_ao4 i_82357343(.A(n_56246), .B(n_32062), .C(n_31934), .D(n_56268)
		, .Z(n_238488294));
	notech_ao4 i_82157345(.A(n_58619), .B(n_31331), .C(n_58646), .D(n_33600)
		, .Z(n_238688296));
	notech_and4 i_82657341(.A(n_238688296), .B(n_171187638), .C(n_238488294)
		, .D(n_170887635), .Z(n_238888298));
	notech_ao4 i_81757348(.A(n_56206), .B(\nbus_11290[2] ), .C(n_56197), .D(n_58802
		), .Z(n_238988299));
	notech_ao4 i_81657349(.A(n_56215), .B(n_33599), .C(n_211833649), .D(n_32656
		), .Z(n_239088300));
	notech_ao4 i_81357351(.A(n_208387996), .B(n_32647), .C(n_56235), .D(n_33598
		), .Z(n_239288302));
	notech_and4 i_82057346(.A(n_239288302), .B(n_239088300), .C(n_238988299)
		, .D(n_170187628), .Z(n_239488304));
	notech_ao4 i_81057354(.A(n_56246), .B(n_32061), .C(n_31933), .D(n_56268)
		, .Z(n_239588305));
	notech_ao4 i_80857356(.A(n_58619), .B(n_31330), .C(n_58646), .D(n_33597)
		, .Z(n_239788307));
	notech_and4 i_81257352(.A(n_239788307), .B(n_169887625), .C(n_239588305)
		, .D(n_169587622), .Z(n_239988309));
	notech_nand3 i_79257371(.A(n_169187618), .B(n_169087617), .C(n_169287619
		), .Z(n_240388313));
	notech_ao4 i_78957374(.A(n_56235), .B(n_33596), .C(n_56215), .D(n_33595)
		, .Z(n_240488314));
	notech_ao4 i_78657377(.A(n_56268), .B(n_31931), .C(n_56257), .D(nbus_11271
		[0]), .Z(n_240788317));
	notech_ao4 i_78457379(.A(n_58619), .B(n_31328), .C(n_58646), .D(n_33594)
		, .Z(n_240988319));
	notech_or4 i_78857375(.A(n_168387610), .B(n_168687613), .C(n_30569), .D(n_30568
		), .Z(n_241188321));
	notech_nor2 i_59555371(.A(n_28867), .B(n_60582), .Z(n_241288322));
	notech_nao3 i_59055376(.A(n_57386), .B(opd[26]), .C(n_57187), .Z(n_241988329
		));
	notech_nor2 i_60355363(.A(n_28867), .B(n_60573), .Z(n_242088330));
	notech_nao3 i_59855368(.A(n_57386), .B(opd[27]), .C(n_57187), .Z(n_243188337
		));
	notech_nao3 i_68655280(.A(n_57386), .B(opd[27]), .C(n_57057), .Z(n_244188345
		));
	notech_nor2 i_71555251(.A(n_443668020), .B(n_60582), .Z(n_244288346));
	notech_ao3 i_71055256(.A(n_57382), .B(opd[26]), .C(n_57130), .Z(n_245088353
		));
	notech_nor2 i_72355243(.A(n_443668020), .B(n_60573), .Z(n_245188354));
	notech_ao3 i_71855248(.A(n_57386), .B(opd[27]), .C(n_57130), .Z(n_245988361
		));
	notech_ao4 i_157854414(.A(n_443968023), .B(n_284131522), .C(n_444068024)
		, .D(n_172669762), .Z(n_246088362));
	notech_ao4 i_157754415(.A(n_119326520), .B(n_5711), .C(n_119226519), .D(n_33195
		), .Z(n_246288364));
	notech_nao3 i_158054412(.A(n_246088362), .B(n_246288364), .C(n_245988361
		), .Z(n_246388365));
	notech_ao4 i_157554417(.A(n_443768021), .B(n_58456), .C(n_443868022), .D
		(n_58938), .Z(n_246488366));
	notech_ao4 i_157154421(.A(n_284231523), .B(n_443968023), .C(n_444068024)
		, .D(n_175169787), .Z(n_246888369));
	notech_ao4 i_157054422(.A(n_119326520), .B(n_5720), .C(n_119226519), .D(n_33198
		), .Z(n_247088371));
	notech_nao3 i_157354419(.A(n_246888369), .B(n_247088371), .C(n_245088353
		), .Z(n_247188372));
	notech_ao4 i_156854424(.A(n_443768021), .B(n_58447), .C(n_443868022), .D
		(\nbus_11290[26] ), .Z(n_247288373));
	notech_ao4 i_154354448(.A(n_284131522), .B(n_303822063), .C(n_172669762)
		, .D(n_299122016), .Z(n_247588376));
	notech_ao4 i_154254449(.A(n_57320), .B(n_5711), .C(n_57319), .D(n_33195)
		, .Z(n_247788378));
	notech_and3 i_154554446(.A(n_247588376), .B(n_247788378), .C(n_244188345
		), .Z(n_247888379));
	notech_ao4 i_154054451(.A(n_57363), .B(n_58456), .C(n_57362), .D(\nbus_11290[27] 
		), .Z(n_247988380));
	notech_ao4 i_153954452(.A(n_31535), .B(n_61697), .C(n_303922064), .D(n_60573
		), .Z(n_248088381));
	notech_ao4 i_142854562(.A(n_284131522), .B(n_28852), .C(n_172669762), .D
		(n_28869), .Z(n_248288383));
	notech_ao4 i_142754563(.A(n_5711), .B(n_388264413), .C(n_388364414), .D(n_33195
		), .Z(n_248488385));
	notech_nand3 i_143054560(.A(n_248288383), .B(n_248488385), .C(n_243188337
		), .Z(n_248588386));
	notech_ao4 i_142554565(.A(n_28874), .B(n_58456), .C(n_28863), .D(n_58938
		), .Z(n_248688387));
	notech_ao4 i_142154569(.A(n_284231523), .B(n_28852), .C(n_175169787), .D
		(n_28869), .Z(n_248988390));
	notech_ao4 i_142054570(.A(n_5720), .B(n_388264413), .C(n_388364414), .D(n_33198
		), .Z(n_249188392));
	notech_nand3 i_142354567(.A(n_248988390), .B(n_249188392), .C(n_241988329
		), .Z(n_249288393));
	notech_ao4 i_141854572(.A(n_28874), .B(n_58447), .C(n_28863), .D(n_58911
		), .Z(n_249388394));
	notech_nor2 i_57749175(.A(n_28867), .B(n_60474), .Z(n_249688397));
	notech_nao3 i_57249180(.A(n_57386), .B(opd[16]), .C(n_57187), .Z(n_250388404
		));
	notech_nor2 i_58549167(.A(n_28867), .B(n_60501), .Z(n_250488405));
	notech_nao3 i_58049172(.A(n_57382), .B(opd[17]), .C(n_57187), .Z(n_251188412
		));
	notech_nor2 i_59349159(.A(n_28867), .B(n_60492), .Z(n_251288413));
	notech_nao3 i_58849164(.A(n_57378), .B(opd[18]), .C(n_57187), .Z(n_251988420
		));
	notech_nand3 i_66249090(.A(n_57378), .B(n_32211), .C(opd[16]), .Z(n_252788428
		));
	notech_nand3 i_67049082(.A(n_57378), .B(n_32211), .C(opd[17]), .Z(n_253588436
		));
	notech_nand3 i_67849074(.A(n_57378), .B(n_32211), .C(opd[18]), .Z(n_254388444
		));
	notech_nand3 i_68649066(.A(n_57378), .B(n_32211), .C(opd[19]), .Z(n_255188452
		));
	notech_or2 i_70149051(.A(n_54741988), .B(n_58784), .Z(n_255688457));
	notech_or4 i_69849054(.A(n_63706), .B(n_376564296), .C(n_61924), .D(n_58256
		), .Z(n_255988460));
	notech_and3 i_71149041(.A(n_57378), .B(n_32224), .C(opd[16]), .Z(n_256488465
		));
	notech_or2 i_70649046(.A(n_443668020), .B(n_60474), .Z(n_257188472));
	notech_and3 i_71949033(.A(n_57382), .B(n_32224), .C(opd[17]), .Z(n_257288473
		));
	notech_or2 i_71449038(.A(n_443668020), .B(n_60501), .Z(n_257988480));
	notech_and3 i_72749025(.A(n_57382), .B(n_32224), .C(opd[18]), .Z(n_258088481
		));
	notech_or2 i_72249030(.A(n_443668020), .B(n_60492), .Z(n_258788488));
	notech_and3 i_73549017(.A(n_57382), .B(n_32224), .C(opd[19]), .Z(n_258888489
		));
	notech_or2 i_73049022(.A(n_443668020), .B(n_60483), .Z(n_259588496));
	notech_or2 i_74549007(.A(n_305244486), .B(n_58784), .Z(n_260088501));
	notech_or4 i_74249010(.A(n_63706), .B(n_61924), .C(n_58256), .D(n_30576)
		, .Z(n_260388504));
	notech_nand2 i_78948963(.A(opd[3]), .B(n_30630), .Z(n_261288513));
	notech_or4 i_78648966(.A(n_60188), .B(n_55831), .C(n_303944473), .D(n_58256
		), .Z(n_261588516));
	notech_ao4 i_186847925(.A(n_74922852), .B(n_30391), .C(n_66222765), .D(n_57163
		), .Z(n_262088521));
	notech_ao4 i_186747926(.A(n_75322856), .B(n_30386), .C(n_75222855), .D(n_30394
		), .Z(n_262188522));
	notech_ao4 i_186547928(.A(n_75522858), .B(n_30387), .C(n_75622859), .D(n_30390
		), .Z(n_262388524));
	notech_and4 i_187047923(.A(n_262388524), .B(n_262188522), .C(n_262088521
		), .D(n_261588516), .Z(n_262588526));
	notech_ao4 i_186247931(.A(n_74522848), .B(n_30393), .C(n_303944473), .D(n_74622849
		), .Z(n_262688527));
	notech_ao4 i_186047933(.A(n_33118), .B(n_323960867), .C(n_338361011), .D
		(n_323860866), .Z(n_262888529));
	notech_and4 i_186447929(.A(n_65022753), .B(n_262888529), .C(n_262688527)
		, .D(n_261288513), .Z(n_263088531));
	notech_ao4 i_182947964(.A(n_74922852), .B(n_29994), .C(n_66222765), .D(n_57112
		), .Z(n_263188532));
	notech_ao4 i_182847965(.A(n_75322856), .B(n_30001), .C(n_75222855), .D(n_29997
		), .Z(n_263288533));
	notech_ao4 i_182647967(.A(n_75522858), .B(n_29998), .C(n_75622859), .D(n_30002
		), .Z(n_263488535));
	notech_and4 i_183147962(.A(n_263488535), .B(n_263288533), .C(n_263188532
		), .D(n_260388504), .Z(n_263688537));
	notech_ao4 i_182347970(.A(n_74522848), .B(n_29993), .C(n_74622849), .D(n_1532
		), .Z(n_263788538));
	notech_ao4 i_182147972(.A(n_33118), .B(n_30191), .C(n_338361011), .D(n_30196
		), .Z(n_263988540));
	notech_and4 i_182547968(.A(n_65022753), .B(n_263988540), .C(n_263788538)
		, .D(n_260088501), .Z(n_264188542));
	notech_ao4 i_181847975(.A(n_443768021), .B(n_58384), .C(n_443868022), .D
		(n_58866), .Z(n_264288543));
	notech_ao4 i_181747976(.A(n_444068024), .B(n_232870324), .C(n_57130), .D
		(n_305478064), .Z(n_264488545));
	notech_nand3 i_182047973(.A(n_264288543), .B(n_264488545), .C(n_259588496
		), .Z(n_264588546));
	notech_ao4 i_181547978(.A(n_119226519), .B(n_33202), .C(n_5356), .D(n_119326520
		), .Z(n_264688547));
	notech_ao4 i_181147982(.A(n_443768021), .B(n_58375), .C(n_443868022), .D
		(n_59077), .Z(n_264988550));
	notech_ao4 i_181047983(.A(n_444068024), .B(n_235370349), .C(n_57130), .D
		(n_265785074), .Z(n_265188552));
	notech_nand3 i_181347980(.A(n_264988550), .B(n_265188552), .C(n_258788488
		), .Z(n_265288553));
	notech_ao4 i_180847985(.A(n_119226519), .B(n_33201), .C(n_5436), .D(n_119326520
		), .Z(n_265388554));
	notech_ao4 i_180447989(.A(n_443768021), .B(n_58366), .C(n_443868022), .D
		(n_59086), .Z(n_265688557));
	notech_ao4 i_180347990(.A(n_237870374), .B(n_444068024), .C(n_57130), .D
		(n_266585082), .Z(n_265888559));
	notech_nand3 i_180647987(.A(n_265688557), .B(n_265888559), .C(n_257988480
		), .Z(n_265988560));
	notech_ao4 i_180147992(.A(n_119226519), .B(n_33200), .C(n_5397), .D(n_119326520
		), .Z(n_266088561));
	notech_ao4 i_179747996(.A(n_443768021), .B(n_58357), .C(n_443868022), .D
		(n_59059), .Z(n_266388564));
	notech_ao4 i_179647997(.A(n_444068024), .B(n_240370399), .C(n_267385090)
		, .D(n_57130), .Z(n_266588566));
	notech_nand3 i_179947994(.A(n_266388564), .B(n_266588566), .C(n_257188472
		), .Z(n_266688567));
	notech_ao4 i_179447999(.A(n_119226519), .B(n_33199), .C(n_5444), .D(n_119326520
		), .Z(n_266788568));
	notech_ao4 i_179048003(.A(n_74922852), .B(n_376764298), .C(n_66222765), 
		.D(n_57130), .Z(n_267088571));
	notech_ao4 i_178948004(.A(n_75322856), .B(n_29680), .C(n_75222855), .D(n_29681
		), .Z(n_267188572));
	notech_ao4 i_178748006(.A(n_75522858), .B(n_29677), .C(n_75622859), .D(n_29678
		), .Z(n_267388574));
	notech_and4 i_179248001(.A(n_267388574), .B(n_267188572), .C(n_267088571
		), .D(n_255988460), .Z(n_267588576));
	notech_ao4 i_178448009(.A(n_74522848), .B(n_376664297), .C(n_74622849), 
		.D(n_94542386), .Z(n_267688577));
	notech_ao4 i_178248011(.A(n_33118), .B(n_376964300), .C(n_338361011), .D
		(n_376864299), .Z(n_267888579));
	notech_and4 i_178648007(.A(n_267888579), .B(n_267688577), .C(n_65022753)
		, .D(n_255688457), .Z(n_268088581));
	notech_ao4 i_177948014(.A(n_319725273), .B(n_303822063), .C(n_232870324)
		, .D(n_299122016), .Z(n_268188582));
	notech_ao4 i_177848015(.A(n_5356), .B(n_57320), .C(n_57319), .D(n_33202)
		, .Z(n_268388584));
	notech_and3 i_178148012(.A(n_268188582), .B(n_268388584), .C(n_255188452
		), .Z(n_268488585));
	notech_ao4 i_177648017(.A(n_57363), .B(n_58384), .C(n_57362), .D(n_58866
		), .Z(n_268588586));
	notech_ao4 i_177548018(.A(n_31527), .B(n_61697), .C(n_303922064), .D(n_60483
		), .Z(n_268688587));
	notech_ao4 i_177248021(.A(n_319825274), .B(n_303822063), .C(n_235370349)
		, .D(n_299122016), .Z(n_268888589));
	notech_ao4 i_177148022(.A(n_5436), .B(n_57320), .C(n_57319), .D(n_33201)
		, .Z(n_269088591));
	notech_and3 i_177448019(.A(n_268888589), .B(n_269088591), .C(n_254388444
		), .Z(n_269188592));
	notech_ao4 i_176948024(.A(n_57363), .B(n_58375), .C(n_57362), .D(n_59077
		), .Z(n_269288593));
	notech_ao4 i_176848025(.A(n_31526), .B(n_61698), .C(n_303922064), .D(nbus_11271
		[18]), .Z(n_269388594));
	notech_ao4 i_176548028(.A(n_319951172), .B(n_303822063), .C(n_237870374)
		, .D(n_299122016), .Z(n_269588596));
	notech_ao4 i_176448029(.A(n_5397), .B(n_57320), .C(n_57319), .D(n_33200)
		, .Z(n_269788598));
	notech_and3 i_176748026(.A(n_269588596), .B(n_269788598), .C(n_253588436
		), .Z(n_269888599));
	notech_ao4 i_176248031(.A(n_57363), .B(n_58366), .C(n_57362), .D(n_59086
		), .Z(n_269988600));
	notech_ao4 i_176148032(.A(n_31525), .B(n_61698), .C(n_303922064), .D(n_60501
		), .Z(n_270088601));
	notech_ao4 i_175848035(.A(n_320051171), .B(n_303822063), .C(n_240370399)
		, .D(n_299122016), .Z(n_270288603));
	notech_ao4 i_175748036(.A(n_5444), .B(n_57320), .C(n_57319), .D(n_33199)
		, .Z(n_270488605));
	notech_and3 i_176048033(.A(n_270288603), .B(n_270488605), .C(n_252788428
		), .Z(n_270588606));
	notech_ao4 i_175548038(.A(n_57363), .B(n_58357), .C(n_57362), .D(n_59059
		), .Z(n_270688607));
	notech_ao4 i_175448039(.A(n_31524), .B(n_61698), .C(n_303922064), .D(n_60474
		), .Z(n_270788608));
	notech_ao4 i_169248101(.A(n_319825274), .B(n_28852), .C(n_235370349), .D
		(n_28869), .Z(n_270988610));
	notech_ao4 i_169148102(.A(n_5436), .B(n_388264413), .C(n_388364414), .D(n_33201
		), .Z(n_271188612));
	notech_nand3 i_169448099(.A(n_270988610), .B(n_271188612), .C(n_251988420
		), .Z(n_271288613));
	notech_ao4 i_168948104(.A(n_28874), .B(n_58375), .C(n_28863), .D(n_59077
		), .Z(n_271388614));
	notech_ao4 i_168548108(.A(n_319951172), .B(n_28852), .C(n_237870374), .D
		(n_28869), .Z(n_271688617));
	notech_ao4 i_168448109(.A(n_5397), .B(n_388264413), .C(n_33200), .D(n_388364414
		), .Z(n_271888619));
	notech_nand3 i_168748106(.A(n_271688617), .B(n_271888619), .C(n_251188412
		), .Z(n_271988620));
	notech_ao4 i_168248111(.A(n_28874), .B(n_58366), .C(n_28863), .D(n_59086
		), .Z(n_272088621));
	notech_ao4 i_167848115(.A(n_320051171), .B(n_28852), .C(n_240370399), .D
		(n_28869), .Z(n_272388624));
	notech_ao4 i_167748116(.A(n_5444), .B(n_388264413), .C(n_388364414), .D(n_33199
		), .Z(n_272588626));
	notech_nand3 i_168048113(.A(n_272388624), .B(n_272588626), .C(n_250388404
		), .Z(n_272688627));
	notech_ao4 i_167548118(.A(n_28874), .B(n_58357), .C(n_28863), .D(n_59059
		), .Z(n_272788628));
	notech_or4 i_4446368(.A(n_58561), .B(n_365964190), .C(n_23760), .D(n_5269
		), .Z(n_273488635));
	notech_or2 i_4146371(.A(n_386164392), .B(\nbus_11290[8] ), .Z(n_273788638
		));
	notech_or4 i_37646042(.A(n_58592), .B(n_384764378), .C(n_384964380), .D(n_5269
		), .Z(n_274688647));
	notech_nand2 i_37346045(.A(n_30354), .B(opd[8]), .Z(n_274988650));
	notech_or4 i_37046048(.A(n_63706), .B(n_440667990), .C(n_63794), .D(nbus_11273
		[8]), .Z(n_275288653));
	notech_or2 i_44645975(.A(n_26935), .B(n_33253), .Z(n_275388654));
	notech_or4 i_44545976(.A(n_162262654), .B(n_26951), .C(n_5269), .D(n_57401
		), .Z(n_275788657));
	notech_nand2 i_44145979(.A(opd[8]), .B(n_305144485), .Z(n_276088660));
	notech_or4 i_43745982(.A(n_63706), .B(n_303844472), .C(n_63794), .D(nbus_11273
		[8]), .Z(n_276388663));
	notech_or2 i_50345929(.A(n_57252), .B(n_33253), .Z(n_276688666));
	notech_or2 i_50045932(.A(n_57110), .B(nbus_11273[8]), .Z(n_276988669));
	notech_or2 i_49745935(.A(n_56896), .B(n_33315), .Z(n_277288672));
	notech_or4 i_49445938(.A(n_63706), .B(n_57388), .C(n_63794), .D(nbus_11273
		[8]), .Z(n_277588675));
	notech_or2 i_55145882(.A(n_28855), .B(n_33253), .Z(n_277688676));
	notech_or4 i_55045883(.A(n_57476), .B(n_3298), .C(n_3290), .D(n_5269), .Z
		(n_277988679));
	notech_nand2 i_54745886(.A(opd[8]), .B(n_305044484), .Z(n_278288682));
	notech_or4 i_54445889(.A(n_63706), .B(n_303744471), .C(n_63778), .D(n_58285
		), .Z(n_278588685));
	notech_nor2 i_57945854(.A(n_5243), .B(n_388264413), .Z(n_278688686));
	notech_nao3 i_57445859(.A(n_57382), .B(opd[31]), .C(n_57187), .Z(n_279388693
		));
	notech_nao3 i_58845845(.A(n_30300), .B(\opa_12[8] ), .C(n_376064291), .Z
		(n_279888698));
	notech_or2 i_58545848(.A(n_58029), .B(n_31481), .Z(n_280188701));
	notech_or4 i_58245851(.A(n_63706), .B(n_57387), .C(n_63778), .D(n_58285)
		, .Z(n_280488704));
	notech_nao3 i_61145825(.A(n_30282), .B(\opa_12[8] ), .C(n_386964400), .Z
		(n_280588705));
	notech_or4 i_61045826(.A(n_57467), .B(n_286263764), .C(n_29560), .D(n_5269
		), .Z(n_280888708));
	notech_or2 i_60745829(.A(n_445268036), .B(n_31481), .Z(n_281188711));
	notech_or4 i_60345832(.A(n_63706), .B(n_445168035), .C(n_63778), .D(n_58285
		), .Z(n_281488714));
	notech_or2 i_61545822(.A(n_303922064), .B(n_60591), .Z(n_282288722));
	notech_or2 i_63045807(.A(n_62642067), .B(n_58285), .Z(n_282388723));
	notech_or2 i_62945808(.A(n_62742068), .B(n_59014), .Z(n_282688726));
	notech_or2 i_62645811(.A(n_446068044), .B(n_33253), .Z(n_282988729));
	notech_or4 i_62345814(.A(n_63706), .B(n_62442065), .C(n_63778), .D(n_58285
		), .Z(n_283288732));
	notech_nor2 i_63845799(.A(n_443668020), .B(n_60591), .Z(n_283388733));
	notech_and3 i_63345804(.A(n_57382), .B(n_32224), .C(opd[31]), .Z(n_284088740
		));
	notech_ao4 i_170944804(.A(n_443968023), .B(n_300822033), .C(n_444068024)
		, .D(n_262470619), .Z(n_284188741));
	notech_ao4 i_170844805(.A(n_5243), .B(n_119326520), .C(n_119226519), .D(n_33206
		), .Z(n_284388743));
	notech_nao3 i_171144802(.A(n_284188741), .B(n_284388743), .C(n_284088740
		), .Z(n_284488744));
	notech_ao4 i_170644807(.A(n_443768021), .B(n_60458), .C(n_443868022), .D
		(n_58983), .Z(n_284588745));
	notech_ao4 i_170244811(.A(n_266870661), .B(n_30601), .C(n_4418), .D(n_266970662
		), .Z(n_284888748));
	notech_ao4 i_170044813(.A(n_267170664), .B(n_442182452), .C(n_335678362)
		, .D(n_57130), .Z(n_285088750));
	notech_and4 i_170444809(.A(n_285088750), .B(n_284888748), .C(n_282988729
		), .D(n_283288732), .Z(n_285288752));
	notech_ao4 i_169744816(.A(n_62142062), .B(n_31481), .C(n_5269), .D(n_445968043
		), .Z(n_285388753));
	notech_and4 i_169944814(.A(n_336078366), .B(n_285388753), .C(n_282388723
		), .D(n_282688726), .Z(n_285688756));
	notech_ao4 i_169344820(.A(n_300822033), .B(n_303822063), .C(n_262470619)
		, .D(n_299122016), .Z(n_285788757));
	notech_ao4 i_169244821(.A(n_57362), .B(n_58983), .C(n_57363), .D(\nbus_11283[31] 
		), .Z(n_285988759));
	notech_and3 i_169544818(.A(n_285788757), .B(n_285988759), .C(n_282288722
		), .Z(n_286088760));
	notech_ao4 i_169044823(.A(n_57319), .B(n_33206), .C(n_5243), .D(n_57320)
		, .Z(n_286188761));
	notech_ao4 i_168944824(.A(n_31539), .B(n_61697), .C(n_386864399), .D(n_31507
		), .Z(n_286288762));
	notech_ao4 i_168644827(.A(n_266870661), .B(n_30599), .C(n_29418), .D(n_266970662
		), .Z(n_286488764));
	notech_ao4 i_168444829(.A(n_267170664), .B(n_29416), .C(n_57059), .D(n_335678362
		), .Z(n_286688766));
	notech_and4 i_168844825(.A(n_286688766), .B(n_286488764), .C(n_281188711
		), .D(n_281488714), .Z(n_286888768));
	notech_ao4 i_168144832(.A(n_444968033), .B(n_59014), .C(n_445068034), .D
		(n_58285), .Z(n_286988769));
	notech_and4 i_168344830(.A(n_336078366), .B(n_280888708), .C(n_286988769
		), .D(n_280588705), .Z(n_287288772));
	notech_ao4 i_167044843(.A(n_334478350), .B(n_266870661), .C(n_334378349)
		, .D(n_266970662), .Z(n_287388773));
	notech_ao4 i_166844845(.A(n_334578351), .B(n_267170664), .C(n_57604), .D
		(n_335678362), .Z(n_287588775));
	notech_and4 i_167244841(.A(n_287588775), .B(n_287388773), .C(n_280188701
		), .D(n_280488704), .Z(n_287788777));
	notech_ao4 i_166544848(.A(n_57237), .B(n_58285), .C(n_57238), .D(n_59014
		), .Z(n_287888778));
	notech_ao4 i_166344850(.A(n_279977810), .B(nbus_11271[8]), .C(n_323378242
		), .D(n_5269), .Z(n_288088780));
	notech_and4 i_166744846(.A(n_336078366), .B(n_288088780), .C(n_287888778
		), .D(n_279888698), .Z(n_288288782));
	notech_ao4 i_166044853(.A(n_300822033), .B(n_28852), .C(n_262470619), .D
		(n_28869), .Z(n_288388783));
	notech_ao4 i_165944854(.A(n_28867), .B(n_60591), .C(n_28863), .D(n_58983
		), .Z(n_288588785));
	notech_nand3 i_166244851(.A(n_288388783), .B(n_288588785), .C(n_279388693
		), .Z(n_288688786));
	notech_ao4 i_165744856(.A(n_388364414), .B(n_33206), .C(n_28874), .D(n_60458
		), .Z(n_288788787));
	notech_ao4 i_157644933(.A(n_28742), .B(n_266870661), .C(n_28743), .D(n_266970662
		), .Z(n_289088790));
	notech_ao4 i_157444935(.A(n_267170664), .B(n_28741), .C(n_57187), .D(n_335678362
		), .Z(n_289288792));
	notech_and4 i_157944931(.A(n_289288792), .B(n_289088790), .C(n_278288682
		), .D(n_278588685), .Z(n_289488794));
	notech_ao4 i_157144938(.A(n_59014), .B(n_303044464), .C(n_302944463), .D
		(n_58285), .Z(n_289588795));
	notech_and4 i_157344936(.A(n_336078366), .B(n_277988679), .C(n_289588795
		), .D(n_277688676), .Z(n_289888798));
	notech_ao4 i_153644972(.A(n_200777063), .B(n_266870661), .C(n_200677062)
		, .D(n_266970662), .Z(n_289988799));
	notech_ao4 i_153444974(.A(n_267170664), .B(n_200577061), .C(n_57152), .D
		(n_335678362), .Z(n_290188801));
	notech_and4 i_153844970(.A(n_290188801), .B(n_289988799), .C(n_277288672
		), .D(n_277588675), .Z(n_290388803));
	notech_ao4 i_153144977(.A(n_58053), .B(n_31481), .C(n_56783), .D(n_31516
		), .Z(n_290488804));
	notech_ao4 i_152944979(.A(n_5269), .B(n_57317), .C(n_57133), .D(n_59014)
		, .Z(n_290688806));
	notech_and4 i_153344975(.A(n_290688806), .B(n_290488804), .C(n_276688666
		), .D(n_276988669), .Z(n_290888808));
	notech_ao4 i_149545011(.A(n_266870661), .B(n_30593), .C(n_266970662), .D
		(n_30592), .Z(n_290988809));
	notech_ao4 i_149345013(.A(n_267170664), .B(n_26821), .C(n_57081), .D(n_335678362
		), .Z(n_291188811));
	notech_and4 i_149745009(.A(n_291188811), .B(n_290988809), .C(n_276088660
		), .D(n_276388663), .Z(n_291388813));
	notech_ao4 i_149045016(.A(n_59014), .B(n_303244466), .C(n_58285), .D(n_303144465
		), .Z(n_291488814));
	notech_and4 i_149245014(.A(n_336078366), .B(n_275788657), .C(n_291488814
		), .D(n_275388654), .Z(n_291788817));
	notech_ao4 i_142945069(.A(n_4533), .B(n_266870661), .C(n_441868002), .D(n_266970662
		), .Z(n_291888818));
	notech_ao4 i_142745071(.A(n_385464385), .B(n_267170664), .C(n_335678362)
		, .D(n_57174), .Z(n_292088820));
	notech_and4 i_143745067(.A(n_292088820), .B(n_291888818), .C(n_274988650
		), .D(n_275288653), .Z(n_292288822));
	notech_ao4 i_142245074(.A(n_441668000), .B(n_59014), .C(n_441768001), .D
		(n_58285), .Z(n_292388823));
	notech_ao4 i_142045076(.A(n_56035), .B(n_32560), .C(n_385664387), .D(n_33253
		), .Z(n_292588825));
	notech_and4 i_142645072(.A(n_336078366), .B(n_292588825), .C(n_274688647
		), .D(n_292388823), .Z(n_292788827));
	notech_ao4 i_109845361(.A(n_266870661), .B(n_23614), .C(n_266970662), .D
		(n_23613), .Z(n_292888828));
	notech_ao4 i_109745362(.A(n_335678362), .B(n_58696), .C(n_386364394), .D
		(n_267470667), .Z(n_292988829));
	notech_ao4 i_109545364(.A(n_386264393), .B(n_31481), .C(n_267170664), .D
		(n_23611), .Z(n_293188831));
	notech_and4 i_110045359(.A(n_293188831), .B(n_292988829), .C(n_292888828
		), .D(n_273788638), .Z(n_293388833));
	notech_ao4 i_109245367(.A(n_23747), .B(n_33253), .C(n_386064391), .D(n_58285
		), .Z(n_293488834));
	notech_ao4 i_109045369(.A(n_56035), .B(n_32537), .C(n_58664), .D(nbus_11271
		[8]), .Z(n_293688836));
	notech_and4 i_109445365(.A(n_293688836), .B(n_273488635), .C(n_293488834
		), .D(n_336078366), .Z(n_293888838));
	notech_and2 i_2043257(.A(n_322089108), .B(n_58116456), .Z(n_293988839)
		);
	notech_and2 i_12343166(.A(n_57622), .B(n_57489), .Z(n_294088840));
	notech_and2 i_1943258(.A(n_56823), .B(n_294288842), .Z(n_294188841));
	notech_or2 i_22843062(.A(n_61816493), .B(n_57467), .Z(n_294288842));
	notech_or2 i_37342917(.A(n_61516490), .B(n_59068), .Z(n_294388843));
	notech_or2 i_6943217(.A(n_56891), .B(n_58238), .Z(n_294988849));
	notech_or4 i_6643220(.A(n_4025), .B(n_60169), .C(n_61607), .D(n_56965), 
		.Z(n_295288852));
	notech_or2 i_6343223(.A(n_56850), .B(nbus_11271[0]), .Z(n_295588855));
	notech_nao3 i_6043226(.A(n_27843), .B(nbus_137[0]), .C(n_56871), .Z(n_295888858
		));
	notech_nao3 i_5743229(.A(n_405982375), .B(imm[32]), .C(n_25713), .Z(n_296188861
		));
	notech_nand2 i_5443232(.A(read_data[8]), .B(n_26316138), .Z(n_296488864)
		);
	notech_nao3 i_5143235(.A(imm[0]), .B(n_382682257), .C(n_61816493), .Z(n_296788867
		));
	notech_or2 i_9443193(.A(n_56891), .B(n_58229), .Z(n_297288872));
	notech_or4 i_9143196(.A(n_4025), .B(n_60169), .C(n_61607), .D(n_56956), 
		.Z(n_297588875));
	notech_or2 i_8843199(.A(n_56850), .B(nbus_11271[1]), .Z(n_297888878));
	notech_nao3 i_8543202(.A(n_58532), .B(nbus_137[1]), .C(n_56871), .Z(n_298188881
		));
	notech_nao3 i_8243205(.A(n_405982375), .B(imm[33]), .C(n_25713), .Z(n_298488884
		));
	notech_nand2 i_7943208(.A(read_data[9]), .B(n_26316138), .Z(n_298788887)
		);
	notech_or2 i_204143267(.A(n_32305), .B(n_61816493), .Z(n_299488894));
	notech_or2 i_12043169(.A(n_56891), .B(nbus_11273[2]), .Z(n_299788897));
	notech_or4 i_11743172(.A(n_4025), .B(n_60163), .C(n_61607), .D(n_58802),
		 .Z(n_300088900));
	notech_or2 i_11443175(.A(n_56850), .B(nbus_11271[2]), .Z(n_300388903));
	notech_nao3 i_11043178(.A(n_58532), .B(nbus_137[2]), .C(n_56871), .Z(n_300788906
		));
	notech_nao3 i_10643181(.A(imm[34]), .B(n_405982375), .C(n_25713), .Z(n_301088909
		));
	notech_nand2 i_10343184(.A(read_data[10]), .B(n_26316138), .Z(n_301388912
		));
	notech_or4 i_16543124(.A(n_340561033), .B(n_32627), .C(n_61607), .D(nbus_11271
		[12]), .Z(n_301888917));
	notech_nand2 i_16443125(.A(resb_shiftbox[4]), .B(n_30417), .Z(n_302188920
		));
	notech_or4 i_16143128(.A(n_4025), .B(n_60163), .C(n_61607), .D(n_56974),
		 .Z(n_302488923));
	notech_or2 i_15843131(.A(n_56850), .B(nbus_11271[4]), .Z(n_302788926));
	notech_or2 i_15343136(.A(n_61516490), .B(n_59050), .Z(n_303388931));
	notech_nand2 i_15043139(.A(read_data[28]), .B(n_26116136), .Z(n_303688934
		));
	notech_nand2 i_14743142(.A(add_src[4]), .B(n_30416), .Z(n_303988937));
	notech_or4 i_18543104(.A(n_58610), .B(n_32627), .C(n_61607), .D(nbus_11271
		[13]), .Z(n_304088938));
	notech_nand2 i_18443105(.A(resb_shiftbox[5]), .B(n_30417), .Z(n_304388941
		));
	notech_nao3 i_17943110(.A(resb_shift4box[5]), .B(n_396382340), .C(n_25670
		), .Z(n_304988946));
	notech_or4 i_17443115(.A(n_32397), .B(n_25485), .C(n_61607), .D(n_31494)
		, .Z(n_305488951));
	notech_nand2 i_17143118(.A(read_data[5]), .B(n_30415), .Z(n_305788954)
		);
	notech_or2 i_16843121(.A(n_26716142), .B(n_31529), .Z(n_306188957));
	notech_or4 i_20643084(.A(n_58610), .B(n_32627), .C(n_61607), .D(nbus_11271
		[14]), .Z(n_306288958));
	notech_nand2 i_20543085(.A(resb_shiftbox[6]), .B(n_30417), .Z(n_306588961
		));
	notech_nao3 i_19943090(.A(resb_shift4box[6]), .B(n_396382340), .C(n_25670
		), .Z(n_307088966));
	notech_or2 i_19443095(.A(n_40216277), .B(n_31496), .Z(n_307588971));
	notech_nand2 i_19143098(.A(read_data[6]), .B(n_30415), .Z(n_307988974)
		);
	notech_or2 i_18843101(.A(n_26716142), .B(n_31530), .Z(n_308288977));
	notech_or4 i_22743063(.A(n_58610), .B(n_32627), .C(n_61607), .D(nbus_11271
		[15]), .Z(n_308388978));
	notech_nand2 i_22643064(.A(resb_shiftbox[7]), .B(n_30417), .Z(n_308688981
		));
	notech_nao3 i_22143069(.A(resb_shift4box[7]), .B(n_396382340), .C(n_25670
		), .Z(n_309188986));
	notech_nor2 i_21643074(.A(n_40216277), .B(n_31499), .Z(n_309788991));
	notech_or2 i_21143079(.A(n_26716142), .B(n_31531), .Z(n_310288996));
	notech_or4 i_24943041(.A(n_28098), .B(n_58610), .C(n_61607), .D(nbus_11271
		[0]), .Z(n_310388997));
	notech_or2 i_24443046(.A(n_60316478), .B(n_31481), .Z(n_311189004));
	notech_nand2 i_23543055(.A(add_src[8]), .B(n_30416), .Z(n_312189013));
	notech_and2 i_180243277(.A(n_446968053), .B(n_294388843), .Z(n_312289014
		));
	notech_ao4 i_140141941(.A(n_56823), .B(n_32312), .C(n_56841), .D(n_31516
		), .Z(n_312389015));
	notech_ao4 i_140041942(.A(n_40616281), .B(n_32309), .C(n_443982453), .D(n_59014
		), .Z(n_312589017));
	notech_and3 i_140441939(.A(n_312389015), .B(n_312589017), .C(n_312189013
		), .Z(n_312689018));
	notech_ao4 i_139841944(.A(n_40116276), .B(n_32873), .C(n_31500), .D(n_40216277
		), .Z(n_312789019));
	notech_ao4 i_139741945(.A(n_56850), .B(nbus_11271[8]), .C(n_40316278), .D
		(n_32711), .Z(n_312889020));
	notech_ao4 i_139241949(.A(n_61116486), .B(n_33144), .C(n_56861), .D(n_32205
		), .Z(n_313189023));
	notech_ao4 i_139141950(.A(n_56891), .B(n_58285), .C(n_56880), .D(n_5269)
		, .Z(n_313389025));
	notech_ao4 i_138941952(.A(n_56929), .B(\nbus_11290[24] ), .C(n_56904), .D
		(n_32165), .Z(n_313589027));
	notech_and4 i_139041951(.A(n_446968053), .B(n_313589027), .C(n_382982260
		), .D(n_310388997), .Z(n_313789029));
	notech_and4 i_139541946(.A(n_313189023), .B(n_313389025), .C(n_311189004
		), .D(n_313789029), .Z(n_313889030));
	notech_ao4 i_137741964(.A(n_56832), .B(n_32325), .C(n_294188841), .D(n_32265
		), .Z(n_313989031));
	notech_ao4 i_137641965(.A(n_30606), .B(n_31539), .C(n_30605), .D(n_31523
		), .Z(n_314189033));
	notech_ao4 i_137341968(.A(n_40616281), .B(n_32307), .C(n_4434), .D(n_31515
		), .Z(n_314389035));
	notech_ao4 i_137241969(.A(n_40316278), .B(n_32710), .C(n_40116276), .D(n_32872
		), .Z(n_314689037));
	notech_ao3 i_137541966(.A(n_314389035), .B(n_314689037), .C(n_309788991)
		, .Z(n_314789038));
	notech_and4 i_138041961(.A(n_313989031), .B(n_314189033), .C(n_310288996
		), .D(n_314789038), .Z(n_314889039));
	notech_ao4 i_136841973(.A(n_56850), .B(nbus_11271[7]), .C(n_4433), .D(\nbus_11290[7] 
		), .Z(n_314989040));
	notech_ao4 i_136741974(.A(n_56914), .B(n_31480), .C(n_61116486), .D(n_32154
		), .Z(n_315189042));
	notech_and3 i_137041971(.A(n_314989040), .B(n_315189042), .C(n_309188986
		), .Z(n_315289043));
	notech_ao4 i_136441977(.A(n_56891), .B(nbus_11273[7]), .C(n_100242443), 
		.D(n_56880), .Z(n_315389044));
	notech_and4 i_136641975(.A(n_315389044), .B(n_312289014), .C(n_308388978
		), .D(n_308688981), .Z(n_315689047));
	notech_ao4 i_135841983(.A(n_56832), .B(n_32324), .C(n_23916114), .D(n_32276
		), .Z(n_315889049));
	notech_ao4 i_135641985(.A(n_31538), .B(n_30606), .C(n_30605), .D(n_31522
		), .Z(n_316089051));
	notech_and4 i_136041981(.A(n_316089051), .B(n_315889049), .C(n_307988974
		), .D(n_308288977), .Z(n_316289053));
	notech_ao4 i_135341988(.A(n_61516490), .B(n_59041), .C(n_40616281), .D(n_32306
		), .Z(n_316389054));
	notech_ao4 i_135241989(.A(n_40316278), .B(n_32709), .C(n_40116276), .D(n_32871
		), .Z(n_316589056));
	notech_and4 i_136141980(.A(n_316389054), .B(n_316589056), .C(n_316289053
		), .D(n_307588971), .Z(n_316789058));
	notech_ao4 i_134841993(.A(n_56850), .B(nbus_11271[6]), .C(n_4433), .D(\nbus_11290[6] 
		), .Z(n_316989059));
	notech_ao4 i_134741994(.A(n_56914), .B(n_31479), .C(n_61116486), .D(n_32153
		), .Z(n_317189061));
	notech_and3 i_135041991(.A(n_316989059), .B(n_317189061), .C(n_307088966
		), .Z(n_317289062));
	notech_ao4 i_134441997(.A(n_56891), .B(n_58265), .C(n_100542446), .D(n_56880
		), .Z(n_317389063));
	notech_and4 i_134641995(.A(n_22216097), .B(n_317389063), .C(n_306288958)
		, .D(n_306588961), .Z(n_317689066));
	notech_ao4 i_133942002(.A(n_56832), .B(n_32322), .C(n_23916114), .D(n_32274
		), .Z(n_317889068));
	notech_ao4 i_133742004(.A(n_30606), .B(n_31537), .C(n_30605), .D(n_31521
		), .Z(n_318089070));
	notech_and4 i_134142000(.A(n_318089070), .B(n_317889068), .C(n_305788954
		), .D(n_306188957), .Z(n_318289072));
	notech_ao4 i_133442007(.A(n_61516490), .B(\nbus_11290[13] ), .C(n_40616281
		), .D(n_32303), .Z(n_318389073));
	notech_ao4 i_133342008(.A(n_40316278), .B(n_32708), .C(n_40116276), .D(n_32870
		), .Z(n_318589075));
	notech_and4 i_134241999(.A(n_318389073), .B(n_318589075), .C(n_318289072
		), .D(n_305488951), .Z(n_318789077));
	notech_ao4 i_132942012(.A(n_56850), .B(nbus_11271[5]), .C(n_4433), .D(\nbus_11290[5] 
		), .Z(n_318989078));
	notech_ao4 i_132842013(.A(n_56914), .B(n_56983), .C(n_61116486), .D(n_32152
		), .Z(n_319189080));
	notech_and3 i_133142010(.A(n_318989078), .B(n_319189080), .C(n_304988946
		), .Z(n_319289081));
	notech_ao4 i_132542016(.A(n_56891), .B(nbus_11273[5]), .C(n_334860976), 
		.D(n_56880), .Z(n_319389082));
	notech_and4 i_132742014(.A(n_22216097), .B(n_319389082), .C(n_304388941)
		, .D(n_304088938), .Z(n_319689085));
	notech_or4 i_132342018(.A(opz[0]), .B(opz[1]), .C(n_31606), .D(n_57444),
		 .Z(n_319889087));
	notech_ao4 i_131942022(.A(n_23916114), .B(n_32300), .C(n_61816493), .D(n_319889087
		), .Z(n_319989088));
	notech_ao4 i_131742024(.A(n_31520), .B(n_30605), .C(n_31528), .D(n_26716142
		), .Z(n_320189090));
	notech_and4 i_132142020(.A(n_320189090), .B(n_319989088), .C(n_303988937
		), .D(n_303688934), .Z(n_320489092));
	notech_ao4 i_131442027(.A(n_40616281), .B(n_32301), .C(n_4434), .D(n_31512
		), .Z(n_320589093));
	notech_ao4 i_131342028(.A(n_40116276), .B(n_32869), .C(n_40216277), .D(n_31493
		), .Z(n_320789095));
	notech_and4 i_132242019(.A(n_320589093), .B(n_320789095), .C(n_320489092
		), .D(n_303388931), .Z(n_320989097));
	notech_ao4 i_130942032(.A(n_4433), .B(\nbus_11290[4] ), .C(n_40316278), 
		.D(n_32707), .Z(n_321089098));
	notech_ao4 i_130742034(.A(n_61116486), .B(n_32151), .C(n_56861), .D(n_32202
		), .Z(n_321289100));
	notech_and4 i_131142030(.A(n_321289100), .B(n_321089098), .C(n_302488923
		), .D(n_302788926), .Z(n_321489102));
	notech_ao4 i_130442037(.A(n_56891), .B(nbus_11273[4]), .C(n_56880), .D(n_334660974
		), .Z(n_321589103));
	notech_and4 i_130642035(.A(n_22216097), .B(n_321589103), .C(n_302188920)
		, .D(n_301888917), .Z(n_321889106));
	notech_or4 i_202343268(.A(instrc[123]), .B(instrc[121]), .C(n_32250), .D
		(n_61816493), .Z(n_322089108));
	notech_or2 i_196043270(.A(n_61816493), .B(n_294088840), .Z(n_322189109)
		);
	notech_ao4 i_127842063(.A(n_322189109), .B(n_33164), .C(n_322089108), .D
		(n_31606), .Z(n_322289110));
	notech_ao4 i_127742064(.A(n_58116456), .B(n_56898), .C(n_23916114), .D(n_32271
		), .Z(n_322389111));
	notech_ao4 i_127542066(.A(n_26716142), .B(n_31526), .C(n_56832), .D(n_32318
		), .Z(n_322589113));
	notech_and4 i_128042061(.A(n_322589113), .B(n_322389111), .C(n_322289110
		), .D(n_301388912), .Z(n_322789115));
	notech_ao4 i_127242069(.A(n_4434), .B(n_31510), .C(n_30606), .D(n_31534)
		, .Z(n_322889116));
	notech_ao4 i_127042071(.A(n_40216277), .B(n_31491), .C(n_61516490), .D(\nbus_11290[10] 
		), .Z(n_323089118));
	notech_and4 i_127442067(.A(n_323089118), .B(n_322889116), .C(n_300788906
		), .D(n_301088909), .Z(n_323289120));
	notech_ao4 i_126642075(.A(n_4433), .B(\nbus_11290[2] ), .C(n_40316278), 
		.D(n_32705), .Z(n_323489122));
	notech_ao4 i_126442077(.A(n_61116486), .B(n_32149), .C(n_56861), .D(n_32200
		), .Z(n_323689124));
	notech_and4 i_126842073(.A(n_323689124), .B(n_323489122), .C(n_300088900
		), .D(n_300388903), .Z(n_323889126));
	notech_ao4 i_126142080(.A(n_57401), .B(n_61816493), .C(n_100842449), .D(n_56880
		), .Z(n_323989127));
	notech_ao4 i_125942082(.A(n_56929), .B(nbus_11271[10]), .C(n_4437), .D(n_32164
		), .Z(n_324189129));
	notech_and4 i_126342078(.A(n_299488894), .B(n_324189129), .C(n_323989127
		), .D(n_299788897), .Z(n_324389131));
	notech_ao4 i_125542086(.A(n_322189109), .B(n_33156), .C(n_322089108), .D
		(n_31605), .Z(n_324589133));
	notech_ao4 i_125442087(.A(n_58116456), .B(n_57104), .C(n_23916114), .D(n_32270
		), .Z(n_324689134));
	notech_ao4 i_125242089(.A(n_26716142), .B(n_31525), .C(n_56832), .D(n_32316
		), .Z(n_324889136));
	notech_and4 i_125742084(.A(n_324889136), .B(n_324689134), .C(n_324589133
		), .D(n_298788887), .Z(n_325089138));
	notech_ao4 i_124942092(.A(n_4434), .B(n_31509), .C(n_30606), .D(n_31533)
		, .Z(n_325189139));
	notech_ao4 i_124742094(.A(n_40216277), .B(n_31490), .C(n_61516490), .D(n_59032
		), .Z(n_325389141));
	notech_and4 i_125142090(.A(n_325389141), .B(n_325189139), .C(n_298188881
		), .D(n_298488884), .Z(n_325589143));
	notech_ao4 i_124342098(.A(n_4433), .B(n_59001), .C(n_40316278), .D(n_32704
		), .Z(n_325789145));
	notech_ao4 i_124142100(.A(n_61116486), .B(n_32148), .C(n_56861), .D(n_32198
		), .Z(n_325989147));
	notech_and4 i_124542096(.A(n_325989147), .B(n_325789145), .C(n_297588875
		), .D(n_297888878), .Z(n_326189149));
	notech_ao4 i_123842103(.A(n_57436), .B(n_61816493), .C(n_334360971), .D(n_56880
		), .Z(n_326289150));
	notech_ao4 i_123642105(.A(n_56929), .B(nbus_11271[9]), .C(n_56904), .D(n_32163
		), .Z(n_326489152));
	notech_and4 i_124042101(.A(n_326489152), .B(n_326289150), .C(n_299488894
		), .D(n_297288872), .Z(n_326689154));
	notech_ao4 i_123242109(.A(n_322189109), .B(n_33174), .C(n_293988839), .D
		(n_31604), .Z(n_326889156));
	notech_ao4 i_123042111(.A(n_26716142), .B(n_31524), .C(n_56832), .D(n_32313
		), .Z(n_327089158));
	notech_and4 i_123442107(.A(n_327089158), .B(n_326889156), .C(n_296488864
		), .D(n_296788867), .Z(n_327289160));
	notech_ao4 i_122742114(.A(n_4434), .B(n_31508), .C(n_31532), .D(n_30606)
		, .Z(n_327389161));
	notech_ao4 i_122542116(.A(n_40216277), .B(n_31489), .C(n_61516490), .D(n_59014
		), .Z(n_327589163));
	notech_and4 i_122942112(.A(n_327589163), .B(n_327389161), .C(n_295888858
		), .D(n_296188861), .Z(n_327789165));
	notech_ao4 i_122142120(.A(n_4433), .B(n_58956), .C(n_40316278), .D(n_32703
		), .Z(n_327989167));
	notech_ao4 i_121942122(.A(n_61116486), .B(n_32147), .C(n_56861), .D(n_32197
		), .Z(n_328189169));
	notech_and4 i_122342118(.A(n_328189169), .B(n_327989167), .C(n_295288852
		), .D(n_295588855), .Z(n_328389171));
	notech_ao4 i_121642125(.A(n_58550), .B(n_61816493), .C(n_56880), .D(n_101142452
		), .Z(n_328489172));
	notech_ao4 i_121442127(.A(n_56929), .B(nbus_11271[8]), .C(n_56904), .D(n_32162
		), .Z(n_328689174));
	notech_and4 i_121842123(.A(n_299488894), .B(n_328689174), .C(n_328489172
		), .D(n_294988849), .Z(n_328889176));
	notech_and2 i_8139995(.A(n_1832), .B(n_332489211), .Z(n_329089178));
	notech_nand2 i_18339896(.A(nbus_135[2]), .B(n_22746), .Z(n_329389181));
	notech_nand3 i_17639903(.A(mul64[2]), .B(n_30648), .C(n_61698), .Z(n_330089188
		));
	notech_nand2 i_16939910(.A(cr0[2]), .B(n_23351), .Z(n_330789195));
	notech_nand2 i_119338915(.A(n_27834), .B(n_58247), .Z(n_332389210));
	notech_ao4 i_119238916(.A(n_22752), .B(n_27834), .C(n_57896), .D(nbus_11291
		[2]), .Z(n_332489211));
	notech_ao4 i_118838920(.A(n_58247), .B(n_329089178), .C(n_22752), .D(n_332389210
		), .Z(n_332589212));
	notech_ao4 i_118738921(.A(n_57998), .B(n_32030), .C(n_58007), .D(nbus_11271
		[2]), .Z(n_332689213));
	notech_ao4 i_118538923(.A(n_57917), .B(nbus_11273[10]), .C(n_22742), .D(n_58802
		), .Z(n_332889215));
	notech_ao4 i_118438924(.A(n_57867), .B(n_33167), .C(n_57907), .D(\nbus_11290[10] 
		), .Z(n_332989216));
	notech_and4 i_119038918(.A(n_332989216), .B(n_332889215), .C(n_332689213
		), .D(n_332589212), .Z(n_333189218));
	notech_ao4 i_118138927(.A(n_57887), .B(n_32492), .C(n_58512), .D(\nbus_11290[2] 
		), .Z(n_333289219));
	notech_ao4 i_118038928(.A(n_57987), .B(n_33688), .C(n_23329), .D(n_32454
		), .Z(n_333389220));
	notech_ao4 i_117838930(.A(n_58492), .B(n_31174), .C(n_58215), .D(n_32424
		), .Z(n_333589222));
	notech_and4 i_118338925(.A(n_333589222), .B(n_333389220), .C(n_333289219
		), .D(n_330789195), .Z(n_333789224));
	notech_ao4 i_117438934(.A(n_23359), .B(n_31221), .C(n_57745), .D(n_32378
		), .Z(n_333989226));
	notech_ao4 i_117338935(.A(n_22979), .B(n_59077), .C(n_23383), .D(n_31202
		), .Z(n_334089227));
	notech_ao4 i_117138937(.A(n_22968), .B(n_32823), .C(n_22967), .D(n_32806
		), .Z(n_334389229));
	notech_and4 i_117638932(.A(n_334389229), .B(n_334089227), .C(n_333989226
		), .D(n_330089188), .Z(n_334589231));
	notech_ao4 i_116738940(.A(n_22977), .B(n_32771), .C(n_22976), .D(n_32346
		), .Z(n_334689232));
	notech_ao4 i_116638941(.A(n_22984), .B(n_32738), .C(n_22980), .D(n_32755
		), .Z(n_334789233));
	notech_ao4 i_116438943(.A(n_22745), .B(n_32840), .C(n_22985), .D(n_33687
		), .Z(n_334989235));
	notech_and4 i_117038938(.A(n_334989235), .B(n_334789233), .C(n_334689232
		), .D(n_329389181), .Z(n_335189237));
	notech_ao3 i_56337539(.A(n_339289277), .B(n_338861016), .C(n_30367), .Z(n_335489239
		));
	notech_and2 i_15737343(.A(n_30867), .B(n_349471379), .Z(n_335589240));
	notech_and4 i_15837342(.A(n_58848), .B(n_346789349), .C(n_2090), .D(n_335489239
		), .Z(n_335689241));
	notech_and4 i_15537345(.A(n_57194), .B(n_22474), .C(n_348271368), .D(n_3455
		), .Z(n_335789242));
	notech_and2 i_15637344(.A(n_1830), .B(n_30681), .Z(n_335889243));
	notech_and4 i_15437346(.A(n_48030), .B(n_315271128), .C(n_338089265), .D
		(n_348171367), .Z(n_335989244));
	notech_ao3 i_15237348(.A(n_23747), .B(n_387864409), .C(n_390664437), .Z(n_336089245
		));
	notech_and3 i_15337347(.A(n_390564436), .B(n_23750), .C(n_387964410), .Z
		(n_336189246));
	notech_and4 i_9137407(.A(n_340989293), .B(n_340789291), .C(n_340589290),
		 .D(n_339989284), .Z(n_336289247));
	notech_ao4 i_9237406(.A(n_79512551), .B(n_447368057), .C(n_80312559), .D
		(n_56002), .Z(n_336389248));
	notech_or4 i_46423(.A(n_30304), .B(n_316160789), .C(n_2091), .D(n_33242)
		, .Z(n_336689251));
	notech_and2 i_5873(.A(sema_rw), .B(n_30540), .Z(n_336789252));
	notech_nor2 i_28137261(.A(n_56603), .B(write_ack), .Z(n_336889253));
	notech_or2 i_29437251(.A(n_2032), .B(read_ack), .Z(n_337589260));
	notech_nao3 i_29537250(.A(over_seg[5]), .B(n_61286), .C(n_345189333), .Z
		(n_338089265));
	notech_or2 i_31137239(.A(n_334460972), .B(n_56965), .Z(n_338589270));
	notech_or2 i_30437242(.A(n_391264443), .B(n_33169), .Z(n_338889273));
	notech_or4 i_30137245(.A(instrc[113]), .B(instrc[114]), .C(n_58707), .D(n_327560903
		), .Z(n_339189276));
	notech_or4 i_42137138(.A(n_314960777), .B(n_61065), .C(n_60163), .D(n_30649
		), .Z(n_339289277));
	notech_or4 i_191537603(.A(n_61877), .B(n_4402), .C(n_61711), .D(n_61864)
		, .Z(n_339389278));
	notech_or4 i_36960(.A(n_32484), .B(n_30343), .C(n_61675), .D(n_33242), .Z
		(n_339489279));
	notech_or4 i_69136902(.A(n_30737), .B(all_cnt[3]), .C(n_31369), .D(n_2815
		), .Z(n_339989284));
	notech_nand3 i_150437651(.A(n_30650), .B(n_62441), .C(n_32353), .Z(n_340489289
		));
	notech_ao4 i_138936291(.A(n_76412520), .B(n_30744), .C(n_336389248), .D(n_80512561
		), .Z(n_340589290));
	notech_ao4 i_138836292(.A(n_30739), .B(n_77012526), .C(n_75912515), .D(n_57436
		), .Z(n_340789291));
	notech_ao4 i_138436294(.A(n_30738), .B(n_77712533), .C(n_447268056), .D(n_30617
		), .Z(n_340989293));
	notech_ao4 i_138336295(.A(n_348489366), .B(n_30681), .C(n_336289247), .D
		(n_340489289), .Z(n_341189295));
	notech_ao4 i_81436811(.A(n_58956), .B(n_336189246), .C(n_58238), .D(n_336089245
		), .Z(n_341489298));
	notech_ao4 i_81236813(.A(n_327760905), .B(n_23511), .C(n_23510), .D(n_327660904
		), .Z(n_341689300));
	notech_and4 i_81636809(.A(n_341689300), .B(n_339189276), .C(n_341489298)
		, .D(n_338889273), .Z(n_341889302));
	notech_ao4 i_80636816(.A(n_58664), .B(nbus_11271[0]), .C(n_391164442), .D
		(n_101142452), .Z(n_341989303));
	notech_ao4 i_80336818(.A(n_56035), .B(n_32529), .C(n_26028), .D(n_61607)
		, .Z(n_342189305));
	notech_and4 i_80936814(.A(n_327860906), .B(n_342189305), .C(n_341989303)
		, .D(n_338589270), .Z(n_342489307));
	notech_or2 i_80236819(.A(n_71912476), .B(n_2081), .Z(n_342589308));
	notech_ao4 i_79436823(.A(n_61838), .B(n_335989244), .C(n_324671211), .D(n_342589308
		), .Z(n_342789310));
	notech_ao4 i_79736821(.A(n_2091), .B(n_30618), .C(n_2033), .D(n_61838), 
		.Z(n_342889311));
	notech_and4 i_79536822(.A(n_342889311), .B(n_342789310), .C(n_337589260)
		, .D(n_56583), .Z(n_343189314));
	notech_ao4 i_78436830(.A(n_2091), .B(n_335889243), .C(n_61838), .D(n_335789242
		), .Z(n_343489317));
	notech_ao4 i_78836827(.A(n_61838), .B(n_345589337), .C(n_4470), .D(n_2081
		), .Z(n_343589318));
	notech_nand3 i_80137512(.A(n_4471), .B(n_343589318), .C(n_339389278), .Z
		(n_343789320));
	notech_and4 i_78236832(.A(n_342889311), .B(n_331471271), .C(n_53429), .D
		(n_56583), .Z(n_344289324));
	notech_ao4 i_77736837(.A(n_61838), .B(n_335689241), .C(n_2091), .D(n_335589240
		), .Z(n_344589327));
	notech_or4 i_77536839(.A(n_336789252), .B(n_30720), .C(n_331771274), .D(n_30629
		), .Z(n_345089332));
	notech_and2 i_166494639(.A(n_348071366), .B(n_3469), .Z(n_345189333));
	notech_nand2 i_11294640(.A(over_seg[5]), .B(n_61281), .Z(n_83245324));
	notech_or4 i_55794641(.A(n_49651676), .B(n_63818), .C(n_61824), .D(n_60152
		), .Z(n_345289334));
	notech_or4 i_55594642(.A(n_49651676), .B(n_349271377), .C(n_61924), .D(n_61959
		), .Z(n_345389335));
	notech_or4 i_55694643(.A(n_49651676), .B(n_60182), .C(n_32646), .D(n_63800
		), .Z(n_345489336));
	notech_and3 i_76194644(.A(n_345489336), .B(n_345389335), .C(n_345289334)
		, .Z(n_345589337));
	notech_and3 i_113394645(.A(n_349471379), .B(n_30681), .C(n_347271361), .Z
		(n_345689338));
	notech_and4 i_113594646(.A(n_348271368), .B(n_345589337), .C(n_346789349
		), .D(n_22474), .Z(n_345789339));
	notech_nand2 i_113994647(.A(n_345989341), .B(n_61085), .Z(n_345889340)
		);
	notech_nand2 i_113694648(.A(n_22481), .B(n_58619), .Z(n_345989341));
	notech_nao3 i_114094651(.A(read_ack), .B(n_26086), .C(n_19603), .Z(n_346289344
		));
	notech_or4 i_113894652(.A(n_61877), .B(n_345789339), .C(n_61711), .D(n_61864
		), .Z(n_346389345));
	notech_and4 i_426941(.A(n_346289344), .B(n_347189353), .C(n_346389345), 
		.D(n_345889340), .Z(n_13955));
	notech_and2 i_9594655(.A(n_22467), .B(n_347071359), .Z(n_346789349));
	notech_or4 i_114394658(.A(opd[2]), .B(opd[3]), .C(n_4343), .D(n_579), .Z
		(n_347089352));
	notech_ao4 i_114494659(.A(n_348571371), .B(n_347089352), .C(n_345689338)
		, .D(n_4340), .Z(n_347189353));
	notech_ao3 i_51360187(.A(n_63790), .B(opc[10]), .C(n_333778343), .Z(n_262863569
		));
	notech_or2 i_19371979(.A(n_119987126), .B(n_57020), .Z(n_347589357));
	notech_or2 i_181671978(.A(n_120087127), .B(n_57020), .Z(n_347689358));
	notech_or2 i_13371976(.A(n_120287129), .B(n_57020), .Z(n_347789359));
	notech_or2 i_19471975(.A(n_120387130), .B(n_57020), .Z(n_347889360));
	notech_or2 i_19871974(.A(n_120487131), .B(n_57020), .Z(n_347989361));
	notech_or2 i_20471973(.A(n_120587132), .B(n_57020), .Z(n_348089362));
	notech_or2 i_15771972(.A(n_120687133), .B(n_57024), .Z(n_348189363));
	notech_or2 i_10312(.A(n_118487111), .B(n_348689368), .Z(n_348289364));
	notech_or4 i_26416(.A(n_61864), .B(n_61607), .C(n_33496), .D(n_315892477
		), .Z(n_348389365));
	notech_nand3 i_32767(.A(n_30650), .B(n_62441), .C(read_ack), .Z(n_348489366
		));
	notech_or4 i_1271952(.A(n_61877), .B(n_61711), .C(n_61864), .D(n_33496),
		 .Z(n_348689368));
	notech_ao3 i_3771927(.A(n_390164432), .B(n_128687213), .C(n_137787304), 
		.Z(n_348789369));
	notech_or4 i_4771917(.A(n_32484), .B(n_30343), .C(n_61651), .D(n_33496),
		 .Z(n_348889370));
	notech_or4 i_206137751(.A(n_2039), .B(n_72112478), .C(n_2081), .D(n_30714
		), .Z(n_56583));
	notech_ao3 i_51460186(.A(opa[10]), .B(n_30351), .C(n_60182), .Z(n_262563566
		));
	notech_or4 i_39460274(.A(n_63706), .B(n_440667990), .C(n_63778), .D(nbus_11273
		[13]), .Z(n_262063562));
	notech_nao3 i_40060271(.A(n_63790), .B(opc[13]), .C(n_441868002), .Z(n_261763559
		));
	notech_and4 i_51493(.A(n_151187438), .B(n_151787444), .C(n_150087427), .D
		(n_152287449), .Z(\nbus_11326[0] ));
	notech_nand2 i_21967(.A(instrc[125]), .B(instrc[126]), .Z(n_37407));
	notech_or4 i_49293(.A(n_159487521), .B(n_160887535), .C(n_161587542), .D
		(n_30556), .Z(\nbus_11305[0] ));
	notech_nand2 i_520739(.A(n_162687553), .B(n_162187548), .Z(n_19592));
	notech_nand2 i_520835(.A(n_163787564), .B(n_163287559), .Z(n_19244));
	notech_nand2 i_520963(.A(n_164887575), .B(n_164387570), .Z(n_18896));
	notech_nand2 i_1517581(.A(n_165987586), .B(n_165587582), .Z(n_11650));
	notech_nand2 i_1417580(.A(n_167087597), .B(n_166587592), .Z(n_11644));
	notech_or4 i_189858145(.A(n_32396), .B(n_59120), .C(n_32397), .D(n_61607
		), .Z(n_213333664));
	notech_nand2 i_3218974(.A(n_209988011), .B(n_208988002), .Z(n_20814));
	notech_nand2 i_3118973(.A(n_210988021), .B(n_210488016), .Z(n_20808));
	notech_nand2 i_3018972(.A(n_211988031), .B(n_211488026), .Z(n_20802));
	notech_nand2 i_2918971(.A(n_212988041), .B(n_212488036), .Z(n_20796));
	notech_nand2 i_2818970(.A(n_214088051), .B(n_213588046), .Z(n_20790));
	notech_nand2 i_2718969(.A(n_215088061), .B(n_214588056), .Z(n_20784));
	notech_nand2 i_2618968(.A(n_216088071), .B(n_215588066), .Z(n_20778));
	notech_nand2 i_2518967(.A(n_217088081), .B(n_216588076), .Z(n_20772));
	notech_nand2 i_2418966(.A(n_218188091), .B(n_217588086), .Z(n_20766));
	notech_nand2 i_2318965(.A(n_219188101), .B(n_218688096), .Z(n_20760));
	notech_nand2 i_2218964(.A(n_220188111), .B(n_219688106), .Z(n_20754));
	notech_nand2 i_2118963(.A(n_221188121), .B(n_220688116), .Z(n_20748));
	notech_nand2 i_2018962(.A(n_222188131), .B(n_221688126), .Z(n_20742));
	notech_nand2 i_1918961(.A(n_223188141), .B(n_222688136), .Z(n_20736));
	notech_nand2 i_1818960(.A(n_224188151), .B(n_223688146), .Z(n_20730));
	notech_nand2 i_1718959(.A(n_225188161), .B(n_224688156), .Z(n_20724));
	notech_nand2 i_1618958(.A(n_226188171), .B(n_225688166), .Z(n_20718));
	notech_nand2 i_1518957(.A(n_227188181), .B(n_226688176), .Z(n_20712));
	notech_nand2 i_1418956(.A(n_228188191), .B(n_227688186), .Z(n_20706));
	notech_nand2 i_1318955(.A(n_229188201), .B(n_228688196), .Z(n_20700));
	notech_nand2 i_1218954(.A(n_230188211), .B(n_229688206), .Z(n_20694));
	notech_nand2 i_1118953(.A(n_231188221), .B(n_230688216), .Z(n_20688));
	notech_nand2 i_1018952(.A(n_232288232), .B(n_231788227), .Z(n_20682));
	notech_nand2 i_918951(.A(n_233388243), .B(n_232888238), .Z(n_20676));
	notech_nand2 i_818950(.A(n_234488254), .B(n_233988249), .Z(n_20670));
	notech_nand2 i_718949(.A(n_235588265), .B(n_235088260), .Z(n_20664));
	notech_nand2 i_618948(.A(n_236688276), .B(n_236188271), .Z(n_20658));
	notech_nand2 i_518947(.A(n_237788287), .B(n_237288282), .Z(n_20652));
	notech_nand2 i_418946(.A(n_238888298), .B(n_238388293), .Z(n_20646));
	notech_nand2 i_318945(.A(n_239988309), .B(n_239488304), .Z(n_20640));
	notech_or4 i_118943(.A(n_168987616), .B(n_240388313), .C(n_30567), .D(n_241188321
		), .Z(n_20628));
	notech_mux2 i_55658136(.S(n_61651), .A(n_209188003), .B(n_32368), .Z(n_212433655
		));
	notech_and2 i_55758135(.A(n_4459), .B(n_167887605), .Z(n_212333654));
	notech_ao4 i_67058130(.A(n_30636), .B(n_61651), .C(n_207787991), .D(n_56226
		), .Z(n_211833649));
	notech_or4 i_141558120(.A(instrc[110]), .B(instrc[111]), .C(n_32155), .D
		(n_32156), .Z(n_210833639));
	notech_nand2 i_153358118(.A(n_335489239), .B(n_167187598), .Z(n_210633637
		));
	notech_nand2 i_40160270(.A(opd[13]), .B(n_30354), .Z(n_261463556));
	notech_or4 i_62194664(.A(n_61711), .B(n_61877), .C(n_83245324), .D(n_345189333
		), .Z(n_348989371));
	notech_or4 i_2820986(.A(n_217484594), .B(n_245188354), .C(n_246388365), 
		.D(n_30570), .Z(n_19034));
	notech_or4 i_2720985(.A(n_30574), .B(n_244288346), .C(n_247188372), .D(n_30571
		), .Z(n_19028));
	notech_nand3 i_2821018(.A(n_248088381), .B(n_247988380), .C(n_247888379)
		, .Z(n_18686));
	notech_or4 i_2821178(.A(n_217484594), .B(n_242088330), .C(n_248588386), 
		.D(n_30572), .Z(n_13502));
	notech_or4 i_2721177(.A(n_30574), .B(n_241288322), .C(n_249288393), .D(n_30573
		), .Z(n_13496));
	notech_nand2 i_420738(.A(n_263088531), .B(n_262588526), .Z(n_19586));
	notech_nand2 i_420834(.A(n_264188542), .B(n_263688537), .Z(n_19238));
	notech_or4 i_2020978(.A(n_258888489), .B(n_261285029), .C(n_264588546), 
		.D(n_30581), .Z(n_18986));
	notech_or4 i_1920977(.A(n_262385040), .B(n_258088481), .C(n_265288553), 
		.D(n_30582), .Z(n_18980));
	notech_or4 i_1820976(.A(n_263485051), .B(n_257288473), .C(n_265988560), 
		.D(n_30584), .Z(n_18974));
	notech_or4 i_1720975(.A(n_264585062), .B(n_256488465), .C(n_266688567), 
		.D(n_30585), .Z(n_18968));
	notech_nand2 i_420962(.A(n_268088581), .B(n_267588576), .Z(n_18890));
	notech_nand3 i_2021010(.A(n_268688587), .B(n_268588586), .C(n_268488585)
		, .Z(n_18638));
	notech_nand3 i_1921009(.A(n_269388594), .B(n_269288593), .C(n_269188592)
		, .Z(n_18632));
	notech_nand3 i_1821008(.A(n_270088601), .B(n_269988600), .C(n_269888599)
		, .Z(n_18626));
	notech_nand3 i_1721007(.A(n_270788608), .B(n_270688607), .C(n_270588606)
		, .Z(n_18620));
	notech_or4 i_1921169(.A(n_262385040), .B(n_251288413), .C(n_271288613), 
		.D(n_30587), .Z(n_13448));
	notech_or4 i_1821168(.A(n_263485051), .B(n_250488405), .C(n_271988620), 
		.D(n_30588), .Z(n_13442));
	notech_or4 i_1721167(.A(n_264585062), .B(n_249688397), .C(n_272688627), 
		.D(n_30589), .Z(n_13436));
	notech_or4 i_35860307(.A(n_63716), .B(n_440667990), .C(n_63794), .D(nbus_11273
		[10]), .Z(n_2609));
	notech_or4 i_3220990(.A(n_293885352), .B(n_283388733), .C(n_284488744), 
		.D(n_30602), .Z(n_19058));
	notech_nand2 i_920967(.A(n_285688756), .B(n_285288752), .Z(n_18920));
	notech_nand3 i_3221022(.A(n_286288762), .B(n_286188761), .C(n_286088760)
		, .Z(n_18710));
	notech_nand2 i_920999(.A(n_287288772), .B(n_286888768), .Z(n_18572));
	notech_nand2 i_921063(.A(n_288288782), .B(n_287788777), .Z(n_16271));
	notech_or4 i_3221182(.A(n_293885352), .B(n_278688686), .C(n_288688786), 
		.D(n_30603), .Z(n_13526));
	notech_nand2 i_921159(.A(n_289888798), .B(n_289488794), .Z(n_13388));
	notech_nand2 i_921351(.A(n_290888808), .B(n_290388803), .Z(n_20432));
	notech_nand2 i_921607(.A(n_291788817), .B(n_291388813), .Z(n_13040));
	notech_nand2 i_921895(.A(n_292788827), .B(n_292288822), .Z(n_12340));
	notech_nand2 i_917575(.A(n_293888838), .B(n_293388833), .Z(n_11614));
	notech_xor2 i_166543357(.A(n_31606), .B(n_320851229), .Z(n_56898));
	notech_and4 i_916199(.A(n_312889020), .B(n_312789019), .C(n_313889030), 
		.D(n_312689018), .Z(n_13665));
	notech_nand3 i_816198(.A(n_315689047), .B(n_314889039), .C(n_315289043),
		 .Z(n_13659));
	notech_nand3 i_716197(.A(n_317689066), .B(n_316789058), .C(n_317289062),
		 .Z(n_13653));
	notech_nand3 i_616196(.A(n_319689085), .B(n_318789077), .C(n_319289081),
		 .Z(n_13647));
	notech_nand3 i_516195(.A(n_321889106), .B(n_320989097), .C(n_321489102),
		 .Z(n_13641));
	notech_and4 i_316193(.A(n_324389131), .B(n_323289120), .C(n_322789115), 
		.D(n_323889126), .Z(n_13629));
	notech_and4 i_216192(.A(n_326689154), .B(n_325589143), .C(n_325089138), 
		.D(n_326189149), .Z(n_13623));
	notech_and4 i_116191(.A(n_328889176), .B(n_328389171), .C(n_327789165), 
		.D(n_327289160), .Z(n_13617));
	notech_nao3 i_36160304(.A(n_63752), .B(opc[10]), .C(n_441868002), .Z(n_260663549
		));
	notech_and2 i_148740131(.A(n_57672), .B(n_30526), .Z(n_57047));
	notech_and4 i_317729(.A(n_335189237), .B(n_334589231), .C(n_333789224), 
		.D(n_333189218), .Z(n_17060));
	notech_nand2 i_50781(.A(n_341189295), .B(n_348289364), .Z(\nbus_11320[0] 
		));
	notech_or4 i_49029(.A(n_56734), .B(n_124545737), .C(n_30312), .D(n_30311
		), .Z(\nbus_11304[0] ));
	notech_nand2 i_117567(.A(n_342489307), .B(n_341889302), .Z(n_11566));
	notech_and4 i_526942(.A(n_3326), .B(n_331471271), .C(n_57016), .D(n_343189314
		), .Z(n_13961));
	notech_or4 i_326940(.A(n_30624), .B(n_343789320), .C(n_30622), .D(n_30625
		), .Z(n_13949));
	notech_or4 i_226939(.A(n_343789320), .B(n_336889253), .C(n_30626), .D(n_345089332
		), .Z(n_13943));
	notech_nand2 i_36260303(.A(n_30354), .B(opd[10]), .Z(n_260363546));
	notech_or2 i_11360528(.A(n_386264393), .B(n_31483), .Z(n_259863541));
	notech_or2 i_11860523(.A(n_58664), .B(nbus_11271[10]), .Z(n_259163535)
		);
	notech_ao4 i_6160579(.A(n_63706), .B(n_61924), .C(n_61052), .D(n_58601),
		 .Z(n_258963533));
	notech_or2 i_6360577(.A(n_57705), .B(n_56820), .Z(n_258763531));
	notech_nand3 i_80659899(.A(n_57714), .B(n_272763658), .C(n_258763531), .Z
		(n_258663530));
	notech_or4 i_80059905(.A(n_61824), .B(n_57535), .C(n_57633), .D(n_32219)
		, .Z(n_258463528));
	notech_and4 i_79159914(.A(n_32310), .B(n_61085), .C(n_32321), .D(n_32204
		), .Z(n_2583));
	notech_and4 i_78659919(.A(n_32310), .B(n_61085), .C(n_32323), .D(n_57211
		), .Z(n_258063525));
	notech_and4 i_78559920(.A(n_32310), .B(n_61085), .C(n_32321), .D(n_57211
		), .Z(n_2579));
	notech_or2 i_77859927(.A(n_384864379), .B(n_30553), .Z(n_257363519));
	notech_or4 i_71259993(.A(n_32269), .B(n_384764378), .C(n_384864379), .D(instrc
		[120]), .Z(n_2570));
	notech_nand2 i_71159994(.A(n_382964360), .B(n_30505), .Z(n_256963516));
	notech_or2 i_137060653(.A(n_57705), .B(instrc[116]), .Z(n_256863515));
	notech_ao4 i_124660658(.A(n_63770), .B(n_61959), .C(n_61052), .D(n_30314
		), .Z(n_256763514));
	notech_ao4 i_124760657(.A(n_63786), .B(n_61959), .C(n_26063), .D(n_61052
		), .Z(n_256563512));
	notech_ao3 i_105260669(.A(n_328160909), .B(n_385064381), .C(n_2579), .Z(n_256463511
		));
	notech_ao4 i_66860671(.A(n_57714), .B(n_31036), .C(n_30212), .D(n_55831)
		, .Z(n_20902));
	notech_nand2 i_66360672(.A(n_56002), .B(n_258663530), .Z(n_20898));
	notech_and3 i_48660681(.A(n_2746), .B(n_2748), .C(n_271663649), .Z(n_30468
		));
	notech_and3 i_48460683(.A(n_2749), .B(n_2751), .C(n_271163644), .Z(n_256363510
		));
	notech_or2 i_47260689(.A(n_57553), .B(n_3299), .Z(n_256263509));
	notech_or2 i_46860691(.A(n_57553), .B(n_366164192), .Z(n_30474));
	notech_or4 i_209460707(.A(n_61797), .B(n_32574), .C(n_63700), .D(n_61924
		), .Z(n_26028));
	notech_and3 i_112362278(.A(n_28238), .B(n_255863505), .C(n_234863345), .Z
		(n_256063507));
	notech_ao4 i_112262279(.A(n_24527), .B(n_33193), .C(n_60449), .D(n_31515
		), .Z(n_255863505));
	notech_ao4 i_112462277(.A(n_24717), .B(n_336060988), .C(n_61085), .D(n_30764
		), .Z(n_255663503));
	notech_ao4 i_112562276(.A(n_381164342), .B(n_31480), .C(n_324060868), .D
		(n_380764338), .Z(n_255563502));
	notech_and4 i_113562266(.A(n_255263499), .B(n_255163498), .C(n_254963496
		), .D(n_254863495), .Z(n_255463501));
	notech_ao4 i_112862273(.A(n_381064341), .B(n_33165), .C(n_380964340), .D
		(n_100242443), .Z(n_255263499));
	notech_ao4 i_112962272(.A(n_324160869), .B(n_24430), .C(n_324560873), .D
		(n_24424), .Z(n_255163498));
	notech_ao4 i_113162270(.A(n_324660874), .B(n_24421), .C(n_324260870), .D
		(n_24431), .Z(n_254963496));
	notech_and2 i_113362268(.A(n_236363360), .B(n_254763494), .Z(n_254863495
		));
	notech_ao4 i_113262269(.A(n_24429), .B(n_324760875), .C(n_324460872), .D
		(n_24425), .Z(n_254763494));
	notech_and4 i_115362248(.A(n_58055), .B(n_254463491), .C(n_254263489), .D
		(n_254163488), .Z(n_254663493));
	notech_ao4 i_114862253(.A(n_336463936), .B(n_24542), .C(n_381764348), .D
		(nbus_11273[10]), .Z(n_254463491));
	notech_ao4 i_115062251(.A(n_381664347), .B(n_59023), .C(n_381564346), .D
		(n_336163933), .Z(n_254263489));
	notech_ao4 i_115162250(.A(n_336363935), .B(n_24541), .C(n_336263934), .D
		(n_24539), .Z(n_254163488));
	notech_and4 i_116062241(.A(n_253863485), .B(n_253763484), .C(n_253563482
		), .D(n_253463481), .Z(n_254063487));
	notech_ao4 i_115462247(.A(n_381464345), .B(n_33204), .C(n_381364344), .D
		(n_353164063), .Z(n_253863485));
	notech_ao4 i_115562246(.A(n_3299), .B(n_24716), .C(n_24528), .D(n_33192)
		, .Z(n_253763484));
	notech_ao4 i_115762244(.A(n_24527), .B(n_33191), .C(n_381264343), .D(n_31483
		), .Z(n_253563482));
	notech_ao4 i_115862243(.A(n_60449), .B(n_31518), .C(n_61085), .D(n_30767
		), .Z(n_253463481));
	notech_and4 i_119162210(.A(n_58055), .B(n_253163478), .C(n_252963476), .D
		(n_252863475), .Z(n_253363480));
	notech_ao4 i_118662215(.A(n_366164192), .B(n_24716), .C(n_24528), .D(n_33190
		), .Z(n_253163478));
	notech_ao4 i_118862213(.A(n_24527), .B(n_33189), .C(n_60449), .D(n_31521
		), .Z(n_252963476));
	notech_ao4 i_118962212(.A(n_31498), .B(n_24542), .C(n_31497), .D(n_24541
		), .Z(n_252863475));
	notech_and4 i_119862203(.A(n_252563472), .B(n_252463471), .C(n_252263469
		), .D(n_252163468), .Z(n_252763474));
	notech_ao4 i_119262209(.A(n_31495), .B(n_24539), .C(n_381464345), .D(n_33213
		), .Z(n_252563472));
	notech_ao4 i_119362208(.A(n_381364344), .B(n_375064281), .C(n_381764348)
		, .D(nbus_11273[13]), .Z(n_252463471));
	notech_ao4 i_119562206(.A(n_381664347), .B(\nbus_11290[13] ), .C(n_381564346
		), .D(n_31475), .Z(n_252263469));
	notech_ao4 i_119662205(.A(n_381264343), .B(n_31486), .C(n_61085), .D(n_30770
		), .Z(n_252163468));
	notech_ao3 i_129962112(.A(n_55802), .B(n_30468), .C(n_239263389), .Z(n_251963466
		));
	notech_ao4 i_130062111(.A(n_31495), .B(n_333978345), .C(n_323978248), .D
		(n_33213), .Z(n_251663463));
	notech_and4 i_130762104(.A(n_251363460), .B(n_251163458), .C(n_239863395
		), .D(n_240163398), .Z(n_251563462));
	notech_ao4 i_130362108(.A(n_57243), .B(nbus_11273[13]), .C(\nbus_11290[13] 
		), .D(n_57244), .Z(n_251363460));
	notech_ao4 i_130562106(.A(n_57068), .B(n_30474), .C(n_58030), .D(n_31486
		), .Z(n_251163458));
	notech_and4 i_134962062(.A(n_30274), .B(n_250863456), .C(n_250663454), .D
		(n_240663403), .Z(n_251063457));
	notech_ao4 i_134562066(.A(n_185962886), .B(n_30891), .C(n_3117), .D(n_30916
		), .Z(n_250863456));
	notech_ao4 i_134762064(.A(n_3116), .B(n_30896), .C(n_3111), .D(n_30914),
		 .Z(n_250663454));
	notech_and4 i_135462057(.A(n_250363451), .B(n_241363409), .C(n_250163449
		), .D(n_240963406), .Z(n_250563453));
	notech_ao4 i_135062061(.A(n_26942), .B(n_334360971), .C(n_58229), .D(n_303544469
		), .Z(n_250363451));
	notech_ao4 i_135262059(.A(n_57081), .B(n_30280), .C(n_26951), .D(n_232763324
		), .Z(n_250163449));
	notech_and4 i_135962052(.A(n_249863446), .B(n_249663444), .C(n_30339), .D
		(n_241963414), .Z(n_250063448));
	notech_ao4 i_135562056(.A(n_3112), .B(n_31126), .C(n_3117), .D(n_31119),
		 .Z(n_249863446));
	notech_ao4 i_135762054(.A(n_31123), .B(n_3114), .C(n_3115), .D(n_31125),
		 .Z(n_249663444));
	notech_and4 i_136562046(.A(n_249363441), .B(n_249163439), .C(n_249063438
		), .D(n_2422), .Z(n_249563443));
	notech_ao4 i_136062051(.A(n_3116), .B(n_31099), .C(n_185962886), .D(n_31098
		), .Z(n_249363441));
	notech_ao4 i_136262049(.A(n_305544489), .B(n_31478), .C(n_3118), .D(n_33135
		), .Z(n_249163439));
	notech_ao4 i_136362048(.A(n_26942), .B(n_334860976), .C(n_57081), .D(n_30338
		), .Z(n_249063438));
	notech_ao4 i_136762044(.A(n_387564406), .B(n_60611), .C(n_305644490), .D
		(n_31506), .Z(n_248763435));
	notech_nand3 i_137262039(.A(n_248363431), .B(n_248563433), .C(n_2435), .Z
		(n_248663434));
	notech_ao4 i_136962042(.A(n_387664407), .B(n_5750), .C(n_58483), .D(n_302744461
		), .Z(n_248563433));
	notech_ao4 i_137062041(.A(n_125326580), .B(n_33194), .C(n_125426581), .D
		(n_5758), .Z(n_248363431));
	notech_and4 i_145661957(.A(n_30274), .B(n_248063428), .C(n_247863426), .D
		(n_2440), .Z(n_248263430));
	notech_ao4 i_145161961(.A(n_177362801), .B(n_30891), .C(n_3129), .D(n_30916
		), .Z(n_248063428));
	notech_ao4 i_145361959(.A(n_30896), .B(n_30707), .C(n_3119), .D(n_30914)
		, .Z(n_247863426));
	notech_and4 i_146161952(.A(n_2475), .B(n_244663418), .C(n_2473), .D(n_2443
		), .Z(n_247763425));
	notech_ao4 i_145761956(.A(n_3293), .B(n_334360971), .C(n_58229), .D(n_233663333
		), .Z(n_2475));
	notech_ao4 i_145961954(.A(n_57187), .B(n_30280), .C(n_3290), .D(n_233463331
		), .Z(n_2473));
	notech_and4 i_146661947(.A(n_30339), .B(n_2470), .C(n_2468), .D(n_245163423
		), .Z(n_2472));
	notech_ao4 i_146261951(.A(n_3122), .B(n_31126), .C(n_3129), .D(n_31119),
		 .Z(n_2470));
	notech_ao4 i_146461949(.A(n_31123), .B(n_3124), .C(n_3126), .D(n_31125),
		 .Z(n_2468));
	notech_and4 i_147261941(.A(n_2465), .B(n_2462), .C(n_2461), .D(n_2454), 
		.Z(n_2467));
	notech_ao4 i_146761946(.A(n_31099), .B(n_30707), .C(n_177362801), .D(n_31098
		), .Z(n_2465));
	notech_ao4 i_146961944(.A(n_178762815), .B(n_56983), .C(n_3295), .D(n_33135
		), .Z(n_2462));
	notech_ao4 i_147061943(.A(n_3293), .B(n_334860976), .C(n_57187), .D(n_30338
		), .Z(n_2461));
	notech_ao4 i_172861687(.A(n_32259), .B(n_232463321), .C(n_60182), .D(n_29891
		), .Z(n_2460));
	notech_or2 i_13163228(.A(n_378364314), .B(n_29557), .Z(n_29342));
	notech_ao4 i_31160(.A(n_28240), .B(nbus_11273[7]), .C(n_331360941), .D(\nbus_11290[7] 
		), .Z(n_28238));
	notech_or2 i_6663291(.A(n_380764338), .B(n_32241), .Z(n_24431));
	notech_nao3 i_6963288(.A(n_24736), .B(n_58570), .C(n_380764338), .Z(n_24429
		));
	notech_or4 i_6763290(.A(n_58583), .B(n_24430), .C(instrc[122]), .D(n_61757
		), .Z(n_24428));
	notech_or4 i_7063287(.A(n_58583), .B(n_380764338), .C(instrc[122]), .D(n_61757
		), .Z(n_24425));
	notech_or2 i_5563302(.A(n_380764338), .B(n_24736), .Z(n_24424));
	notech_or2 i_5663301(.A(n_380864339), .B(n_24736), .Z(n_24421));
	notech_or4 i_69862685(.A(n_177362801), .B(n_60163), .C(n_32247), .D(nbus_11273
		[5]), .Z(n_2454));
	notech_nao3 i_70162682(.A(n_63770), .B(opc[5]), .C(n_3119), .Z(n_245163423
		));
	notech_or4 i_67962704(.A(n_3298), .B(n_190662933), .C(n_57476), .D(n_59001
		), .Z(n_244663418));
	notech_or2 i_68262701(.A(n_3295), .B(n_33103), .Z(n_2443));
	notech_or2 i_68562698(.A(n_178762815), .B(n_56956), .Z(n_2440));
	notech_or2 i_62862755(.A(n_302844462), .B(n_58992), .Z(n_2435));
	notech_ao3 i_63362750(.A(opc_10[30]), .B(n_63780), .C(n_387764408), .Z(n_2428
		));
	notech_or2 i_62062763(.A(n_3113), .B(n_31122), .Z(n_2422));
	notech_nao3 i_62362760(.A(n_63790), .B(opc[5]), .C(n_3111), .Z(n_241963414
		));
	notech_or4 i_60162782(.A(n_162262654), .B(n_57401), .C(n_288444319), .D(n_59001
		), .Z(n_241363409));
	notech_or2 i_60462779(.A(n_3118), .B(n_33103), .Z(n_240963406));
	notech_nand2 i_60762776(.A(n_30665), .B(opd[1]), .Z(n_240663403));
	notech_or4 i_54362839(.A(n_63698), .B(n_57393), .C(n_63780), .D(nbus_11273
		[13]), .Z(n_240163398));
	notech_or4 i_54662836(.A(n_58550), .B(n_256563512), .C(n_324078249), .D(n_375064281
		), .Z(n_239863395));
	notech_nao3 i_54962833(.A(n_63790), .B(opc[13]), .C(n_333778343), .Z(n_239563392
		));
	notech_ao3 i_55062832(.A(n_61025), .B(n_30351), .C(n_60182), .Z(n_239263389
		));
	notech_or4 i_34563022(.A(n_61052), .B(n_24430), .C(\nbus_11290[7] ), .D(n_58570
		), .Z(n_236363360));
	notech_nao3 i_35863009(.A(n_3479), .B(n_61275), .C(n_32186), .Z(n_234863345
		));
	notech_or4 i_95062442(.A(n_61823), .B(n_57535), .C(n_30698), .D(n_32224)
		, .Z(n_234763344));
	notech_nand2 i_94362449(.A(n_115942600), .B(n_32224), .Z(n_234363340));
	notech_ao4 i_10663251(.A(n_332363895), .B(n_30919), .C(n_60163), .D(n_58229
		), .Z(n_234063337));
	notech_ao4 i_10763250(.A(n_332363895), .B(n_30920), .C(n_60163), .D(n_59005
		), .Z(n_233863335));
	notech_nao3 i_121169333(.A(n_57480), .B(n_30674), .C(n_190662933), .Z(n_233663333
		));
	notech_nao3 i_121069334(.A(n_32247), .B(n_30674), .C(n_190662933), .Z(n_233563332
		));
	notech_mux2 i_14263217(.S(n_32247), .A(n_234063337), .B(n_233863335), .Z
		(n_233463331));
	notech_ao4 i_10863249(.A(n_26957), .B(n_30919), .C(n_60163), .D(n_58229)
		, .Z(n_233163328));
	notech_ao4 i_10963248(.A(n_26957), .B(n_30920), .C(n_60163), .D(n_59005)
		, .Z(n_232963326));
	notech_mux2 i_14763212(.S(n_32272), .A(n_233163328), .B(n_232963326), .Z
		(n_232763324));
	notech_ao4 i_6063297(.A(n_63740), .B(n_61959), .C(n_29891), .D(n_61052),
		 .Z(n_232463321));
	notech_or2 i_128063348(.A(n_380764338), .B(n_30314), .Z(n_24430));
	notech_and4 i_117465005(.A(n_232063318), .B(n_231863316), .C(n_231763315
		), .D(n_209963112), .Z(n_232363320));
	notech_ao4 i_116965010(.A(n_55975), .B(n_32069), .C(n_55966), .D(n_33188
		), .Z(n_232063318));
	notech_ao4 i_117165008(.A(n_331560943), .B(n_3299), .C(n_55946), .D(n_31518
		), .Z(n_231863316));
	notech_ao4 i_117265007(.A(n_26397), .B(n_336463936), .C(n_26394), .D(n_336363935
		), .Z(n_231763315));
	notech_and4 i_118164998(.A(n_231463313), .B(n_231363312), .C(n_231163310
		), .D(n_231063309), .Z(n_231663314));
	notech_ao4 i_117565004(.A(n_26396), .B(n_336263934), .C(n_378964320), .D
		(n_33204), .Z(n_231463313));
	notech_ao4 i_117665003(.A(n_378864319), .B(n_353164063), .C(n_58303), .D
		(n_378764318), .Z(n_231363312));
	notech_ao4 i_117865001(.A(n_378664317), .B(n_59023), .C(n_378564316), .D
		(n_336163933), .Z(n_231163310));
	notech_ao4 i_117965000(.A(n_378464315), .B(n_31483), .C(n_61087), .D(n_30789
		), .Z(n_231063309));
	notech_and4 i_136664824(.A(n_230763306), .B(n_230563304), .C(n_230463303
		), .D(n_211663127), .Z(n_230963308));
	notech_ao4 i_136164829(.A(n_57006), .B(n_31518), .C(n_336463936), .D(n_334278348
		), .Z(n_230763306));
	notech_ao4 i_136364827(.A(n_336363935), .B(n_334078346), .C(n_336263934)
		, .D(n_334178347), .Z(n_230563304));
	notech_ao4 i_136464826(.A(n_57274), .B(n_33204), .C(n_353164063), .D(n_57275
		), .Z(n_230463303));
	notech_and4 i_137264818(.A(n_230163300), .B(n_229963298), .C(n_229863297
		), .D(n_212363134), .Z(n_230363302));
	notech_ao4 i_136764823(.A(n_59023), .B(n_30320), .C(n_336163933), .D(n_57394
		), .Z(n_230163300));
	notech_ao4 i_136964821(.A(n_58025), .B(n_31483), .C(n_61085), .D(n_30816
		), .Z(n_229963298));
	notech_ao4 i_137064820(.A(n_55913), .B(n_33187), .C(n_55793), .D(n_33186
		), .Z(n_229863297));
	notech_and4 i_140264788(.A(n_229563294), .B(n_229363292), .C(n_229263291
		), .D(n_213063141), .Z(n_229763296));
	notech_ao4 i_139764793(.A(n_57006), .B(n_31521), .C(n_31498), .D(n_334278348
		), .Z(n_229563294));
	notech_ao4 i_139964791(.A(n_31495), .B(n_334178347), .C(n_31497), .D(n_334078346
		), .Z(n_229363292));
	notech_ao4 i_140064790(.A(n_375064281), .B(n_57275), .C(n_57274), .D(n_33213
		), .Z(n_229263291));
	notech_and4 i_140864782(.A(n_228963288), .B(n_228763286), .C(n_228663285
		), .D(n_213763148), .Z(n_229163290));
	notech_ao4 i_140364787(.A(n_57128), .B(nbus_11273[13]), .C(n_31475), .D(n_57394
		), .Z(n_228963288));
	notech_ao4 i_140564785(.A(n_58025), .B(n_31486), .C(n_61087), .D(n_30820
		), .Z(n_228763286));
	notech_ao4 i_140664784(.A(n_55913), .B(n_33185), .C(n_55793), .D(n_33184
		), .Z(n_228663285));
	notech_and4 i_143564755(.A(n_228363282), .B(n_228163280), .C(n_214563155
		), .D(n_214863158), .Z(n_228563284));
	notech_ao4 i_143164759(.A(n_336463936), .B(n_200777063), .C(n_336363935)
		, .D(n_200677062), .Z(n_228363282));
	notech_ao4 i_143364757(.A(n_57252), .B(n_33204), .C(n_353164063), .D(n_57317
		), .Z(n_228163280));
	notech_and4 i_144064750(.A(n_227863277), .B(n_227663275), .C(n_215163161
		), .D(n_215463164), .Z(n_228063279));
	notech_ao4 i_143664754(.A(n_57133), .B(n_59023), .C(n_336163933), .D(n_57388
		), .Z(n_227863277));
	notech_ao4 i_143864752(.A(n_58053), .B(n_31483), .C(n_56896), .D(n_33108
		), .Z(n_227663275));
	notech_ao4 i_145064740(.A(n_56783), .B(n_31521), .C(n_31498), .D(n_200777063
		), .Z(n_227463273));
	notech_ao4 i_145164739(.A(n_31497), .B(n_200677062), .C(n_375064281), .D
		(n_57317), .Z(n_227263271));
	notech_and4 i_145864732(.A(n_226963268), .B(n_226763266), .C(n_217263172
		), .D(n_217563175), .Z(n_227163270));
	notech_ao4 i_145464736(.A(n_57133), .B(n_58965), .C(n_58330), .D(n_57110
		), .Z(n_226963268));
	notech_ao4 i_145664734(.A(n_57152), .B(n_30474), .C(n_58053), .D(n_31486
		), .Z(n_226763266));
	notech_and4 i_158664606(.A(n_226463263), .B(n_226263261), .C(n_226163260
		), .D(n_217863178), .Z(n_226663265));
	notech_ao4 i_158164611(.A(n_333260960), .B(n_33183), .C(n_55884), .D(n_33182
		), .Z(n_226463263));
	notech_ao4 i_158364609(.A(n_336463936), .B(n_28368), .C(n_57006), .D(n_31518
		), .Z(n_226263261));
	notech_ao4 i_158464608(.A(n_336363935), .B(n_28367), .C(n_336263934), .D
		(n_28365), .Z(n_226163260));
	notech_and4 i_159264600(.A(n_225863257), .B(n_225663255), .C(n_225563254
		), .D(n_218563184), .Z(n_226063259));
	notech_ao4 i_158764605(.A(n_353164063), .B(n_444668030), .C(n_58303), .D
		(n_444368027), .Z(n_225863257));
	notech_ao4 i_158964603(.A(n_444468028), .B(n_59023), .C(n_336163933), .D
		(n_444768031), .Z(n_225663255));
	notech_ao4 i_159064602(.A(n_444868032), .B(n_31483), .C(n_61087), .D(n_30845
		), .Z(n_225563254));
	notech_and4 i_162264570(.A(n_225263251), .B(n_225063249), .C(n_224963248
		), .D(n_219263191), .Z(n_225463253));
	notech_ao4 i_161764575(.A(n_333260960), .B(n_33181), .C(n_55884), .D(n_33180
		), .Z(n_225263251));
	notech_ao4 i_161964573(.A(n_31498), .B(n_28368), .C(n_57001), .D(n_31521
		), .Z(n_225063249));
	notech_ao4 i_162064572(.A(n_31495), .B(n_28365), .C(n_31497), .D(n_28367
		), .Z(n_224963248));
	notech_and4 i_162864564(.A(n_224663245), .B(n_224463243), .C(n_224363242
		), .D(n_219863197), .Z(n_224863247));
	notech_ao4 i_162364569(.A(n_444568029), .B(n_33213), .C(n_58965), .D(n_444468028
		), .Z(n_224663245));
	notech_ao4 i_162564567(.A(n_444368027), .B(n_58330), .C(n_31475), .D(n_444768031
		), .Z(n_224463243));
	notech_ao4 i_162664566(.A(n_444868032), .B(n_31486), .C(n_61087), .D(n_30848
		), .Z(n_224363242));
	notech_and4 i_171864474(.A(n_224063239), .B(n_223863237), .C(n_256363510
		), .D(n_220763206), .Z(n_224263241));
	notech_ao4 i_171464478(.A(n_336463936), .B(n_334478350), .C(n_336363935)
		, .D(n_334378349), .Z(n_224063239));
	notech_ao4 i_171664476(.A(n_33204), .B(n_323478243), .C(n_353164063), .D
		(n_323378242), .Z(n_223863237));
	notech_and4 i_172364469(.A(n_223563234), .B(n_223363232), .C(n_221063209
		), .D(n_221363212), .Z(n_223763236));
	notech_ao4 i_171964473(.A(n_57238), .B(n_59023), .C(n_336163933), .D(n_57387
		), .Z(n_223563234));
	notech_ao4 i_172164471(.A(n_58029), .B(n_31483), .C(n_279977810), .D(nbus_11271
		[10]), .Z(n_223363232));
	notech_nand2 i_183864355(.A(n_222963228), .B(n_221763216), .Z(n_223063229
		));
	notech_ao4 i_183764356(.A(n_31497), .B(n_29418), .C(n_375064281), .D(n_57611
		), .Z(n_222963228));
	notech_or4 i_184464349(.A(n_222363222), .B(n_222063219), .C(n_30754), .D
		(n_30755), .Z(n_222863227));
	notech_ao4 i_184064353(.A(n_58965), .B(n_444968033), .C(n_445068034), .D
		(n_58330), .Z(n_222663225));
	notech_ao4 i_184264351(.A(n_57059), .B(n_30474), .C(n_445268036), .D(n_31486
		), .Z(n_222463223));
	notech_nao3 i_2266134(.A(n_30269), .B(n_57467), .C(n_378364314), .Z(n_29341
		));
	notech_or4 i_2766129(.A(n_318060808), .B(n_2577), .C(n_378364314), .D(n_29557
		), .Z(n_29340));
	notech_or2 i_2366133(.A(n_378364314), .B(n_57467), .Z(n_29338));
	notech_or2 i_2666130(.A(n_378364314), .B(n_32244), .Z(n_29337));
	notech_nor2 i_96365205(.A(n_31475), .B(n_445168035), .Z(n_222363222));
	notech_ao3 i_96665202(.A(n_30282), .B(\opa_12[13] ), .C(n_386964400), .Z
		(n_222063219));
	notech_or4 i_96965199(.A(n_61924), .B(n_31624), .C(n_30269), .D(n_29560)
		, .Z(n_221763216));
	notech_ao3 i_97065198(.A(opa[13]), .B(n_29417), .C(n_60182), .Z(n_221463213
		));
	notech_or2 i_83065338(.A(n_57604), .B(n_256263509), .Z(n_221363212));
	notech_or2 i_83365335(.A(n_57237), .B(n_58303), .Z(n_221063209));
	notech_or4 i_83665332(.A(n_61924), .B(n_31621), .C(n_30319), .D(n_323578244
		), .Z(n_220763206));
	notech_or2 i_73365435(.A(n_375064281), .B(n_444668030), .Z(n_219863197)
		);
	notech_or2 i_74065428(.A(n_366164192), .B(n_331760945), .Z(n_219263191)
		);
	notech_or2 i_69165477(.A(n_444568029), .B(n_33204), .Z(n_218563184));
	notech_or2 i_69865470(.A(n_3299), .B(n_331760945), .Z(n_217863178));
	notech_or4 i_53465634(.A(n_63720), .B(n_57388), .C(n_63780), .D(n_58330)
		, .Z(n_217563175));
	notech_or2 i_53765631(.A(n_57252), .B(n_33213), .Z(n_217263172));
	notech_or4 i_54065628(.A(n_192776985), .B(n_61924), .C(n_31624), .D(n_58279
		), .Z(n_216963169));
	notech_or2 i_51065657(.A(n_57152), .B(n_256263509), .Z(n_215463164));
	notech_or2 i_51365654(.A(n_57110), .B(n_58303), .Z(n_215163161));
	notech_or4 i_51765651(.A(n_192776985), .B(n_61928), .C(n_31621), .D(n_58279
		), .Z(n_214863158));
	notech_nand3 i_52065648(.A(n_30524), .B(n_61609), .C(read_data[10]), .Z(n_214563155
		));
	notech_nand2 i_47265693(.A(opb[13]), .B(n_57129), .Z(n_213763148));
	notech_or2 i_47965686(.A(n_366164192), .B(n_328860916), .Z(n_213063141)
		);
	notech_or2 i_42965735(.A(n_57128), .B(n_58303), .Z(n_212363134));
	notech_or2 i_43665728(.A(n_3299), .B(n_328860916), .Z(n_211663127));
	notech_or2 i_22665931(.A(n_55955), .B(n_30987), .Z(n_209963112));
	notech_ao4 i_171067648(.A(n_56407), .B(n_58303), .C(n_61647), .D(n_32602
		), .Z(n_209563109));
	notech_ao4 i_169467663(.A(n_56407), .B(n_58330), .C(n_61651), .D(n_32605
		), .Z(n_209363108));
	notech_ao4 i_145967879(.A(n_59114), .B(n_32952), .C(n_56387), .D(n_32954
		), .Z(n_209163106));
	notech_ao4 i_132068016(.A(n_326560893), .B(n_3115), .C(n_326460892), .D(n_3112
		), .Z(n_208963104));
	notech_and4 i_131968017(.A(n_208063095), .B(n_186862895), .C(n_208563100
		), .D(n_186962896), .Z(n_208863103));
	notech_ao3 i_131568021(.A(n_208363098), .B(n_186562892), .C(n_186462891)
		, .Z(n_208563100));
	notech_and4 i_131368023(.A(n_186362890), .B(n_326860896), .C(n_186162888
		), .D(n_186262889), .Z(n_208363098));
	notech_ao4 i_131668020(.A(n_326660894), .B(n_3113), .C(n_326360891), .D(n_3111
		), .Z(n_208063095));
	notech_ao4 i_129368040(.A(n_325560883), .B(n_3115), .C(n_325460882), .D(n_3112
		), .Z(n_207863093));
	notech_and4 i_129268041(.A(n_206663084), .B(n_185462881), .C(n_207363089
		), .D(n_185562882), .Z(n_207663092));
	notech_ao3 i_128868045(.A(n_206963087), .B(n_185162878), .C(n_184962877)
		, .Z(n_207363089));
	notech_and4 i_128568047(.A(n_184862876), .B(n_325860886), .C(n_184662874
		), .D(n_184762875), .Z(n_206963087));
	notech_ao4 i_128968044(.A(n_325660884), .B(n_3113), .C(n_325360881), .D(n_3111
		), .Z(n_206663084));
	notech_ao4 i_126368064(.A(n_324360871), .B(n_3115), .C(n_324760875), .D(n_3112
		), .Z(n_206463082));
	notech_and4 i_126268065(.A(n_184062868), .B(n_205563073), .C(n_206063078
		), .D(n_184162869), .Z(n_206363081));
	notech_and4 i_125868069(.A(n_183562863), .B(n_183662864), .C(n_183762865
		), .D(n_205763075), .Z(n_206063078));
	notech_and3 i_125568072(.A(n_324860876), .B(n_183362861), .C(n_183462862
		), .Z(n_205763075));
	notech_ao4 i_125968068(.A(n_324260870), .B(n_3113), .C(n_324560873), .D(n_3111
		), .Z(n_205563073));
	notech_ao3 i_121868108(.A(n_182862856), .B(n_182962857), .C(n_205163069)
		, .Z(n_205363071));
	notech_or4 i_121668110(.A(n_182562853), .B(n_182662854), .C(n_182762855)
		, .D(n_204863066), .Z(n_205163069));
	notech_or4 i_121368113(.A(n_182262850), .B(n_30747), .C(n_182362851), .D
		(n_182462852), .Z(n_204863066));
	notech_nao3 i_115368169(.A(n_181762845), .B(n_181662844), .C(n_203863059
		), .Z(n_204163061));
	notech_or4 i_115168171(.A(n_181462842), .B(n_181562843), .C(n_181362841)
		, .D(n_203563056), .Z(n_203863059));
	notech_nand3 i_114868174(.A(n_181162839), .B(n_30468), .C(n_181262840), 
		.Z(n_203563056));
	notech_nao3 i_113368189(.A(n_202963050), .B(n_180662834), .C(n_180562833
		), .Z(n_203163052));
	notech_and4 i_113168191(.A(n_180262830), .B(n_180362831), .C(n_180462832
		), .D(n_377364304), .Z(n_202963050));
	notech_and4 i_109268228(.A(n_327860906), .B(n_179162819), .C(n_202263043
		), .D(n_179462822), .Z(n_202463045));
	notech_ao4 i_109068230(.A(n_3295), .B(n_33169), .C(n_101142452), .D(n_3293
		), .Z(n_202263043));
	notech_ao4 i_109368227(.A(n_58956), .B(n_178962817), .C(n_56965), .D(n_178762815
		), .Z(n_201963040));
	notech_and4 i_107468246(.A(n_200463028), .B(n_201363034), .C(n_178462812
		), .D(n_178162809), .Z(n_201663037));
	notech_ao3 i_106768250(.A(n_201063032), .B(n_177962807), .C(n_178062808)
		, .Z(n_201363034));
	notech_and4 i_106568252(.A(n_200863030), .B(n_177862806), .C(n_177562803
		), .D(n_326860896), .Z(n_201063032));
	notech_ao4 i_106368254(.A(n_3295), .B(n_33167), .C(n_100842449), .D(n_3293
		), .Z(n_200863030));
	notech_ao4 i_107168248(.A(n_326760895), .B(n_3124), .C(n_326360891), .D(n_3119
		), .Z(n_200463028));
	notech_and4 i_104568270(.A(n_199063017), .B(n_199863023), .C(n_177062798
		), .D(n_176762795), .Z(n_200263026));
	notech_ao3 i_104168274(.A(n_199463021), .B(n_176562793), .C(n_176662794)
		, .Z(n_199863023));
	notech_and4 i_103868276(.A(n_199263019), .B(n_176462792), .C(n_325860886
		), .D(n_176162789), .Z(n_199463021));
	notech_ao4 i_103668278(.A(n_3295), .B(n_33166), .C(n_100542446), .D(n_3293
		), .Z(n_199263019));
	notech_ao4 i_104368272(.A(n_325760885), .B(n_3124), .C(n_325360881), .D(n_3119
		), .Z(n_199063017));
	notech_nao3 i_101968295(.A(n_175762785), .B(n_198563012), .C(n_175462782
		), .Z(n_198763014));
	notech_and4 i_101668298(.A(n_175162779), .B(n_175362781), .C(n_198263009
		), .D(n_175262780), .Z(n_198563012));
	notech_and3 i_101368301(.A(n_324860876), .B(n_174862776), .C(n_198163008
		), .Z(n_198263009));
	notech_ao4 i_101268302(.A(n_3295), .B(n_33165), .C(n_100242443), .D(n_3293
		), .Z(n_198163008));
	notech_ao4 i_101868296(.A(n_324460872), .B(n_3124), .C(n_324560873), .D(n_3119
		), .Z(n_197963006));
	notech_ao4 i_92668377(.A(n_31498), .B(n_28742), .C(n_31497), .D(n_28743)
		, .Z(n_197863005));
	notech_or4 i_92368380(.A(n_174162769), .B(n_173962767), .C(n_197262999),
		 .D(n_174062768), .Z(n_197563002));
	notech_nand3 i_92068383(.A(n_197162998), .B(n_173662764), .C(n_30468), .Z
		(n_197262999));
	notech_ao4 i_91968384(.A(n_28855), .B(n_33213), .C(n_375064281), .D(n_28860
		), .Z(n_197162998));
	notech_and4 i_90468398(.A(n_172962759), .B(n_196562992), .C(n_173062760)
		, .D(n_173162761), .Z(n_196862995));
	notech_and3 i_90168401(.A(n_172462756), .B(n_196462991), .C(n_377364304)
		, .Z(n_196562992));
	notech_ao4 i_90068402(.A(n_28855), .B(n_33215), .C(n_97342414), .D(n_28860
		), .Z(n_196462991));
	notech_ao4 i_83968456(.A(n_326760895), .B(n_29678), .C(n_326560893), .D(n_29677
		), .Z(n_196162988));
	notech_and4 i_83768457(.A(n_195662983), .B(n_195462981), .C(n_195362980)
		, .D(n_195862985), .Z(n_196062987));
	notech_and3 i_83468460(.A(n_326860896), .B(n_170862740), .C(n_171562747)
		, .Z(n_195862985));
	notech_ao4 i_83368461(.A(n_326060888), .B(n_57130), .C(n_376964300), .D(n_33167
		), .Z(n_195662983));
	notech_ao4 i_83268462(.A(n_100842449), .B(n_376864299), .C(n_326160889),
		 .D(n_94542386), .Z(n_195462981));
	notech_ao4 i_83168463(.A(n_325960887), .B(n_376564296), .C(n_326360891),
		 .D(n_376764298), .Z(n_195362980));
	notech_ao4 i_84068455(.A(n_326460892), .B(n_29681), .C(n_326660894), .D(n_29680
		), .Z(n_195262979));
	notech_and4 i_74568546(.A(n_194962976), .B(n_194862975), .C(n_170662738)
		, .D(n_194662973), .Z(n_195162978));
	notech_ao4 i_73968552(.A(n_446068044), .B(n_33204), .C(n_445968043), .D(n_353164063
		), .Z(n_194962976));
	notech_ao4 i_73868553(.A(n_4418), .B(n_336363935), .C(n_442182452), .D(n_336263934
		), .Z(n_194862975));
	notech_nor2 i_73768554(.A(n_169762729), .B(n_30747), .Z(n_194662973));
	notech_ao4 i_74168550(.A(n_57136), .B(n_256263509), .C(n_62442065), .D(n_336163933
		), .Z(n_194462971));
	notech_ao4 i_74068551(.A(n_62642067), .B(n_58303), .C(n_62742068), .D(n_59023
		), .Z(n_194362970));
	notech_and4 i_68568606(.A(n_194062967), .B(n_193962966), .C(n_169562727)
		, .D(n_193762964), .Z(n_194262969));
	notech_ao4 i_67968612(.A(n_446068044), .B(n_33213), .C(n_445968043), .D(n_375064281
		), .Z(n_194062967));
	notech_ao4 i_67868613(.A(n_4418), .B(n_31497), .C(n_442182452), .D(n_31495
		), .Z(n_193962966));
	notech_nor2 i_67768614(.A(n_168662718), .B(n_30559), .Z(n_193762964));
	notech_ao4 i_68168610(.A(n_57136), .B(n_30474), .C(n_62442065), .D(n_31475
		), .Z(n_193562962));
	notech_ao4 i_68068611(.A(n_62642067), .B(n_58330), .C(n_62742068), .D(n_58965
		), .Z(n_193462961));
	notech_and4 i_47368815(.A(n_193162958), .B(n_193062957), .C(n_168462716)
		, .D(n_192862955), .Z(n_193362960));
	notech_ao4 i_46768821(.A(n_304744481), .B(n_33213), .C(n_304644480), .D(n_375064281
		), .Z(n_193162958));
	notech_ao4 i_46668822(.A(n_30075), .B(n_31497), .C(n_30078), .D(n_31495)
		, .Z(n_193062957));
	notech_nor2 i_46568823(.A(n_167562707), .B(n_30559), .Z(n_192862955));
	notech_ao4 i_46968819(.A(n_57112), .B(n_30474), .C(n_72542166), .D(n_31475
		), .Z(n_192662953));
	notech_ao4 i_46868820(.A(n_72742168), .B(n_58330), .C(n_4924), .D(n_58965
		), .Z(n_192562952));
	notech_and4 i_29568985(.A(n_192262949), .B(n_192162948), .C(n_191962946)
		, .D(n_167362705), .Z(n_192462951));
	notech_ao4 i_28968991(.A(n_442168005), .B(n_33204), .C(n_442268006), .D(n_353164063
		), .Z(n_192262949));
	notech_ao4 i_28868992(.A(n_445668040), .B(n_336363935), .C(n_445868042),
		 .D(n_336263934), .Z(n_192162948));
	notech_and2 i_28768993(.A(n_166462696), .B(n_256363510), .Z(n_191962946)
		);
	notech_ao4 i_29168989(.A(n_57163), .B(n_256263509), .C(n_91142352), .D(n_336163933
		), .Z(n_191762944));
	notech_ao4 i_29068990(.A(n_91442355), .B(nbus_11273[10]), .C(n_91542356)
		, .D(n_59023), .Z(n_191662943));
	notech_and4 i_22769045(.A(n_191362940), .B(n_191262939), .C(n_191062937)
		, .D(n_166262694), .Z(n_191562942));
	notech_ao4 i_22169051(.A(n_442168005), .B(n_33213), .C(n_442268006), .D(n_375064281
		), .Z(n_191362940));
	notech_ao4 i_22069052(.A(n_445668040), .B(n_31497), .C(n_445868042), .D(n_31495
		), .Z(n_191262939));
	notech_and2 i_21969053(.A(n_165362685), .B(n_30468), .Z(n_191062937));
	notech_ao4 i_22369049(.A(n_57163), .B(n_30474), .C(n_91142352), .D(n_31475
		), .Z(n_190862935));
	notech_ao4 i_22269050(.A(n_91442355), .B(n_58330), .C(n_91542356), .D(n_58965
		), .Z(n_190762934));
	notech_and3 i_105669292(.A(n_57544), .B(n_3292), .C(n_3310), .Z(n_190662933
		));
	notech_and4 i_8169182(.A(n_189762924), .B(n_164062672), .C(n_163962671),
		 .D(n_163862670), .Z(n_190362930));
	notech_and4 i_7969184(.A(n_163762669), .B(n_163662668), .C(n_189462921),
		 .D(n_163562667), .Z(n_189762924));
	notech_ao4 i_7569188(.A(n_58583), .B(n_30257), .C(n_30333), .D(n_30249),
		 .Z(n_189462921));
	notech_nao3 i_6169202(.A(n_63818), .B(instrc[124]), .C(n_163062662), .Z(n_189162918
		));
	notech_ao4 i_144669286(.A(n_57633), .B(n_2810), .C(n_30798), .D(n_32208)
		, .Z(n_188862915));
	notech_ao3 i_4669217(.A(n_57705), .B(n_57686), .C(n_57714), .Z(n_188662913
		));
	notech_nand2 i_1127350(.A(n_209563109), .B(n_188262909), .Z(n_188562912)
		);
	notech_nao3 i_170967649(.A(n_3498), .B(n_60605), .C(n_56428), .Z(n_188262909
		));
	notech_nand2 i_1427353(.A(n_209363108), .B(n_187862905), .Z(n_188162908)
		);
	notech_nao3 i_169267664(.A(n_3501), .B(n_60605), .C(n_56428), .Z(n_187862905
		));
	notech_nand3 i_1427481(.A(n_209163106), .B(n_187662903), .C(n_187362900)
		, .Z(n_187762904));
	notech_or2 i_145767881(.A(n_309892426), .B(n_58965), .Z(n_187662903));
	notech_nao3 i_145867880(.A(n_3565), .B(opb[31]), .C(n_56428), .Z(n_187362900
		));
	notech_nand3 i_321601(.A(n_208963104), .B(n_208863103), .C(n_186062887),
		 .Z(n_187262899));
	notech_or2 i_130168034(.A(n_100842449), .B(n_26942), .Z(n_186962896));
	notech_or4 i_130468032(.A(n_60182), .B(n_26957), .C(n_185962886), .D(n_58247
		), .Z(n_186862895));
	notech_or4 i_130768029(.A(n_60163), .B(n_185962886), .C(n_57401), .D(\nbus_11290[2] 
		), .Z(n_186562892));
	notech_nor2 i_129968035(.A(n_326160889), .B(n_185962886), .Z(n_186462891
		));
	notech_nao3 i_130568031(.A(n_63776), .B(opc_10[2]), .C(n_3117), .Z(n_186362890
		));
	notech_nand2 i_129868036(.A(opd[2]), .B(n_30665), .Z(n_186262889));
	notech_or2 i_129668037(.A(n_326060888), .B(n_57081), .Z(n_186162888));
	notech_or2 i_130268033(.A(n_3118), .B(n_33167), .Z(n_186062887));
	notech_and2 i_106869341(.A(n_288444319), .B(n_26951), .Z(n_185962886));
	notech_nand3 i_721605(.A(n_207863093), .B(n_207663092), .C(n_184562873),
		 .Z(n_185862885));
	notech_or2 i_126968058(.A(n_100542446), .B(n_26942), .Z(n_185562882));
	notech_or4 i_127568056(.A(n_63716), .B(n_3116), .C(n_61924), .D(n_58265)
		, .Z(n_185462881));
	notech_or4 i_127868053(.A(n_60163), .B(n_185962886), .C(n_57401), .D(\nbus_11290[6] 
		), .Z(n_185162878));
	notech_nor2 i_126868059(.A(n_325160879), .B(n_185962886), .Z(n_184962877
		));
	notech_nao3 i_127668055(.A(n_63748), .B(opc_10[6]), .C(n_3117), .Z(n_184862876
		));
	notech_nand2 i_126768060(.A(opd[6]), .B(n_30665), .Z(n_184762875));
	notech_or2 i_126668061(.A(n_325060878), .B(n_57081), .Z(n_184662874));
	notech_or2 i_127468057(.A(n_3118), .B(n_33166), .Z(n_184562873));
	notech_nand3 i_821606(.A(n_206463082), .B(n_206363081), .C(n_183262860),
		 .Z(n_184462872));
	notech_or2 i_124468082(.A(n_100242443), .B(n_26942), .Z(n_184162869));
	notech_or4 i_124668080(.A(n_63716), .B(n_3116), .C(n_61924), .D(nbus_11273
		[7]), .Z(n_184062868));
	notech_or2 i_125068077(.A(n_324460872), .B(n_3114), .Z(n_183762865));
	notech_or4 i_124368083(.A(n_63716), .B(n_185962886), .C(n_63780), .D(n_58275
		), .Z(n_183662864));
	notech_nao3 i_124768079(.A(n_63796), .B(opc_10[7]), .C(n_3117), .Z(n_183562863
		));
	notech_nand2 i_124268084(.A(n_30665), .B(opd[7]), .Z(n_183462862));
	notech_or2 i_124168085(.A(n_323760865), .B(n_57081), .Z(n_183362861));
	notech_or2 i_124568081(.A(n_3118), .B(n_33165), .Z(n_183262860));
	notech_nand3 i_1121609(.A(n_183062858), .B(n_205363071), .C(n_182162849)
		, .Z(n_183162859));
	notech_or2 i_120368119(.A(n_26935), .B(n_33204), .Z(n_183062858));
	notech_nand2 i_120168121(.A(n_30522), .B(opa[10]), .Z(n_182962857));
	notech_or4 i_120268120(.A(n_162262654), .B(n_57401), .C(n_26951), .D(n_353164063
		), .Z(n_182862856));
	notech_and3 i_120468118(.A(n_63796), .B(opc[10]), .C(n_26823), .Z(n_182762855
		));
	notech_ao3 i_120668116(.A(opa[10]), .B(n_26822), .C(n_60182), .Z(n_182662854
		));
	notech_nor2 i_119968123(.A(n_303844472), .B(n_336163933), .Z(n_182562853
		));
	notech_ao3 i_120568117(.A(n_63794), .B(opc_10[10]), .C(n_26821), .Z(n_182462852
		));
	notech_and2 i_119868124(.A(n_305144485), .B(opd[10]), .Z(n_182362851));
	notech_nor2 i_119768125(.A(n_57081), .B(n_256263509), .Z(n_182262850));
	notech_nand2 i_120068122(.A(n_30523), .B(opb[10]), .Z(n_182162849));
	notech_or4 i_1421612(.A(n_181862846), .B(n_204163061), .C(n_181962847), 
		.D(n_181062838), .Z(n_182062848));
	notech_nor2 i_114368179(.A(n_26935), .B(n_33213), .Z(n_181962847));
	notech_and2 i_114168181(.A(n_30522), .B(opa[13]), .Z(n_181862846));
	notech_or4 i_114268180(.A(n_162262654), .B(n_57401), .C(n_26951), .D(n_375064281
		), .Z(n_181762845));
	notech_nand3 i_114468178(.A(n_63796), .B(opc[13]), .C(n_26823), .Z(n_181662844
		));
	notech_ao3 i_114668176(.A(opa[13]), .B(n_26822), .C(n_60182), .Z(n_181562843
		));
	notech_nor2 i_113968183(.A(n_303844472), .B(n_31475), .Z(n_181462842));
	notech_ao3 i_114568177(.A(n_63794), .B(opc_10[13]), .C(n_26821), .Z(n_181362841
		));
	notech_nand2 i_113868184(.A(n_305144485), .B(opd[13]), .Z(n_181262840)
		);
	notech_or2 i_113768185(.A(n_57081), .B(n_30474), .Z(n_181162839));
	notech_and2 i_114068182(.A(n_30523), .B(opb[13]), .Z(n_181062838));
	notech_or4 i_1521613(.A(n_180762835), .B(n_203163052), .C(n_180862836), 
		.D(n_180062828), .Z(n_180962837));
	notech_nor2 i_112468198(.A(n_26935), .B(n_33215), .Z(n_180862836));
	notech_and2 i_112768195(.A(opb[14]), .B(n_179962827), .Z(n_180762835));
	notech_or4 i_112368199(.A(n_162262654), .B(n_57401), .C(n_26951), .D(n_97342414
		), .Z(n_180662834));
	notech_and3 i_112568197(.A(n_63770), .B(opc[14]), .C(n_26823), .Z(n_180562833
		));
	notech_nao3 i_112668196(.A(n_63796), .B(opc_10[14]), .C(n_26821), .Z(n_180462832
		));
	notech_nand2 i_112268200(.A(n_305144485), .B(opd[14]), .Z(n_180362831)
		);
	notech_or2 i_112168201(.A(n_57081), .B(n_377064301), .Z(n_180262830));
	notech_nand3 i_112068202(.A(n_301744451), .B(n_3118), .C(n_302744461), .Z
		(n_180162829));
	notech_and2 i_112868194(.A(opa[14]), .B(n_180162829), .Z(n_180062828));
	notech_nand3 i_111968203(.A(n_301844452), .B(n_26942), .C(n_302844462), 
		.Z(n_179962827));
	notech_and4 i_121151(.A(n_202463045), .B(n_201963040), .C(n_179762825), 
		.D(n_178862816), .Z(n_179862826));
	notech_nand2 i_108868232(.A(opa[0]), .B(n_179062818), .Z(n_179762825));
	notech_nao3 i_108668234(.A(n_63794), .B(opc_10[0]), .C(n_3129), .Z(n_179462822
		));
	notech_or4 i_108168239(.A(instrc[113]), .B(instrc[114]), .C(n_32217), .D
		(n_327560903), .Z(n_179162819));
	notech_nao3 i_108068240(.A(n_28874), .B(n_28855), .C(n_3296), .Z(n_179062818
		));
	notech_and3 i_107968241(.A(n_3294), .B(n_28863), .C(n_28860), .Z(n_178962817
		));
	notech_nao3 i_108568235(.A(n_63796), .B(opc[0]), .C(n_3119), .Z(n_178862816
		));
	notech_and2 i_43169359(.A(n_28854), .B(n_164862680), .Z(n_178762815));
	notech_nao3 i_321153(.A(n_178562813), .B(n_201663037), .C(n_177462802), 
		.Z(n_178662814));
	notech_or4 i_106068257(.A(n_332363895), .B(n_177362801), .C(n_326560893)
		, .D(n_57476), .Z(n_178562813));
	notech_or4 i_105368262(.A(n_60182), .B(n_177362801), .C(n_58247), .D(n_332363895
		), .Z(n_178462812));
	notech_or4 i_105868259(.A(n_60163), .B(n_177362801), .C(n_58247), .D(n_32247
		), .Z(n_178162809));
	notech_nor2 i_105268263(.A(n_326160889), .B(n_177362801), .Z(n_178062808
		));
	notech_or2 i_105168264(.A(n_178762815), .B(n_58802), .Z(n_177962807));
	notech_nao3 i_105468261(.A(n_63792), .B(opc_10[2]), .C(n_3129), .Z(n_177862806
		));
	notech_or4 i_104868267(.A(instrc[113]), .B(n_60431), .C(n_32217), .D(n_326060888
		), .Z(n_177562803));
	notech_ao3 i_106168256(.A(n_57476), .B(n_3127), .C(n_326460892), .Z(n_177462802
		));
	notech_and2 i_106969340(.A(n_3290), .B(n_190662933), .Z(n_177362801));
	notech_nao3 i_721157(.A(n_177162799), .B(n_200263026), .C(n_176062788), 
		.Z(n_177262800));
	notech_or4 i_103368281(.A(n_61052), .B(\nbus_11290[6] ), .C(n_57476), .D
		(n_30707), .Z(n_177162799));
	notech_or4 i_102868286(.A(n_63706), .B(n_61924), .C(n_58265), .D(n_30707
		), .Z(n_177062798));
	notech_or4 i_103168283(.A(n_60170), .B(n_177362801), .C(n_58265), .D(n_32247
		), .Z(n_176762795));
	notech_nor2 i_102768287(.A(n_325160879), .B(n_177362801), .Z(n_176662794
		));
	notech_or2 i_102668288(.A(n_178762815), .B(n_31479), .Z(n_176562793));
	notech_nao3 i_102968285(.A(n_63740), .B(opc_10[6]), .C(n_3129), .Z(n_176462792
		));
	notech_or4 i_102368291(.A(instrc[113]), .B(n_60431), .C(n_32217), .D(n_325060878
		), .Z(n_176162789));
	notech_ao3 i_103468280(.A(n_57476), .B(n_3127), .C(n_325460882), .Z(n_176062788
		));
	notech_or4 i_821158(.A(n_174762775), .B(n_198763014), .C(n_175862786), .D
		(n_30756), .Z(n_175962787));
	notech_nor2 i_100968305(.A(n_324360871), .B(n_3126), .Z(n_175862786));
	notech_or4 i_100468310(.A(n_63716), .B(n_61924), .C(n_58275), .D(n_30707
		), .Z(n_175762785));
	notech_nor2 i_100768307(.A(n_324260870), .B(n_3123), .Z(n_175462782));
	notech_or4 i_100368311(.A(n_63718), .B(n_177362801), .C(n_63758), .D(n_58275
		), .Z(n_175362781));
	notech_or2 i_100268312(.A(n_178762815), .B(n_31480), .Z(n_175262780));
	notech_nao3 i_100568309(.A(n_63770), .B(opc_10[7]), .C(n_3129), .Z(n_175162779
		));
	notech_or4 i_99968315(.A(n_60440), .B(n_60431), .C(n_32217), .D(n_323760865
		), .Z(n_174862776));
	notech_ao3 i_101068304(.A(n_57476), .B(n_3127), .C(n_324760875), .Z(n_174762775
		));
	notech_or4 i_1421164(.A(n_174262770), .B(n_197563002), .C(n_174362771), 
		.D(n_30757), .Z(n_174662774));
	notech_nor2 i_91368389(.A(n_302944463), .B(n_58330), .Z(n_174362771));
	notech_and2 i_91268390(.A(n_30631), .B(opb[13]), .Z(n_174262770));
	notech_nor2 i_91168391(.A(n_303744471), .B(n_31475), .Z(n_174162769));
	notech_and2 i_91068392(.A(n_305044484), .B(opd[13]), .Z(n_174062768));
	notech_ao3 i_91568387(.A(n_63768), .B(opc_10[13]), .C(n_28741), .Z(n_173962767
		));
	notech_or2 i_90768395(.A(n_57189), .B(n_30474), .Z(n_173662764));
	notech_nao3 i_1521165(.A(n_173262762), .B(n_196862995), .C(n_172162753),
		 .Z(n_173562763));
	notech_nand2 i_89368408(.A(n_305044484), .B(opd[14]), .Z(n_173262762));
	notech_nao3 i_89568406(.A(n_63770), .B(opc_10[14]), .C(n_28741), .Z(n_173162761
		));
	notech_nand2 i_89868404(.A(opb[14]), .B(n_172362755), .Z(n_173062760));
	notech_nand2 i_89768405(.A(opa[14]), .B(n_172262754), .Z(n_172962759));
	notech_or2 i_89068411(.A(n_57189), .B(n_377064301), .Z(n_172462756));
	notech_nand3 i_88968412(.A(n_3294), .B(n_3293), .C(n_28863), .Z(n_172362755
		));
	notech_nao3 i_88868413(.A(n_3295), .B(n_28874), .C(n_3296), .Z(n_172262754
		));
	notech_ao3 i_89468407(.A(n_63790), .B(opc[14]), .C(n_28743), .Z(n_172162753
		));
	notech_nand3 i_320961(.A(n_196162988), .B(n_195262979), .C(n_196062987),
		 .Z(n_172062752));
	notech_or2 i_82568469(.A(n_54741988), .B(n_58802), .Z(n_171562747));
	notech_nao3 i_81768476(.A(n_63768), .B(opc_10[2]), .C(n_376664297), .Z(n_170862740
		));
	notech_nand3 i_1120969(.A(n_194462971), .B(n_194362970), .C(n_195162978)
		, .Z(n_170762739));
	notech_or2 i_73668555(.A(n_62142062), .B(n_31483), .Z(n_170662738));
	notech_ao3 i_72768564(.A(opa[10]), .B(n_442082451), .C(n_60182), .Z(n_169762729
		));
	notech_nand3 i_1420972(.A(n_193562962), .B(n_193462961), .C(n_194262969)
		, .Z(n_169662728));
	notech_or2 i_67668615(.A(n_62142062), .B(n_31486), .Z(n_169562727));
	notech_ao3 i_66768624(.A(opa[13]), .B(n_442082451), .C(n_60182), .Z(n_168662718
		));
	notech_nand3 i_1420844(.A(n_192662953), .B(n_192562952), .C(n_193362960)
		, .Z(n_168562717));
	notech_or2 i_46468824(.A(n_4922), .B(n_31486), .Z(n_168462716));
	notech_ao3 i_45568833(.A(opa[13]), .B(n_30076), .C(n_60188), .Z(n_167562707
		));
	notech_nand3 i_1120745(.A(n_191762944), .B(n_191662943), .C(n_192462951)
		, .Z(n_167462706));
	notech_or2 i_28668994(.A(n_90742348), .B(n_31483), .Z(n_167362705));
	notech_or4 i_27569003(.A(n_91142352), .B(n_55831), .C(n_60189), .D(n_58303
		), .Z(n_166462696));
	notech_nand3 i_1420748(.A(n_190862935), .B(n_190762934), .C(n_191562942)
		, .Z(n_166362695));
	notech_or2 i_21869054(.A(n_90742348), .B(n_31486), .Z(n_166262694));
	notech_or4 i_20969063(.A(n_91142352), .B(n_55831), .C(n_60189), .D(n_58330
		), .Z(n_165362685));
	notech_nao3 i_13869126(.A(n_57476), .B(n_30674), .C(n_3291), .Z(n_165262684
		));
	notech_or4 i_12269142(.A(n_61824), .B(n_57535), .C(n_57662), .D(n_32208)
		, .Z(n_165062682));
	notech_nand2 i_10969154(.A(n_115442595), .B(n_32216), .Z(n_164962681));
	notech_nand2 i_10169162(.A(n_115942600), .B(n_32216), .Z(n_164862680));
	notech_nand2 i_9969164(.A(n_115942600), .B(n_32208), .Z(n_164762679));
	notech_ao4 i_25769367(.A(n_32208), .B(n_30316), .C(n_57562), .D(n_57633)
		, .Z(n_164562677));
	notech_and4 i_49803(.A(n_164262674), .B(n_163162663), .C(n_164162673), .D
		(n_190362930), .Z(n_164362675));
	notech_or4 i_6969194(.A(n_56792), .B(n_162262654), .C(n_163062662), .D(n_58583
		), .Z(n_164262674));
	notech_nand3 i_6869195(.A(instrc[116]), .B(n_188662913), .C(n_162962661)
		, .Z(n_164162673));
	notech_nao3 i_6769196(.A(n_63790), .B(n_26957), .C(n_188862915), .Z(n_164062672
		));
	notech_or4 i_7269191(.A(n_30551), .B(n_322660854), .C(n_30332), .D(n_30550
		), .Z(n_163962671));
	notech_or4 i_7169192(.A(n_30551), .B(n_30234), .C(instrc[107]), .D(n_371764248
		), .Z(n_163862670));
	notech_nao3 i_6669197(.A(n_30869), .B(n_143460302), .C(n_26662), .Z(n_163762669
		));
	notech_nao3 i_6569198(.A(n_30869), .B(n_143360301), .C(n_26663), .Z(n_163662668
		));
	notech_or2 i_6469199(.A(n_57081), .B(n_114845640), .Z(n_163562667));
	notech_or4 i_113273405(.A(n_314960777), .B(n_32627), .C(n_61052), .D(n_61838
		), .Z(n_97090337));
	notech_or4 i_113773400(.A(n_61797), .B(n_2152), .C(n_61775), .D(n_63800)
		, .Z(n_97590342));
	notech_or4 i_113873399(.A(n_61797), .B(n_2152), .C(\opcode[0] ), .D(n_63800
		), .Z(n_97690343));
	notech_or4 i_113973398(.A(n_61838), .B(n_61797), .C(n_32628), .D(n_60152
		), .Z(n_97790344));
	notech_or4 i_114073397(.A(n_61838), .B(n_61797), .C(n_32391), .D(n_60154
		), .Z(n_97890345));
	notech_or4 i_20850(.A(instrc[123]), .B(n_61964), .C(n_32250), .D(n_124890615
		), .Z(n_97990346));
	notech_or4 i_18745(.A(n_58583), .B(n_124890615), .C(instrc[122]), .D(n_61757
		), .Z(n_98090347));
	notech_or4 i_18741(.A(n_32269), .B(n_124890615), .C(n_61757), .D(n_23389
		), .Z(n_98190348));
	notech_or4 i_17354(.A(n_124190608), .B(\opcode[1] ), .C(n_63762), .D(n_61775
		), .Z(n_98290349));
	notech_or4 i_17352(.A(n_124190608), .B(\opcode[1] ), .C(n_63762), .D(\opcode[0] 
		), .Z(n_98390350));
	notech_or4 i_17351(.A(n_124190608), .B(n_63762), .C(n_61953), .D(\opcode[0] 
		), .Z(n_98490351));
	notech_or4 i_17350(.A(n_124190608), .B(n_63762), .C(n_61775), .D(n_61953
		), .Z(n_98590352));
	notech_or4 i_17005(.A(n_314960777), .B(n_61065), .C(n_61052), .D(n_61837
		), .Z(n_113490501));
	notech_nao3 i_181772720(.A(n_579), .B(n_19698), .C(n_32484), .Z(n_113590502
		));
	notech_or4 i_6574529(.A(from_acu[0]), .B(from_acu[3]), .C(n_32934), .D(n_32933
		), .Z(n_114090507));
	notech_or4 i_6474530(.A(n_32934), .B(from_acu[3]), .C(from_acu[1]), .D(n_32932
		), .Z(n_114290509));
	notech_or4 i_831057(.A(from_acu[3]), .B(from_acu[2]), .C(from_acu[1]), .D
		(from_acu[0]), .Z(n_114590512));
	notech_or4 i_6374531(.A(from_acu[1]), .B(from_acu[0]), .C(from_acu[3]), 
		.D(n_30726), .Z(n_114790514));
	notech_or4 i_6274532(.A(from_acu[3]), .B(from_acu[2]), .C(n_32933), .D(n_32932
		), .Z(n_114990516));
	notech_or4 i_6074534(.A(from_acu[3]), .B(from_acu[2]), .C(n_32933), .D(from_acu
		[0]), .Z(n_115090517));
	notech_or4 i_5974535(.A(from_acu[3]), .B(from_acu[2]), .C(n_32932), .D(from_acu
		[1]), .Z(n_115190518));
	notech_and4 i_5774537(.A(from_acu[1]), .B(from_acu[0]), .C(from_acu[2]),
		 .D(n_32935), .Z(n_115290519));
	notech_ao4 i_172172816(.A(n_54271), .B(n_31882), .C(n_54153), .D(n_31658
		), .Z(n_115390520));
	notech_ao4 i_172072817(.A(n_54291), .B(n_31818), .C(n_54281), .D(n_31947
		), .Z(n_115490521));
	notech_ao4 i_171872819(.A(n_54311), .B(n_31423), .C(n_54301), .D(n_32011
		), .Z(n_115690523));
	notech_ao4 i_171772820(.A(n_54330), .B(n_31979), .C(n_31914), .D(n_54321
		), .Z(n_115790524));
	notech_ao4 i_171572822(.A(n_54271), .B(n_31883), .C(n_54153), .D(n_31659
		), .Z(n_115990526));
	notech_ao4 i_171472823(.A(n_54291), .B(n_31819), .C(n_54281), .D(n_31948
		), .Z(n_116090527));
	notech_ao4 i_171272825(.A(n_54311), .B(n_31424), .C(n_54301), .D(n_32012
		), .Z(n_116290529));
	notech_ao4 i_171172826(.A(n_54330), .B(n_31980), .C(n_31915), .D(n_54321
		), .Z(n_116390530));
	notech_ao4 i_170372834(.A(n_54271), .B(n_31885), .C(n_54153), .D(n_31661
		), .Z(n_116590532));
	notech_ao4 i_170272835(.A(n_54291), .B(n_31821), .C(n_54281), .D(n_31950
		), .Z(n_116690533));
	notech_ao4 i_170072837(.A(n_54311), .B(n_31426), .C(n_54301), .D(n_32014
		), .Z(n_116890535));
	notech_ao4 i_169972838(.A(n_54330), .B(n_31982), .C(n_31917), .D(n_54321
		), .Z(n_116990536));
	notech_ao4 i_169772840(.A(n_54271), .B(n_31886), .C(n_54153), .D(n_31662
		), .Z(n_117190538));
	notech_ao4 i_169672841(.A(n_54291), .B(n_31822), .C(n_54281), .D(n_31951
		), .Z(n_117290539));
	notech_ao4 i_169472843(.A(n_54311), .B(n_31427), .C(n_54301), .D(n_32015
		), .Z(n_117490541));
	notech_ao4 i_169372844(.A(n_54330), .B(n_31983), .C(n_31918), .D(n_54321
		), .Z(n_117590542));
	notech_ao4 i_169172846(.A(n_54270), .B(n_31887), .C(n_54152), .D(n_31663
		), .Z(n_117790544));
	notech_ao4 i_169072847(.A(n_54290), .B(n_31823), .C(n_54280), .D(n_31952
		), .Z(n_117890545));
	notech_ao4 i_168872849(.A(n_54310), .B(n_31428), .C(n_54300), .D(n_32016
		), .Z(n_118090547));
	notech_ao4 i_168772850(.A(n_54329), .B(n_31984), .C(n_31919), .D(n_54320
		), .Z(n_118190548));
	notech_ao4 i_168572852(.A(n_54270), .B(n_31888), .C(n_54152), .D(n_31664
		), .Z(n_118390550));
	notech_ao4 i_168472853(.A(n_54290), .B(n_31824), .C(n_54280), .D(n_31953
		), .Z(n_118490551));
	notech_ao4 i_168272855(.A(n_54310), .B(n_31429), .C(n_54300), .D(n_32017
		), .Z(n_118690553));
	notech_ao4 i_168172856(.A(n_54329), .B(n_31985), .C(n_31920), .D(n_54320
		), .Z(n_118790554));
	notech_ao4 i_136073177(.A(n_293792280), .B(n_31261), .C(n_57436), .D(n_30967
		), .Z(n_118990556));
	notech_ao4 i_135973178(.A(n_292192264), .B(n_101142452), .C(n_292292265)
		, .D(n_31294), .Z(n_119090557));
	notech_ao4 i_135873179(.A(n_293792280), .B(n_31262), .C(n_57436), .D(n_30969
		), .Z(n_119190558));
	notech_ao4 i_135773180(.A(n_334360971), .B(n_292192264), .C(n_292292265)
		, .D(n_31295), .Z(n_119290559));
	notech_ao4 i_135673181(.A(n_293792280), .B(n_31263), .C(n_57436), .D(n_30971
		), .Z(n_119390560));
	notech_ao4 i_135573182(.A(n_292192264), .B(n_100842449), .C(n_292292265)
		, .D(n_31296), .Z(n_119490561));
	notech_ao4 i_135473183(.A(n_293792280), .B(n_31264), .C(n_57436), .D(n_30973
		), .Z(n_119590562));
	notech_ao4 i_135373184(.A(n_338361011), .B(n_292192264), .C(n_292292265)
		, .D(n_31297), .Z(n_119690563));
	notech_ao4 i_135273185(.A(n_293792280), .B(n_31265), .C(n_57436), .D(n_30975
		), .Z(n_119790564));
	notech_ao4 i_135173186(.A(n_292192264), .B(n_334660974), .C(n_292292265)
		, .D(n_31298), .Z(n_119890565));
	notech_ao4 i_135073187(.A(n_293792280), .B(n_31266), .C(n_57436), .D(n_30977
		), .Z(n_119990566));
	notech_ao4 i_134973188(.A(n_292192264), .B(n_334860976), .C(n_292292265)
		, .D(n_31299), .Z(n_120090567));
	notech_ao4 i_134873189(.A(n_293792280), .B(n_31267), .C(n_57436), .D(n_30979
		), .Z(n_120190568));
	notech_ao4 i_134773190(.A(n_292192264), .B(n_100542446), .C(n_292292265)
		, .D(n_31300), .Z(n_120290569));
	notech_ao4 i_134673191(.A(n_293792280), .B(n_31268), .C(n_57423), .D(n_30981
		), .Z(n_120390570));
	notech_ao4 i_134573192(.A(n_292192264), .B(n_100242443), .C(n_292292265)
		, .D(n_31301), .Z(n_120490571));
	notech_ao4 i_134473193(.A(n_293792280), .B(n_31269), .C(n_57423), .D(n_30983
		), .Z(n_120590572));
	notech_ao4 i_134373194(.A(n_5269), .B(n_292192264), .C(n_292292265), .D(n_31302
		), .Z(n_120690573));
	notech_ao4 i_134273195(.A(n_293792280), .B(n_31270), .C(n_57423), .D(n_30985
		), .Z(n_120790574));
	notech_ao4 i_134173196(.A(n_99942440), .B(n_292192264), .C(n_292292265),
		 .D(n_31303), .Z(n_120890575));
	notech_ao4 i_133273205(.A(n_293792280), .B(n_31275), .C(n_57423), .D(n_30995
		), .Z(n_120990576));
	notech_ao4 i_133173206(.A(n_97342414), .B(n_292192264), .C(n_292292265),
		 .D(n_31308), .Z(n_121090577));
	notech_ao4 i_132873209(.A(n_293792280), .B(n_31277), .C(n_57423), .D(n_30999
		), .Z(n_121190578));
	notech_ao4 i_132773210(.A(n_292192264), .B(n_5444), .C(n_292292265), .D(n_31310
		), .Z(n_121290579));
	notech_ao4 i_132673211(.A(n_55207), .B(n_31278), .C(n_57423), .D(n_31002
		), .Z(n_121390580));
	notech_ao4 i_132573212(.A(n_55227), .B(n_5397), .C(n_55218), .D(n_31311)
		, .Z(n_121490581));
	notech_ao4 i_132473213(.A(n_55207), .B(n_31279), .C(n_57423), .D(n_31004
		), .Z(n_121590582));
	notech_ao4 i_132373214(.A(n_55227), .B(n_5436), .C(n_55218), .D(n_31312)
		, .Z(n_121690583));
	notech_ao4 i_132273215(.A(n_55207), .B(n_31280), .C(n_57423), .D(n_31006
		), .Z(n_121790584));
	notech_ao4 i_132173216(.A(n_55227), .B(n_5356), .C(n_55218), .D(n_31313)
		, .Z(n_121890585));
	notech_ao4 i_132073217(.A(n_55207), .B(n_31281), .C(n_57423), .D(n_31008
		), .Z(n_121990586));
	notech_ao4 i_131973218(.A(n_55227), .B(n_59466), .C(n_55218), .D(n_31314
		), .Z(n_122090587));
	notech_ao4 i_131873219(.A(n_55207), .B(n_31282), .C(n_57423), .D(n_31010
		), .Z(n_122190588));
	notech_ao4 i_131773220(.A(n_55227), .B(n_59465), .C(n_55218), .D(n_31315
		), .Z(n_122290589));
	notech_ao4 i_131673221(.A(n_55207), .B(n_31283), .C(n_57423), .D(n_31012
		), .Z(n_122390590));
	notech_ao4 i_131573222(.A(n_55227), .B(n_59464), .C(n_55218), .D(n_31316
		), .Z(n_122490591));
	notech_ao4 i_131473223(.A(n_55207), .B(n_31284), .C(n_57423), .D(n_31014
		), .Z(n_122590592));
	notech_ao4 i_131373224(.A(n_55227), .B(n_109226419), .C(n_55218), .D(n_31317
		), .Z(n_122690593));
	notech_ao4 i_131273225(.A(n_31285), .B(n_55207), .C(n_31016), .D(n_57423
		), .Z(n_122790594));
	notech_ao4 i_131173226(.A(n_106826395), .B(n_55227), .C(n_55218), .D(n_31318
		), .Z(n_122890595));
	notech_ao4 i_131073227(.A(n_55207), .B(n_31286), .C(n_57423), .D(n_31018
		), .Z(n_122990596));
	notech_ao4 i_130973228(.A(n_101026337), .B(n_55227), .C(n_55218), .D(n_31319
		), .Z(n_123090597));
	notech_ao4 i_130873229(.A(n_55207), .B(n_31287), .C(n_57423), .D(n_31020
		), .Z(n_123190598));
	notech_ao4 i_130773230(.A(n_55227), .B(n_5720), .C(n_55218), .D(n_31320)
		, .Z(n_123290599));
	notech_ao4 i_130673231(.A(n_55207), .B(n_31288), .C(n_57423), .D(n_31022
		), .Z(n_123390600));
	notech_ao4 i_130573232(.A(n_55227), .B(n_5711), .C(n_292292265), .D(n_31321
		), .Z(n_123490601));
	notech_ao4 i_130473233(.A(n_55207), .B(n_31289), .C(n_57423), .D(n_31024
		), .Z(n_123590602));
	notech_ao4 i_130373234(.A(n_55227), .B(n_4427), .C(n_55218), .D(n_31322)
		, .Z(n_123690603));
	notech_ao4 i_130073237(.A(n_55207), .B(n_31292), .C(n_57423), .D(n_31030
		), .Z(n_123790604));
	notech_ao4 i_129973238(.A(n_55227), .B(n_5243), .C(n_55218), .D(n_31325)
		, .Z(n_123890605));
	notech_or4 i_79474516(.A(n_32184), .B(n_61837), .C(n_32576), .D(n_63800)
		, .Z(n_124190608));
	notech_or4 i_195174502(.A(n_61739), .B(n_25713), .C(n_61609), .D(n_61864
		), .Z(n_124890615));
	notech_nao3 i_30171964(.A(n_195191311), .B(n_316260790), .C(n_61877), .Z
		(n_125190618));
	notech_or2 i_5571909(.A(n_28092), .B(n_28097), .Z(n_125290619));
	notech_or4 i_8271882(.A(n_61877), .B(n_61711), .C(n_61864), .D(n_57799),
		 .Z(n_125390620));
	notech_ao3 i_8371881(.A(n_61085), .B(n_61651), .C(n_315892477), .Z(n_125490621
		));
	notech_or4 i_46921(.A(n_30669), .B(n_30722), .C(n_125490621), .D(n_30670
		), .Z(n_8555));
	notech_ao3 i_8671878(.A(n_1836), .B(n_19680), .C(n_2091), .Z(n_125590622
		));
	notech_or4 i_47832(.A(n_2004), .B(n_30669), .C(n_30722), .D(n_125590622)
		, .Z(n_10020));
	notech_or4 i_29071689(.A(n_314960777), .B(n_61065), .C(n_61837), .D(n_60154
		), .Z(n_125690623));
	notech_nand2 i_29271687(.A(n_4401), .B(n_30648), .Z(n_125790624));
	notech_or4 i_29371686(.A(n_61877), .B(n_61717), .C(n_61864), .D(n_125990626
		), .Z(n_125890625));
	notech_and3 i_29171688(.A(n_32590), .B(n_1817), .C(n_125790624), .Z(n_125990626
		));
	notech_nao3 i_46995(.A(n_125690623), .B(n_125890625), .C(n_30722), .Z(\nbus_11285[0] 
		));
	notech_nand3 i_29571684(.A(n_284331524), .B(n_194984376), .C(n_295192294
		), .Z(n_126090627));
	notech_and2 i_30071679(.A(n_126290629), .B(eval_flag), .Z(n_126190628)
		);
	notech_nand2 i_29671683(.A(n_2036), .B(n_125390620), .Z(n_126290629));
	notech_nor2 i_29871681(.A(n_28007), .B(n_2152), .Z(n_126390630));
	notech_and3 i_29971680(.A(n_61085), .B(n_61651), .C(n_126090627), .Z(n_126490631
		));
	notech_or4 i_48586(.A(n_126390630), .B(n_30670), .C(n_126490631), .D(n_126190628
		), .Z(n_11366));
	notech_or4 i_44771533(.A(n_314960777), .B(n_61739), .C(n_2152), .D(n_27842
		), .Z(n_126590632));
	notech_or4 i_44671534(.A(n_32628), .B(n_32394), .C(n_61837), .D(n_60154)
		, .Z(n_126690633));
	notech_nand3 i_52234(.A(n_223991593), .B(n_126690633), .C(n_126590632), 
		.Z(n_16830));
	notech_or4 i_46071520(.A(n_61718), .B(n_61878), .C(n_61864), .D(n_363850921
		), .Z(n_126790634));
	notech_nao3 i_46178(.A(n_126790634), .B(n_364350916), .C(n_30722), .Z(n_7370
		));
	notech_nao3 i_46471516(.A(over_seg[5]), .B(n_61275), .C(n_348071366), .Z
		(n_126890635));
	notech_and2 i_46371517(.A(n_348171367), .B(n_126890635), .Z(n_127190638)
		);
	notech_ao4 i_53032(.A(n_61837), .B(n_127190638), .C(n_83245324), .D(n_57717
		), .Z(n_18288));
	notech_ao4 i_52988(.A(n_348489366), .B(n_30383), .C(n_348689368), .D(n_118487111
		), .Z(\nbus_11345[0] ));
	notech_or4 i_49371487(.A(n_32628), .B(n_32394), .C(n_60189), .D(n_61837)
		, .Z(n_127390640));
	notech_nao3 i_50732(.A(n_125690623), .B(n_127390640), .C(n_30722), .Z(n_14262
		));
	notech_or2 i_49671484(.A(n_2091), .B(n_30867), .Z(n_127490641));
	notech_nand3 i_48555(.A(n_2018), .B(n_53429), .C(n_127490641), .Z(n_11332
		));
	notech_or4 i_46258(.A(n_30671), .B(n_30722), .C(n_53445), .D(n_30672), .Z
		(\nbus_11272[0] ));
	notech_and2 i_54971431(.A(imm[8]), .B(n_57236), .Z(n_127590642));
	notech_and2 i_55171429(.A(imm[9]), .B(n_57236), .Z(n_127690643));
	notech_and2 i_55371427(.A(imm[10]), .B(n_57236), .Z(n_127790644));
	notech_and2 i_56371417(.A(imm[15]), .B(n_57236), .Z(n_127890645));
	notech_mux2 i_3878(.S(n_61651), .A(n_19680), .B(n_30651), .Z(n_10023));
	notech_xor2 i_58771393(.A(pipe_mul[0]), .B(pipe_mul[1]), .Z(n_128090647)
		);
	notech_nao3 i_59671384(.A(n_545), .B(mul64[31]), .C(n_61052), .Z(n_128690653
		));
	notech_nao3 i_59771383(.A(n_541), .B(mul64[7]), .C(n_60189), .Z(n_128790654
		));
	notech_nand2 i_60171379(.A(n_537), .B(n_30667), .Z(n_128890655));
	notech_ao4 i_5471910(.A(n_60189), .B(mul64[7]), .C(\opcode[1] ), .D(n_63762
		), .Z(n_128990656));
	notech_or4 i_60371377(.A(n_151990886), .B(n_151690883), .C(n_152890895),
		 .D(n_151390880), .Z(n_129090657));
	notech_ao4 i_1071954(.A(n_61052), .B(mul64[31]), .C(n_63762), .D(n_61953
		), .Z(n_129190658));
	notech_ao4 i_59371387(.A(n_1858), .B(mul64[15]), .C(n_32627), .D(n_315160779
		), .Z(n_129290659));
	notech_or4 i_63771344(.A(n_312460752), .B(n_2952), .C(n_61065), .D(n_129490661
		), .Z(n_129390660));
	notech_and4 i_60271378(.A(n_128790654), .B(n_128690653), .C(n_128890655)
		, .D(n_129090657), .Z(n_129490661));
	notech_nand2 i_6287(.A(n_129390660), .B(n_153190898), .Z(n_8438));
	notech_ao4 i_3215646(.A(n_249536174), .B(n_31539), .C(n_194891308), .D(n_31963
		), .Z(n_14492));
	notech_ao4 i_3115645(.A(n_249536174), .B(n_31538), .C(n_194891308), .D(n_31962
		), .Z(n_14487));
	notech_ao4 i_2915643(.A(n_249536174), .B(n_31536), .C(n_194891308), .D(n_31960
		), .Z(n_14477));
	notech_ao4 i_2815642(.A(n_249536174), .B(n_31535), .C(n_194891308), .D(n_31959
		), .Z(n_14472));
	notech_ao4 i_2715641(.A(n_249536174), .B(n_31534), .C(n_194891308), .D(n_31958
		), .Z(n_14467));
	notech_ao4 i_2615640(.A(n_249536174), .B(n_31533), .C(n_194891308), .D(n_31957
		), .Z(n_14462));
	notech_ao4 i_2515639(.A(n_249536174), .B(n_31532), .C(n_194891308), .D(n_31956
		), .Z(n_14457));
	notech_ao4 i_2415638(.A(n_249536174), .B(n_31531), .C(n_194891308), .D(n_31955
		), .Z(n_14452));
	notech_ao4 i_2315637(.A(n_249536174), .B(n_31530), .C(n_194891308), .D(n_31954
		), .Z(n_14447));
	notech_ao4 i_2215636(.A(n_249536174), .B(n_31529), .C(n_194891308), .D(n_31953
		), .Z(n_14442));
	notech_ao4 i_2115635(.A(n_249536174), .B(n_31528), .C(n_194891308), .D(n_31952
		), .Z(n_14437));
	notech_ao4 i_2015634(.A(n_249536174), .B(n_31527), .C(n_194891308), .D(n_31951
		), .Z(n_14432));
	notech_ao4 i_1815632(.A(n_249536174), .B(n_31525), .C(n_194891308), .D(n_31949
		), .Z(n_14422));
	notech_ao4 i_1715631(.A(n_249536174), .B(n_31524), .C(n_194891308), .D(n_31948
		), .Z(n_14417));
	notech_ao4 i_1615630(.A(n_249536174), .B(n_31523), .C(n_194891308), .D(n_31947
		), .Z(n_14412));
	notech_ao4 i_1515629(.A(n_55588), .B(n_31522), .C(n_55579), .D(n_31946),
		 .Z(n_14407));
	notech_ao4 i_1415628(.A(n_55588), .B(n_31521), .C(n_55579), .D(n_31945),
		 .Z(n_14402));
	notech_ao4 i_1315627(.A(n_55588), .B(n_31520), .C(n_55579), .D(n_31944),
		 .Z(n_14397));
	notech_ao4 i_1215626(.A(n_55588), .B(n_31519), .C(n_55579), .D(n_31943),
		 .Z(n_14392));
	notech_ao4 i_1115625(.A(n_55588), .B(n_31518), .C(n_55579), .D(n_31941),
		 .Z(n_14387));
	notech_ao4 i_1015624(.A(n_55588), .B(n_31517), .C(n_55579), .D(n_31940),
		 .Z(n_14382));
	notech_ao4 i_915623(.A(n_55588), .B(n_31516), .C(n_55579), .D(n_31939), 
		.Z(n_14377));
	notech_ao4 i_815622(.A(n_55588), .B(n_31515), .C(n_55579), .D(n_31938), 
		.Z(n_14372));
	notech_ao4 i_715621(.A(n_55588), .B(n_31514), .C(n_55579), .D(n_31937), 
		.Z(n_14367));
	notech_ao4 i_615620(.A(n_55588), .B(n_31513), .C(n_55579), .D(n_31936), 
		.Z(n_14362));
	notech_ao4 i_515619(.A(n_55588), .B(n_31512), .C(n_194891308), .D(n_31935
		), .Z(n_14357));
	notech_ao4 i_415618(.A(n_55588), .B(n_31511), .C(n_31934), .D(n_55579), 
		.Z(n_14352));
	notech_ao4 i_315617(.A(n_55588), .B(n_31510), .C(n_55579), .D(n_31933), 
		.Z(n_14347));
	notech_ao4 i_215616(.A(n_55588), .B(n_31509), .C(n_55579), .D(n_31932), 
		.Z(n_14342));
	notech_ao4 i_115615(.A(n_55579), .B(n_31931), .C(n_55588), .D(n_31508), 
		.Z(n_14337));
	notech_nand2 i_3127498(.A(n_153390900), .B(n_153290899), .Z(n_7934));
	notech_nand2 i_1827485(.A(n_153590902), .B(n_153490901), .Z(n_7869));
	notech_nand2 i_1527482(.A(n_153790904), .B(n_153690903), .Z(n_7854));
	notech_nand2 i_1127478(.A(n_153990906), .B(n_153890905), .Z(n_7834));
	notech_nand2 i_1027477(.A(n_154190908), .B(n_154090907), .Z(n_7829));
	notech_nand2 i_927476(.A(n_154390910), .B(n_154290909), .Z(n_7824));
	notech_nand2 i_827475(.A(n_154590912), .B(n_154490911), .Z(n_7819));
	notech_nand2 i_727474(.A(n_154790914), .B(n_154690913), .Z(n_7814));
	notech_nand2 i_227469(.A(n_154990916), .B(n_154890915), .Z(n_7789));
	notech_nand2 i_81271171(.A(divr_1[61]), .B(n_61609), .Z(n_139390760));
	notech_nand2 i_6227401(.A(n_155090917), .B(n_139390760), .Z(n_16807));
	notech_nand2 i_81771166(.A(divr_1[60]), .B(n_61609), .Z(n_139690763));
	notech_nand2 i_6127400(.A(n_155190918), .B(n_139690763), .Z(n_16802));
	notech_nand2 i_82271161(.A(divr_1[59]), .B(n_61609), .Z(n_139990766));
	notech_nand2 i_6027399(.A(n_155290919), .B(n_139990766), .Z(n_16797));
	notech_nand2 i_82771156(.A(divr_1[58]), .B(n_61609), .Z(n_140290769));
	notech_nand2 i_5927398(.A(n_155390920), .B(n_140290769), .Z(n_16792));
	notech_nand2 i_83271151(.A(divr_1[57]), .B(n_61609), .Z(n_140590772));
	notech_nand2 i_5827397(.A(n_155490921), .B(n_140590772), .Z(n_16787));
	notech_nand2 i_83771146(.A(divr_1[56]), .B(n_61607), .Z(n_140890775));
	notech_nand2 i_5727396(.A(n_155590922), .B(n_140890775), .Z(n_16782));
	notech_nand2 i_84271141(.A(divr_1[55]), .B(n_61607), .Z(n_141190778));
	notech_nand2 i_5627395(.A(n_155690923), .B(n_141190778), .Z(n_16777));
	notech_nand2 i_84771136(.A(divr_1[54]), .B(n_61607), .Z(n_141490781));
	notech_nand2 i_5527394(.A(n_155790924), .B(n_141490781), .Z(n_16772));
	notech_nand2 i_85271131(.A(divr_1[52]), .B(n_61609), .Z(n_141790784));
	notech_nand2 i_5327392(.A(n_155890925), .B(n_141790784), .Z(n_16762));
	notech_nand2 i_85771126(.A(divr_1[51]), .B(n_61609), .Z(n_142090787));
	notech_nand2 i_5227391(.A(n_155990926), .B(n_142090787), .Z(n_16757));
	notech_nand2 i_86771116(.A(divr_1[49]), .B(n_61609), .Z(n_142390790));
	notech_nand2 i_5027389(.A(n_156090927), .B(n_142390790), .Z(n_16747));
	notech_nand2 i_87271111(.A(divr_1[48]), .B(n_61618), .Z(n_142690793));
	notech_nand2 i_4927388(.A(n_156190928), .B(n_142690793), .Z(n_16742));
	notech_nand2 i_87771106(.A(divr_1[47]), .B(n_61618), .Z(n_142990796));
	notech_nand2 i_4827387(.A(n_156290929), .B(n_142990796), .Z(n_16737));
	notech_nand2 i_88271101(.A(divr_1[45]), .B(n_61618), .Z(n_143290799));
	notech_nand2 i_4627385(.A(n_156390930), .B(n_143290799), .Z(n_16727));
	notech_nand2 i_88771096(.A(divr_1[44]), .B(n_61618), .Z(n_143590802));
	notech_nand2 i_4527384(.A(n_156490931), .B(n_143590802), .Z(n_16722));
	notech_or2 i_12571980(.A(n_127890645), .B(n_57024), .Z(\nbus_11309[15] )
		);
	notech_nand2 i_104970934(.A(add_src[15]), .B(n_30668), .Z(n_143890805)
		);
	notech_ao4 i_104870935(.A(n_57024), .B(n_127890645), .C(n_56321), .D(n_349385901
		), .Z(n_144790814));
	notech_nao3 i_1612910(.A(n_157190938), .B(n_143890805), .C(n_144790814),
		 .Z(n_21382));
	notech_or2 i_20571985(.A(n_127790644), .B(n_57024), .Z(\nbus_11309[10] )
		);
	notech_nand2 i_114470839(.A(add_src[10]), .B(n_30668), .Z(n_144890815)
		);
	notech_ao4 i_114370840(.A(n_57024), .B(n_127790644), .C(n_56321), .D(n_349385901
		), .Z(n_145790824));
	notech_nao3 i_1112905(.A(n_157990946), .B(n_144890815), .C(n_145790824),
		 .Z(n_21357));
	notech_or2 i_20371986(.A(n_127690643), .B(n_57024), .Z(\nbus_11309[9] )
		);
	notech_nand2 i_116370820(.A(add_src[9]), .B(n_30668), .Z(n_145890825));
	notech_ao4 i_116270821(.A(n_57020), .B(n_127690643), .C(n_56321), .D(n_349385901
		), .Z(n_146790834));
	notech_nao3 i_1012904(.A(n_158790954), .B(n_145890825), .C(n_146790834),
		 .Z(n_21352));
	notech_or2 i_19171987(.A(n_127590642), .B(n_57020), .Z(\nbus_11309[8] )
		);
	notech_nand2 i_118270801(.A(add_src[8]), .B(n_30668), .Z(n_146890835));
	notech_ao4 i_118170802(.A(n_127590642), .B(n_57020), .C(n_56321), .D(n_349385901
		), .Z(n_147790844));
	notech_nao3 i_912903(.A(n_159590962), .B(n_146890835), .C(n_147790844), 
		.Z(n_21347));
	notech_or4 i_37833(.A(n_61837), .B(n_61824), .C(n_61797), .D(n_61775), .Z
		(n_149390860));
	notech_or4 i_62371358(.A(mul64[42]), .B(mul64[43]), .C(mul64[40]), .D(mul64
		[41]), .Z(n_150190868));
	notech_or4 i_62471357(.A(mul64[47]), .B(mul64[46]), .C(mul64[44]), .D(mul64
		[45]), .Z(n_150490871));
	notech_or4 i_62571356(.A(mul64[50]), .B(mul64[51]), .C(mul64[48]), .D(mul64
		[49]), .Z(n_150890875));
	notech_or4 i_62671355(.A(mul64[54]), .B(mul64[55]), .C(mul64[52]), .D(mul64
		[53]), .Z(n_151190878));
	notech_or4 i_63471347(.A(n_151190878), .B(n_150890875), .C(n_150490871),
		 .D(n_150190868), .Z(n_151390880));
	notech_or4 i_62771354(.A(mul64[58]), .B(mul64[59]), .C(mul64[56]), .D(mul64
		[57]), .Z(n_151690883));
	notech_or4 i_62871353(.A(mul64[62]), .B(mul64[63]), .C(mul64[60]), .D(mul64
		[61]), .Z(n_151990886));
	notech_and4 i_62171360(.A(n_33714), .B(n_33712), .C(n_33713), .D(n_33711
		), .Z(n_152390890));
	notech_or4 i_62271359(.A(mul64[38]), .B(mul64[39]), .C(mul64[37]), .D(mul64
		[36]), .Z(n_152690893));
	notech_nao3 i_63371348(.A(n_152390890), .B(n_30675), .C(n_129190658), .Z
		(n_152890895));
	notech_or4 i_63971342(.A(n_32589), .B(n_60189), .C(n_32627), .D(n_33754)
		, .Z(n_153090897));
	notech_ao4 i_64071341(.A(n_153090897), .B(n_33381), .C(n_129290659), .D(n_33717
		), .Z(n_153190898));
	notech_ao4 i_75071232(.A(n_309892426), .B(n_58992), .C(n_24298), .D(n_33718
		), .Z(n_153290899));
	notech_ao4 i_75171231(.A(n_59114), .B(n_32969), .C(n_56387), .D(n_32971)
		, .Z(n_153390900));
	notech_ao4 i_75771225(.A(n_309892426), .B(n_59086), .C(n_24298), .D(n_33719
		), .Z(n_153490901));
	notech_ao4 i_75871224(.A(n_59114), .B(n_32956), .C(n_56387), .D(n_32958)
		, .Z(n_153590902));
	notech_ao4 i_76471218(.A(n_309892426), .B(\nbus_11290[14] ), .C(n_24298)
		, .D(n_33720), .Z(n_153690903));
	notech_ao4 i_76571217(.A(n_59114), .B(n_32953), .C(n_56387), .D(n_32955)
		, .Z(n_153790904));
	notech_ao4 i_77171211(.A(n_309892426), .B(\nbus_11290[10] ), .C(n_24298)
		, .D(n_33721), .Z(n_153890905));
	notech_ao4 i_77271210(.A(n_59114), .B(n_32949), .C(n_56387), .D(n_32951)
		, .Z(n_153990906));
	notech_ao4 i_77971204(.A(n_309892426), .B(n_59032), .C(n_24298), .D(n_33722
		), .Z(n_154090907));
	notech_ao4 i_78071203(.A(n_59114), .B(n_32948), .C(n_56387), .D(n_32950)
		, .Z(n_154190908));
	notech_ao4 i_78671197(.A(n_309892426), .B(\nbus_11290[8] ), .C(n_24298),
		 .D(n_33723), .Z(n_154290909));
	notech_ao4 i_78771196(.A(n_59114), .B(n_32947), .C(n_56383), .D(n_32949)
		, .Z(n_154390910));
	notech_ao4 i_79371190(.A(n_309892426), .B(\nbus_11290[7] ), .C(n_24298),
		 .D(n_33724), .Z(n_154490911));
	notech_ao4 i_79471189(.A(n_59114), .B(n_32946), .C(n_56383), .D(n_32948)
		, .Z(n_154590912));
	notech_ao4 i_80071183(.A(n_309892426), .B(\nbus_11290[6] ), .C(n_24298),
		 .D(n_33725), .Z(n_154690913));
	notech_ao4 i_80171182(.A(n_59114), .B(n_32945), .C(n_56383), .D(n_32947)
		, .Z(n_154790914));
	notech_ao4 i_80771176(.A(n_309892426), .B(n_59005), .C(n_24298), .D(n_33726
		), .Z(n_154890915));
	notech_ao4 i_80871175(.A(n_59115), .B(n_32940), .C(n_56387), .D(n_32942)
		, .Z(n_154990916));
	notech_ao4 i_81371170(.A(n_24216), .B(n_33727), .C(n_56411), .D(n_60620)
		, .Z(n_155090917));
	notech_ao4 i_81871165(.A(n_24216), .B(n_33728), .C(n_56411), .D(nbus_11271
		[28]), .Z(n_155190918));
	notech_ao4 i_82371160(.A(n_24216), .B(n_33729), .C(n_56411), .D(n_60573)
		, .Z(n_155290919));
	notech_ao4 i_82871155(.A(n_24216), .B(n_33730), .C(n_56411), .D(n_60582)
		, .Z(n_155390920));
	notech_ao4 i_83371150(.A(n_24216), .B(n_33731), .C(n_56411), .D(n_60510)
		, .Z(n_155490921));
	notech_ao4 i_83871145(.A(n_24216), .B(n_33732), .C(n_56412), .D(n_60519)
		, .Z(n_155590922));
	notech_ao4 i_84371140(.A(n_24216), .B(n_33733), .C(n_56412), .D(n_60528)
		, .Z(n_155690923));
	notech_ao4 i_84871135(.A(n_24216), .B(n_33734), .C(n_56412), .D(nbus_11271
		[22]), .Z(n_155790924));
	notech_ao4 i_85371130(.A(n_24216), .B(n_33735), .C(n_56412), .D(nbus_11271
		[20]), .Z(n_155890925));
	notech_ao4 i_85871125(.A(n_24216), .B(n_33736), .C(n_56412), .D(nbus_11271
		[19]), .Z(n_155990926));
	notech_ao4 i_86871115(.A(n_24216), .B(n_33737), .C(n_56412), .D(nbus_11271
		[17]), .Z(n_156090927));
	notech_ao4 i_87371110(.A(n_24216), .B(n_33738), .C(n_56412), .D(nbus_11271
		[16]), .Z(n_156190928));
	notech_ao4 i_87871105(.A(n_24216), .B(n_33739), .C(n_56412), .D(nbus_11271
		[15]), .Z(n_156290929));
	notech_ao4 i_88371100(.A(n_24216), .B(n_33740), .C(n_56412), .D(nbus_11271
		[13]), .Z(n_156390930));
	notech_ao4 i_88871095(.A(n_24216), .B(n_33741), .C(n_56412), .D(nbus_11271
		[12]), .Z(n_156490931));
	notech_ao4 i_105070933(.A(n_2129), .B(n_32896), .C(n_2128), .D(n_32867),
		 .Z(n_156590932));
	notech_ao4 i_105170932(.A(n_4350), .B(n_33743), .C(n_56330), .D(n_33742)
		, .Z(n_156690933));
	notech_ao4 i_105270931(.A(n_4353), .B(nbus_11271[15]), .C(n_24142), .D(n_33744
		), .Z(n_156890935));
	notech_ao4 i_105370930(.A(n_2127), .B(n_31523), .C(n_4352), .D(n_58348),
		 .Z(n_156990936));
	notech_and4 i_105670927(.A(n_156990936), .B(n_156890935), .C(n_156690933
		), .D(n_156590932), .Z(n_157190938));
	notech_ao4 i_114570838(.A(n_2129), .B(n_32891), .C(n_2128), .D(n_32862),
		 .Z(n_157390940));
	notech_ao4 i_114670837(.A(n_56359), .B(nbus_11271[10]), .C(n_56330), .D(n_33745
		), .Z(n_157490941));
	notech_ao4 i_114770836(.A(n_56718), .B(n_33747), .C(n_56341), .D(n_33746
		), .Z(n_157690943));
	notech_ao4 i_114870835(.A(n_2127), .B(n_31518), .C(n_56350), .D(n_58303)
		, .Z(n_157790944));
	notech_and4 i_115170832(.A(n_157790944), .B(n_157690943), .C(n_157490941
		), .D(n_157390940), .Z(n_157990946));
	notech_ao4 i_116470819(.A(n_2129), .B(n_32890), .C(n_2128), .D(n_32861),
		 .Z(n_158190948));
	notech_ao4 i_116570818(.A(n_56359), .B(nbus_11271[9]), .C(n_56330), .D(n_33748
		), .Z(n_158290949));
	notech_ao4 i_116670817(.A(n_56718), .B(n_33750), .C(n_56341), .D(n_33749
		), .Z(n_158490951));
	notech_ao4 i_116770816(.A(n_2127), .B(n_31517), .C(n_56350), .D(nbus_11273
		[9]), .Z(n_158590952));
	notech_and4 i_117070813(.A(n_158590952), .B(n_158490951), .C(n_158290949
		), .D(n_158190948), .Z(n_158790954));
	notech_ao4 i_118370800(.A(n_2129), .B(n_32889), .C(n_2128), .D(n_32860),
		 .Z(n_158990956));
	notech_ao4 i_118470799(.A(n_56359), .B(nbus_11271[8]), .C(n_56330), .D(n_33751
		), .Z(n_159090957));
	notech_ao4 i_118570798(.A(n_56718), .B(n_33753), .C(n_56341), .D(n_33752
		), .Z(n_159290959));
	notech_ao4 i_118670797(.A(n_2127), .B(n_31516), .C(n_56350), .D(n_58285)
		, .Z(n_159390960));
	notech_and4 i_118970794(.A(n_159390960), .B(n_159290959), .C(n_159090957
		), .D(n_158990956), .Z(n_159590962));
	notech_and2 i_15669109(.A(imm[29]), .B(n_57236), .Z(n_159890965));
	notech_nao3 i_134567991(.A(n_3584), .B(opb[31]), .C(n_56428), .Z(n_160090967
		));
	notech_nand2 i_3327500(.A(n_180191168), .B(n_160090967), .Z(n_7944));
	notech_nao3 i_135167985(.A(n_3583), .B(opb[31]), .C(n_56428), .Z(n_160390970
		));
	notech_or4 i_135067986(.A(n_61878), .B(n_2112), .C(n_61718), .D(n_58983)
		, .Z(n_160690973));
	notech_nand3 i_3227499(.A(n_180291169), .B(n_160690973), .C(n_160390970)
		, .Z(n_7939));
	notech_nao3 i_135867978(.A(n_3581), .B(opb[31]), .C(n_56428), .Z(n_160790974
		));
	notech_nor2 i_135767979(.A(n_59115), .B(n_32968), .Z(n_161090977));
	notech_nao3 i_3027497(.A(n_180491171), .B(n_160790974), .C(n_161090977),
		 .Z(n_7929));
	notech_nao3 i_136567971(.A(n_3580), .B(opb[31]), .C(n_56429), .Z(n_161190978
		));
	notech_nor2 i_136467972(.A(n_59115), .B(n_32967), .Z(n_161490981));
	notech_nao3 i_2927496(.A(n_180691173), .B(n_161190978), .C(n_161490981),
		 .Z(n_7924));
	notech_nao3 i_137267964(.A(n_3579), .B(opb[31]), .C(n_56429), .Z(n_161590982
		));
	notech_nor2 i_137167965(.A(n_59115), .B(n_32966), .Z(n_161890985));
	notech_nao3 i_2827495(.A(n_180891175), .B(n_161590982), .C(n_161890985),
		 .Z(n_7919));
	notech_nao3 i_137967957(.A(n_3578), .B(opb[31]), .C(n_56429), .Z(n_161990986
		));
	notech_nor2 i_137867958(.A(n_59115), .B(n_32965), .Z(n_162290989));
	notech_nao3 i_2727494(.A(n_181091177), .B(n_161990986), .C(n_162290989),
		 .Z(n_7914));
	notech_nao3 i_138667950(.A(n_3577), .B(opb[31]), .C(n_56429), .Z(n_162390990
		));
	notech_nor2 i_138567951(.A(n_59115), .B(n_32964), .Z(n_162690993));
	notech_nao3 i_2627493(.A(n_181291179), .B(n_162390990), .C(n_162690993),
		 .Z(n_7909));
	notech_nao3 i_139367943(.A(n_3576), .B(opb[31]), .C(n_56429), .Z(n_162790994
		));
	notech_nor2 i_139267944(.A(n_59115), .B(n_32963), .Z(n_163090997));
	notech_nao3 i_2527492(.A(n_181491181), .B(n_162790994), .C(n_163090997),
		 .Z(n_7904));
	notech_nao3 i_140067936(.A(n_3575), .B(opb[31]), .C(n_56429), .Z(n_163190998
		));
	notech_nor2 i_139967937(.A(n_59115), .B(n_32962), .Z(n_163491001));
	notech_nao3 i_2427491(.A(n_181891183), .B(n_163190998), .C(n_163491001),
		 .Z(n_7899));
	notech_nao3 i_140767929(.A(n_3574), .B(opb[31]), .C(n_56429), .Z(n_163591002
		));
	notech_nor2 i_140667930(.A(n_59115), .B(n_32961), .Z(n_163891005));
	notech_nao3 i_2327490(.A(n_182191185), .B(n_163591002), .C(n_163891005),
		 .Z(n_7894));
	notech_nao3 i_141467922(.A(n_3573), .B(opb[31]), .C(n_56429), .Z(n_163991006
		));
	notech_nor2 i_141367923(.A(n_59115), .B(n_32960), .Z(n_164291009));
	notech_nao3 i_2227489(.A(n_182391187), .B(n_163991006), .C(n_164291009),
		 .Z(n_7889));
	notech_nao3 i_142167915(.A(n_3572), .B(opb[31]), .C(n_56429), .Z(n_164391010
		));
	notech_nor2 i_142067916(.A(n_59115), .B(n_32959), .Z(n_164691013));
	notech_nao3 i_2127488(.A(n_182591189), .B(n_164391010), .C(n_164691013),
		 .Z(n_7884));
	notech_nao3 i_142867908(.A(n_3571), .B(opb[31]), .C(n_56429), .Z(n_164791014
		));
	notech_nor2 i_142767909(.A(n_59115), .B(n_32958), .Z(n_165091017));
	notech_nao3 i_2027487(.A(n_182791191), .B(n_164791014), .C(n_165091017),
		 .Z(n_7879));
	notech_nao3 i_143567901(.A(n_3570), .B(opb[31]), .C(n_56429), .Z(n_165191018
		));
	notech_nor2 i_143467902(.A(n_59115), .B(n_32957), .Z(n_165491021));
	notech_nao3 i_1927486(.A(n_182991193), .B(n_165191018), .C(n_165491021),
		 .Z(n_7874));
	notech_nao3 i_144267894(.A(n_3568), .B(n_60629), .C(n_56429), .Z(n_165591022
		));
	notech_nor2 i_144167895(.A(n_59115), .B(n_32955), .Z(n_165891025));
	notech_nao3 i_1727484(.A(n_183291195), .B(n_165591022), .C(n_165891025),
		 .Z(n_7864));
	notech_nao3 i_147467866(.A(n_3557), .B(n_60629), .C(n_56429), .Z(n_165991026
		));
	notech_nor2 i_147267867(.A(n_59115), .B(n_32944), .Z(n_166291029));
	notech_nao3 i_627473(.A(n_183491197), .B(n_165991026), .C(n_166291029), 
		.Z(n_7809));
	notech_nao3 i_148167859(.A(n_3556), .B(n_60629), .C(n_56429), .Z(n_166391030
		));
	notech_nor2 i_148067860(.A(n_59115), .B(n_32943), .Z(n_166691033));
	notech_nao3 i_527472(.A(n_183691199), .B(n_166391030), .C(n_166691033), 
		.Z(n_7804));
	notech_nao3 i_148867852(.A(n_3555), .B(n_60629), .C(n_56429), .Z(n_166791034
		));
	notech_nor2 i_148767853(.A(n_59115), .B(n_32942), .Z(n_167091037));
	notech_nao3 i_427471(.A(n_183891201), .B(n_166791034), .C(n_167091037), 
		.Z(n_7799));
	notech_nao3 i_149567845(.A(n_3554), .B(n_60629), .C(n_56429), .Z(n_167191038
		));
	notech_nor2 i_149467846(.A(n_59114), .B(n_32941), .Z(n_167491041));
	notech_nao3 i_327470(.A(n_184091203), .B(n_167191038), .C(n_167491041), 
		.Z(n_7794));
	notech_nao3 i_150267839(.A(n_3552), .B(n_60629), .C(n_56429), .Z(n_167591042
		));
	notech_nand2 i_127468(.A(n_184291205), .B(n_167591042), .Z(n_7784));
	notech_nao3 i_150767834(.A(n_3551), .B(n_60605), .C(n_56429), .Z(n_167891045
		));
	notech_nand2 i_6427403(.A(n_184391206), .B(n_167891045), .Z(n_16817));
	notech_nao3 i_151367829(.A(n_3550), .B(n_60605), .C(n_56429), .Z(n_168191048
		));
	notech_nand2 i_6327402(.A(n_184491207), .B(n_168191048), .Z(n_16812));
	notech_nao3 i_151867824(.A(n_3541), .B(n_60605), .C(n_56416), .Z(n_168491051
		));
	notech_nand2 i_5427393(.A(n_184591208), .B(n_168491051), .Z(n_16767));
	notech_nao3 i_152367819(.A(n_3534), .B(n_60607), .C(n_56416), .Z(n_168791054
		));
	notech_nand2 i_4727386(.A(n_184691209), .B(n_168791054), .Z(n_16732));
	notech_nao3 i_152867814(.A(n_3531), .B(n_60607), .C(n_56416), .Z(n_169091057
		));
	notech_nand2 i_4427383(.A(n_184791210), .B(n_169091057), .Z(n_16717));
	notech_nao3 i_153367809(.A(n_3530), .B(n_60607), .C(n_56416), .Z(n_169391060
		));
	notech_nand2 i_4327382(.A(n_184891211), .B(n_169391060), .Z(n_16712));
	notech_nao3 i_153967804(.A(n_3529), .B(n_60607), .C(n_56416), .Z(n_169691063
		));
	notech_nand2 i_4227381(.A(n_184991212), .B(n_169691063), .Z(n_16707));
	notech_nao3 i_154567799(.A(n_3528), .B(n_60607), .C(n_56422), .Z(n_169991066
		));
	notech_nand2 i_4127380(.A(n_185091213), .B(n_169991066), .Z(n_16702));
	notech_nao3 i_155067794(.A(n_3527), .B(n_60607), .C(n_56422), .Z(n_170291069
		));
	notech_nand2 i_4027379(.A(n_185191214), .B(n_170291069), .Z(n_16697));
	notech_nao3 i_155567789(.A(n_3526), .B(n_60607), .C(n_56422), .Z(n_170591072
		));
	notech_nand2 i_3927378(.A(n_185291215), .B(n_170591072), .Z(n_16692));
	notech_nao3 i_156067784(.A(n_3525), .B(n_60607), .C(n_56422), .Z(n_170891075
		));
	notech_nand2 i_3827377(.A(n_185391216), .B(n_170891075), .Z(n_16687));
	notech_nao3 i_156667779(.A(n_3524), .B(n_60607), .C(n_56416), .Z(n_171191078
		));
	notech_nand2 i_3727376(.A(n_185491217), .B(n_171191078), .Z(n_16682));
	notech_nao3 i_157267774(.A(n_3523), .B(n_60607), .C(n_56416), .Z(n_171491081
		));
	notech_nand2 i_3627375(.A(n_185591218), .B(n_171491081), .Z(n_16677));
	notech_nao3 i_157767769(.A(n_3522), .B(n_60607), .C(n_56416), .Z(n_171791084
		));
	notech_nand2 i_3527374(.A(n_185991219), .B(n_171791084), .Z(n_16672));
	notech_nao3 i_158367764(.A(n_3521), .B(n_60607), .C(n_56416), .Z(n_172091087
		));
	notech_nand2 i_3427373(.A(n_186091220), .B(n_172091087), .Z(n_16667));
	notech_nao3 i_159067759(.A(n_3520), .B(n_60607), .C(n_56416), .Z(n_172391090
		));
	notech_nand2 i_3327372(.A(n_186191221), .B(n_172391090), .Z(n_16662));
	notech_nao3 i_159667754(.A(n_3519), .B(n_60607), .C(n_56416), .Z(n_172691093
		));
	notech_nand2 i_3227371(.A(n_186291222), .B(n_172691093), .Z(n_16657));
	notech_nao3 i_160167749(.A(n_3518), .B(n_60600), .C(n_56416), .Z(n_172991096
		));
	notech_nand2 i_3127370(.A(n_186391223), .B(n_172991096), .Z(n_16652));
	notech_nao3 i_160667744(.A(n_3517), .B(n_60600), .C(n_56416), .Z(n_173291099
		));
	notech_nand2 i_3027369(.A(n_186491224), .B(n_173291099), .Z(n_16647));
	notech_nao3 i_161667734(.A(n_3515), .B(n_60600), .C(n_56416), .Z(n_173591102
		));
	notech_nand2 i_2827367(.A(n_186591225), .B(n_173591102), .Z(n_16637));
	notech_nao3 i_162667724(.A(n_3513), .B(n_60602), .C(n_56422), .Z(n_173891105
		));
	notech_nand2 i_2627365(.A(n_186691226), .B(n_173891105), .Z(n_16627));
	notech_nao3 i_164867704(.A(n_3509), .B(n_60602), .C(n_56422), .Z(n_174191108
		));
	notech_nand2 i_2227361(.A(n_186791227), .B(n_174191108), .Z(n_16607));
	notech_nao3 i_165367699(.A(n_3508), .B(n_60602), .C(n_56422), .Z(n_174491111
		));
	notech_nand2 i_2127360(.A(n_186891228), .B(n_174491111), .Z(n_16602));
	notech_nao3 i_165867694(.A(n_3507), .B(n_60600), .C(n_56422), .Z(n_174791114
		));
	notech_nand2 i_2027359(.A(n_186991229), .B(n_174791114), .Z(n_16597));
	notech_nao3 i_166367689(.A(n_3506), .B(n_60600), .C(n_56422), .Z(n_175091117
		));
	notech_nand2 i_1927358(.A(n_187091230), .B(n_175091117), .Z(n_16592));
	notech_nao3 i_166867684(.A(n_3505), .B(n_60600), .C(n_56422), .Z(n_175391120
		));
	notech_nand2 i_1827357(.A(n_187191231), .B(n_175391120), .Z(n_16587));
	notech_nao3 i_167467679(.A(n_3504), .B(n_60600), .C(n_56428), .Z(n_175691123
		));
	notech_nand2 i_1727356(.A(n_187291232), .B(n_175691123), .Z(n_16582));
	notech_nao3 i_168767669(.A(n_3502), .B(n_60600), .C(n_56428), .Z(n_175991126
		));
	notech_nand2 i_1527354(.A(n_187391233), .B(n_175991126), .Z(n_16572));
	notech_nao3 i_171467644(.A(n_3497), .B(n_60600), .C(n_56422), .Z(n_176291129
		));
	notech_nand2 i_1027349(.A(n_187491234), .B(n_176291129), .Z(n_16547));
	notech_nao3 i_171967639(.A(n_3496), .B(n_60602), .C(n_56428), .Z(n_176591132
		));
	notech_nand2 i_927348(.A(n_187591235), .B(n_176591132), .Z(n_16542));
	notech_nao3 i_172567634(.A(n_3495), .B(n_60602), .C(n_56422), .Z(n_176891135
		));
	notech_nand2 i_827347(.A(n_187691236), .B(n_176891135), .Z(n_16537));
	notech_nao3 i_173467629(.A(n_3494), .B(n_60602), .C(n_56422), .Z(n_177191138
		));
	notech_nand2 i_727346(.A(n_187791237), .B(n_177191138), .Z(n_16532));
	notech_nao3 i_173967624(.A(n_3493), .B(n_60605), .C(n_56422), .Z(n_177491141
		));
	notech_nand2 i_627345(.A(n_187891238), .B(n_177491141), .Z(n_16527));
	notech_nao3 i_174567619(.A(n_3492), .B(n_60602), .C(n_56422), .Z(n_177791144
		));
	notech_nand2 i_527344(.A(n_187991239), .B(n_177791144), .Z(n_16522));
	notech_nao3 i_175267614(.A(n_3491), .B(n_60602), .C(n_56422), .Z(n_178091147
		));
	notech_nand2 i_427343(.A(n_188091240), .B(n_178091147), .Z(n_16517));
	notech_nao3 i_175767609(.A(n_3490), .B(n_60602), .C(n_56422), .Z(n_178391150
		));
	notech_nand2 i_327342(.A(n_188191241), .B(n_178391150), .Z(n_16512));
	notech_nao3 i_176267604(.A(n_3489), .B(n_60602), .C(n_56422), .Z(n_178691153
		));
	notech_nand2 i_227341(.A(n_188291242), .B(n_178691153), .Z(n_16507));
	notech_nao3 i_177767589(.A(n_3488), .B(n_60602), .C(n_56422), .Z(n_178991156
		));
	notech_nand2 i_127340(.A(n_188391243), .B(n_178991156), .Z(n_16502));
	notech_ao4 i_180967557(.A(n_57024), .B(n_159890965), .C(n_56321), .D(n_384582276
		), .Z(n_179291159));
	notech_or2 i_19969316(.A(n_159890965), .B(n_57024), .Z(\nbus_11309[29] )
		);
	notech_nand2 i_3012924(.A(n_189091250), .B(n_30676), .Z(n_21452));
	notech_ao4 i_134667990(.A(n_59104), .B(n_32971), .C(n_56387), .D(n_32973
		), .Z(n_180191168));
	notech_ao4 i_135267984(.A(n_59104), .B(n_32970), .C(n_56387), .D(n_32972
		), .Z(n_180291169));
	notech_ao4 i_135967977(.A(n_56387), .B(n_32970), .C(n_309892426), .D(n_58947
		), .Z(n_180491171));
	notech_ao4 i_136667970(.A(n_56387), .B(n_32969), .C(n_309892426), .D(n_58929
		), .Z(n_180691173));
	notech_ao4 i_137367963(.A(n_56388), .B(n_32968), .C(n_309892426), .D(n_58938
		), .Z(n_180891175));
	notech_ao4 i_138067956(.A(n_56388), .B(n_32967), .C(n_309892426), .D(n_58911
		), .Z(n_181091177));
	notech_ao4 i_138767949(.A(n_56388), .B(n_32966), .C(n_56368), .D(n_58920
		), .Z(n_181291179));
	notech_ao4 i_139467942(.A(n_56388), .B(n_32965), .C(n_56368), .D(n_58893
		), .Z(n_181491181));
	notech_ao4 i_140167935(.A(n_56388), .B(n_32964), .C(n_56368), .D(n_58902
		), .Z(n_181891183));
	notech_ao4 i_140867928(.A(n_56388), .B(n_32963), .C(n_56368), .D(n_58875
		), .Z(n_182191185));
	notech_ao4 i_141567921(.A(n_56388), .B(n_32962), .C(n_56368), .D(n_58884
		), .Z(n_182391187));
	notech_ao4 i_142267914(.A(n_56388), .B(n_32961), .C(n_56368), .D(n_58857
		), .Z(n_182591189));
	notech_ao4 i_142967907(.A(n_56388), .B(n_32960), .C(n_56368), .D(n_58866
		), .Z(n_182791191));
	notech_ao4 i_143667900(.A(n_56388), .B(n_32959), .C(n_56368), .D(n_59077
		), .Z(n_182991193));
	notech_ao4 i_144367893(.A(n_56387), .B(n_32957), .C(n_56368), .D(n_59059
		), .Z(n_183291195));
	notech_ao4 i_147567865(.A(n_56388), .B(n_32946), .C(n_56368), .D(\nbus_11290[5] 
		), .Z(n_183491197));
	notech_ao4 i_148267858(.A(n_56388), .B(n_32945), .C(n_56368), .D(\nbus_11290[4] 
		), .Z(n_183691199));
	notech_ao4 i_148967851(.A(n_56388), .B(n_32944), .C(n_56368), .D(\nbus_11290[3] 
		), .Z(n_183891201));
	notech_ao4 i_149667844(.A(n_56388), .B(n_32943), .C(n_56368), .D(\nbus_11290[2] 
		), .Z(n_184091203));
	notech_ao4 i_150367838(.A(n_56368), .B(n_58956), .C(n_56383), .D(n_32941
		), .Z(n_184291205));
	notech_ao4 i_150867833(.A(n_309192421), .B(n_60591), .C(n_61651), .D(n_32645
		), .Z(n_184391206));
	notech_ao4 i_151467828(.A(n_56411), .B(n_60611), .C(n_61651), .D(n_32644
		), .Z(n_184491207));
	notech_ao4 i_151967823(.A(n_56412), .B(nbus_11271[21]), .C(n_61647), .D(n_32643
		), .Z(n_184591208));
	notech_ao4 i_152467818(.A(n_56412), .B(nbus_11271[14]), .C(n_61647), .D(n_32642
		), .Z(n_184691209));
	notech_ao4 i_152967813(.A(n_56412), .B(nbus_11271[11]), .C(n_61647), .D(n_32641
		), .Z(n_184791210));
	notech_ao4 i_153467808(.A(n_56412), .B(nbus_11271[10]), .C(n_61647), .D(n_32640
		), .Z(n_184891211));
	notech_ao4 i_154067803(.A(n_56407), .B(nbus_11271[9]), .C(n_61647), .D(n_32639
		), .Z(n_184991212));
	notech_ao4 i_154667798(.A(n_56404), .B(nbus_11271[8]), .C(n_61647), .D(n_32638
		), .Z(n_185091213));
	notech_ao4 i_155167793(.A(n_56404), .B(nbus_11271[7]), .C(n_61647), .D(n_32637
		), .Z(n_185191214));
	notech_ao4 i_155667788(.A(n_56404), .B(nbus_11271[6]), .C(n_61647), .D(n_32636
		), .Z(n_185291215));
	notech_ao4 i_156167783(.A(n_56404), .B(nbus_11271[5]), .C(n_61647), .D(n_32635
		), .Z(n_185391216));
	notech_ao4 i_156867778(.A(n_56404), .B(nbus_11271[4]), .C(n_61647), .D(n_32634
		), .Z(n_185491217));
	notech_ao4 i_157367773(.A(n_56404), .B(nbus_11271[3]), .C(n_61651), .D(n_32632
		), .Z(n_185591218));
	notech_ao4 i_157867768(.A(n_56404), .B(nbus_11271[2]), .C(n_61652), .D(n_32631
		), .Z(n_185991219));
	notech_ao4 i_158467763(.A(n_56404), .B(nbus_11271[1]), .C(n_61652), .D(n_32630
		), .Z(n_186091220));
	notech_ao4 i_159167758(.A(n_56403), .B(nbus_11271[0]), .C(n_61652), .D(n_32626
		), .Z(n_186191221));
	notech_ao4 i_159767753(.A(n_56403), .B(n_60458), .C(n_61652), .D(n_32625
		), .Z(n_186291222));
	notech_ao4 i_160267748(.A(n_56403), .B(n_58483), .C(n_61652), .D(n_32624
		), .Z(n_186391223));
	notech_ao4 i_160767743(.A(n_56403), .B(n_58474), .C(n_61656), .D(n_32623
		), .Z(n_186491224));
	notech_ao4 i_161767733(.A(n_56403), .B(n_58456), .C(n_61656), .D(n_32621
		), .Z(n_186591225));
	notech_ao4 i_162767723(.A(n_56403), .B(n_58438), .C(n_61652), .D(n_32619
		), .Z(n_186691226));
	notech_ao4 i_164967703(.A(n_56403), .B(n_58402), .C(n_61652), .D(n_32613
		), .Z(n_186791227));
	notech_ao4 i_165467698(.A(n_56404), .B(n_58393), .C(n_61652), .D(n_32612
		), .Z(n_186891228));
	notech_ao4 i_165967693(.A(n_56407), .B(n_58384), .C(n_61651), .D(n_32611
		), .Z(n_186991229));
	notech_ao4 i_166467688(.A(n_56407), .B(n_58375), .C(n_61652), .D(n_32610
		), .Z(n_187091230));
	notech_ao4 i_166967683(.A(n_56407), .B(n_58366), .C(n_61651), .D(n_32609
		), .Z(n_187191231));
	notech_ao4 i_167767678(.A(n_56407), .B(n_58357), .C(n_61651), .D(n_32608
		), .Z(n_187291232));
	notech_ao4 i_168867668(.A(n_56407), .B(n_58339), .C(n_61651), .D(n_32606
		), .Z(n_187391233));
	notech_ao4 i_171567643(.A(n_56407), .B(n_58294), .C(n_61652), .D(n_32601
		), .Z(n_187491234));
	notech_ao4 i_172067638(.A(n_56407), .B(n_58285), .C(n_61652), .D(n_32600
		), .Z(n_187591235));
	notech_ao4 i_173067633(.A(n_56407), .B(n_58275), .C(n_61652), .D(n_32599
		), .Z(n_187691236));
	notech_ao4 i_173567628(.A(n_56404), .B(nbus_11273[6]), .C(n_61652), .D(n_32598
		), .Z(n_187791237));
	notech_ao4 i_174067623(.A(n_56404), .B(nbus_11273[5]), .C(n_61652), .D(n_32597
		), .Z(n_187891238));
	notech_ao4 i_174667618(.A(n_56404), .B(nbus_11273[4]), .C(n_61647), .D(n_32596
		), .Z(n_187991239));
	notech_ao4 i_175367613(.A(n_56404), .B(n_58256), .C(n_61643), .D(n_32595
		), .Z(n_188091240));
	notech_ao4 i_175867608(.A(n_56407), .B(n_58247), .C(n_61643), .D(n_32594
		), .Z(n_188191241));
	notech_ao4 i_176367603(.A(n_56407), .B(n_58229), .C(n_61643), .D(n_32593
		), .Z(n_188291242));
	notech_ao4 i_177867588(.A(n_56404), .B(nbus_11273[0]), .C(n_61642), .D(n_32592
		), .Z(n_188391243));
	notech_ao4 i_181067556(.A(n_4348), .B(n_31537), .C(n_112042561), .D(n_32343
		), .Z(n_188491244));
	notech_ao4 i_181167555(.A(n_56359), .B(n_60620), .C(n_56330), .D(n_33755
		), .Z(n_188591245));
	notech_ao4 i_181267554(.A(n_56718), .B(n_33757), .C(n_56341), .D(n_33756
		), .Z(n_188791247));
	notech_ao4 i_181367553(.A(n_56350), .B(n_58474), .C(n_4351), .D(n_32910)
		, .Z(n_188891248));
	notech_and4 i_181667550(.A(n_188891248), .B(n_188791247), .C(n_188591245
		), .D(n_188491244), .Z(n_189091250));
	notech_ao4 i_11163246(.A(n_336760995), .B(n_57656), .C(n_56965), .D(n_331960947
		), .Z(n_189191251));
	notech_ao4 i_14863211(.A(nbus_11273[0]), .B(n_331860946), .C(n_58956), .D
		(n_189591255), .Z(n_189291252));
	notech_and4 i_14963210(.A(n_191391273), .B(n_191591275), .C(n_191491274)
		, .D(n_191691276), .Z(n_189391253));
	notech_and2 i_11063247(.A(n_57742), .B(n_1847), .Z(n_189591255));
	notech_nand2 i_12663233(.A(n_192091280), .B(n_189891258), .Z(n_189791257
		));
	notech_nand2 i_57662807(.A(n_30389), .B(\opa_12[0] ), .Z(n_189891258));
	notech_nand2 i_56762816(.A(regs_4_2[0]), .B(n_30359), .Z(n_190791267));
	notech_or4 i_56162821(.A(n_61838), .B(n_189391253), .C(n_339461022), .D(n_191791277
		), .Z(n_191291272));
	notech_nao3 i_57462809(.A(n_247980969), .B(opb[0]), .C(n_26618), .Z(n_191391273
		));
	notech_nand3 i_57562808(.A(n_247980969), .B(n_30389), .C(opa[0]), .Z(n_191491274
		));
	notech_or4 i_57262811(.A(n_56002), .B(n_331960947), .C(n_61933), .D(nbus_11271
		[0]), .Z(n_191591275));
	notech_nand2 i_57362810(.A(n_32323), .B(n_189791257), .Z(n_191691276));
	notech_and2 i_2563332(.A(n_63800), .B(n_32215), .Z(n_191791277));
	notech_ao4 i_12063239(.A(n_327760905), .B(n_56002), .C(n_101142452), .D(n_26618
		), .Z(n_192091280));
	notech_or4 i_132762084(.A(n_61841), .B(n_339461022), .C(n_61824), .D(n_57199
		), .Z(n_192391283));
	notech_ao4 i_132162090(.A(n_61841), .B(n_189291252), .C(n_189191251), .D
		(n_192391283), .Z(n_192491284));
	notech_ao4 i_132062091(.A(n_101142452), .B(n_332660954), .C(n_33169), .D
		(n_332360951), .Z(n_192691286));
	notech_and3 i_132362088(.A(n_191291272), .B(n_192491284), .C(n_192691286
		), .Z(n_192791287));
	notech_ao4 i_131762094(.A(n_55966), .B(n_33758), .C(n_61085), .D(n_30776
		), .Z(n_192891288));
	notech_ao4 i_131662095(.A(n_55946), .B(n_31508), .C(n_55955), .D(n_30967
		), .Z(n_193091290));
	notech_ao4 i_3058091(.A(n_61718), .B(n_317460802), .C(n_193691296), .D(n_2039
		), .Z(n_193491294));
	notech_ao4 i_3158090(.A(n_19612), .B(n_72012477), .C(n_193891298), .D(n_26133
		), .Z(n_193691296));
	notech_ao4 i_3258089(.A(n_30304), .B(n_316160789), .C(n_349371378), .D(n_194091300
		), .Z(n_193891298));
	notech_and2 i_3358088(.A(n_347671363), .B(n_30681), .Z(n_194091300));
	notech_mux2 i_24258161(.S(n_61642), .A(n_19595), .B(n_195191311), .Z(n_194891308
		));
	notech_and2 i_75457409(.A(n_349171376), .B(n_59516), .Z(n_195191311));
	notech_ao3 i_8558036(.A(Daddrs_8[1]), .B(n_61642), .C(n_58848), .Z(n_195491314
		));
	notech_nor2 i_8258039(.A(n_56246), .B(n_32060), .Z(n_195791317));
	notech_ao3 i_7958042(.A(Daddrs_3[1]), .B(n_58628), .C(n_56226), .Z(n_196091320
		));
	notech_nand3 i_7458047(.A(n_210633637), .B(opd[1]), .C(n_61642), .Z(n_196191321
		));
	notech_or4 i_7558046(.A(n_61718), .B(n_61878), .C(n_56794), .D(n_59005),
		 .Z(n_196291322));
	notech_nand2 i_7658045(.A(Daddrs_1[1]), .B(n_56188), .Z(n_196391323));
	notech_nand3 i_49657657(.A(n_30367), .B(n_61643), .C(ecx[0]), .Z(n_196891328
		));
	notech_nand3 i_50157652(.A(n_30367), .B(n_61643), .C(ecx[1]), .Z(n_197391333
		));
	notech_nand3 i_50657647(.A(n_30367), .B(n_61643), .C(ecx[2]), .Z(n_197891338
		));
	notech_nand3 i_51157642(.A(n_30367), .B(n_61642), .C(ecx[3]), .Z(n_198391343
		));
	notech_nand3 i_51657637(.A(n_30367), .B(n_61642), .C(ecx[4]), .Z(n_198891348
		));
	notech_nand3 i_52157632(.A(n_30367), .B(n_61642), .C(ecx[5]), .Z(n_199391353
		));
	notech_nand3 i_52657627(.A(n_30367), .B(n_61642), .C(ecx[6]), .Z(n_199891358
		));
	notech_nand3 i_53157622(.A(n_30367), .B(n_61642), .C(ecx[7]), .Z(n_200391363
		));
	notech_nand3 i_53657617(.A(n_30367), .B(n_61642), .C(ecx[8]), .Z(n_200891368
		));
	notech_nand3 i_54257612(.A(n_30367), .B(n_61642), .C(ecx[9]), .Z(n_201391373
		));
	notech_nand3 i_54757607(.A(n_30367), .B(n_61642), .C(ecx[10]), .Z(n_201991378
		));
	notech_nand3 i_55257602(.A(n_61642), .B(n_30367), .C(ecx[11]), .Z(n_202491383
		));
	notech_nand3 i_55957597(.A(n_61642), .B(n_30367), .C(ecx[12]), .Z(n_202991388
		));
	notech_nand3 i_56457592(.A(n_61642), .B(n_30367), .C(ecx[13]), .Z(n_203491393
		));
	notech_nand3 i_56957587(.A(n_61643), .B(n_30367), .C(ecx[14]), .Z(n_203991398
		));
	notech_nand3 i_57457582(.A(n_61643), .B(n_58839), .C(ecx[15]), .Z(n_204491403
		));
	notech_nand3 i_57957577(.A(n_58839), .B(n_61643), .C(ecx[16]), .Z(n_204991408
		));
	notech_nand3 i_58457572(.A(n_58839), .B(n_61643), .C(ecx[17]), .Z(n_205491413
		));
	notech_nand3 i_58957567(.A(n_58839), .B(n_61643), .C(ecx[18]), .Z(n_205991418
		));
	notech_nand3 i_59457562(.A(n_58839), .B(n_61647), .C(ecx[19]), .Z(n_206491423
		));
	notech_and3 i_59957557(.A(n_58839), .B(n_61647), .C(ecx[20]), .Z(n_206991428
		));
	notech_nand3 i_60457552(.A(n_58839), .B(n_61643), .C(ecx[21]), .Z(n_207491433
		));
	notech_and3 i_60957547(.A(n_58839), .B(n_61643), .C(ecx[22]), .Z(n_207991438
		));
	notech_nand3 i_61457542(.A(n_58839), .B(n_61643), .C(ecx[23]), .Z(n_208491443
		));
	notech_and3 i_61957537(.A(n_58839), .B(n_61642), .C(ecx[24]), .Z(n_208991448
		));
	notech_and3 i_62457532(.A(n_58839), .B(n_61643), .C(ecx[25]), .Z(n_209591453
		));
	notech_nand3 i_62957527(.A(n_58839), .B(n_61642), .C(ecx[26]), .Z(n_210091458
		));
	notech_nand3 i_63557522(.A(n_58839), .B(n_61642), .C(ecx[27]), .Z(n_210591463
		));
	notech_nand3 i_64157517(.A(n_58839), .B(n_61642), .C(ecx[28]), .Z(n_211091468
		));
	notech_nand3 i_64757512(.A(n_58839), .B(n_61643), .C(ecx[29]), .Z(n_211591473
		));
	notech_nand3 i_65357507(.A(n_58839), .B(n_61643), .C(ecx[30]), .Z(n_212091478
		));
	notech_nand3 i_65857502(.A(n_58839), .B(n_61643), .C(ecx[31]), .Z(n_212591483
		));
	notech_or4 i_124356943(.A(n_61076), .B(n_32627), .C(n_60170), .D(n_61618
		), .Z(n_212691484));
	notech_ao4 i_80558126(.A(n_27924), .B(n_25705), .C(n_212691484), .D(n_210833639
		), .Z(n_213091485));
	notech_ao4 i_124156945(.A(n_4461), .B(n_60591), .C(n_4460), .D(n_58983),
		 .Z(n_213191486));
	notech_ao4 i_124056946(.A(n_61643), .B(n_32699), .C(n_390164432), .D(n_31834
		), .Z(n_213391488));
	notech_ao4 i_123856948(.A(n_4461), .B(n_60611), .C(n_4460), .D(n_58992),
		 .Z(n_213491489));
	notech_ao4 i_123756949(.A(n_61643), .B(n_32698), .C(n_390164432), .D(n_31833
		), .Z(n_213691491));
	notech_ao4 i_123556951(.A(n_4461), .B(nbus_11271[29]), .C(n_4460), .D(n_58947
		), .Z(n_213791492));
	notech_ao4 i_123456952(.A(n_61669), .B(n_32696), .C(n_390164432), .D(n_31832
		), .Z(n_213991494));
	notech_ao4 i_123256954(.A(n_4461), .B(n_60564), .C(n_4460), .D(n_58929),
		 .Z(n_214191495));
	notech_ao4 i_123156955(.A(n_61669), .B(n_32695), .C(n_390164432), .D(n_31831
		), .Z(n_214391497));
	notech_ao4 i_122956957(.A(n_4461), .B(nbus_11271[27]), .C(n_4460), .D(n_58938
		), .Z(n_214491498));
	notech_ao4 i_122856958(.A(n_61669), .B(n_32694), .C(n_390164432), .D(n_31830
		), .Z(n_214691500));
	notech_ao4 i_122556960(.A(n_4461), .B(nbus_11271[26]), .C(n_4460), .D(n_58911
		), .Z(n_214791501));
	notech_ao4 i_122256961(.A(n_61665), .B(n_32693), .C(n_390164432), .D(n_31829
		), .Z(n_214991503));
	notech_ao4 i_122056963(.A(n_4461), .B(n_60510), .C(n_4460), .D(n_58920),
		 .Z(n_215091504));
	notech_ao4 i_121956964(.A(n_61665), .B(n_32692), .C(n_390164432), .D(n_31828
		), .Z(n_215291506));
	notech_ao4 i_121756966(.A(n_4461), .B(n_60519), .C(n_4460), .D(n_58893),
		 .Z(n_215391507));
	notech_ao4 i_121656967(.A(n_61669), .B(n_32691), .C(n_390164432), .D(n_31827
		), .Z(n_215591509));
	notech_ao4 i_121356969(.A(n_4461), .B(nbus_11271[23]), .C(n_4460), .D(n_58902
		), .Z(n_215691510));
	notech_ao4 i_121256970(.A(n_61669), .B(n_32690), .C(n_390164432), .D(n_31826
		), .Z(n_215891512));
	notech_ao4 i_121056972(.A(n_4461), .B(n_60537), .C(n_4460), .D(n_58875),
		 .Z(n_215991513));
	notech_ao4 i_120956973(.A(n_61669), .B(n_32688), .C(n_390164432), .D(n_31825
		), .Z(n_216191515));
	notech_ao4 i_120756975(.A(n_4461), .B(n_60546), .C(n_4460), .D(n_58884),
		 .Z(n_216291516));
	notech_ao4 i_120656976(.A(n_61669), .B(n_32687), .C(n_390164432), .D(n_31824
		), .Z(n_216491518));
	notech_ao4 i_120456978(.A(n_4461), .B(n_60555), .C(n_4460), .D(n_58857),
		 .Z(n_216591519));
	notech_ao4 i_120356979(.A(n_61669), .B(n_32686), .C(n_390164432), .D(n_31823
		), .Z(n_216791521));
	notech_ao4 i_120156981(.A(n_4461), .B(n_60483), .C(n_4460), .D(n_58866),
		 .Z(n_216891522));
	notech_ao4 i_120056982(.A(n_61665), .B(n_32685), .C(n_390164432), .D(n_31822
		), .Z(n_217091524));
	notech_ao4 i_119856984(.A(n_4461), .B(n_60492), .C(n_4460), .D(n_59077),
		 .Z(n_217191525));
	notech_ao4 i_119756985(.A(n_61665), .B(n_32683), .C(n_390164432), .D(n_31821
		), .Z(n_217391527));
	notech_ao4 i_119556987(.A(n_4461), .B(n_60501), .C(n_4460), .D(n_59086),
		 .Z(n_217491528));
	notech_ao4 i_119456988(.A(n_61665), .B(n_32682), .C(n_390164432), .D(n_31820
		), .Z(n_217691530));
	notech_ao4 i_119256990(.A(n_4461), .B(n_60474), .C(n_4460), .D(n_59059),
		 .Z(n_217791531));
	notech_ao4 i_118856991(.A(n_61665), .B(n_32681), .C(n_58673), .D(n_31819
		), .Z(n_217991533));
	notech_ao4 i_118656993(.A(n_58637), .B(nbus_11271[15]), .C(n_58655), .D(n_59068
		), .Z(n_218091534));
	notech_ao4 i_118556994(.A(n_61665), .B(n_32680), .C(n_58673), .D(n_31818
		), .Z(n_218291536));
	notech_ao4 i_118356996(.A(n_58637), .B(nbus_11271[14]), .C(n_58655), .D(n_59041
		), .Z(n_218391537));
	notech_ao4 i_118256997(.A(n_61665), .B(n_32679), .C(n_58673), .D(n_31817
		), .Z(n_218591539));
	notech_ao4 i_118056999(.A(n_58637), .B(nbus_11271[13]), .C(n_58655), .D(n_58965
		), .Z(n_218691540));
	notech_ao4 i_117957000(.A(n_61665), .B(n_32678), .C(n_58673), .D(n_31816
		), .Z(n_218891542));
	notech_ao4 i_117757002(.A(n_58637), .B(nbus_11271[12]), .C(n_58655), .D(n_59050
		), .Z(n_218991543));
	notech_ao4 i_117657003(.A(n_61665), .B(n_32677), .C(n_58673), .D(n_31815
		), .Z(n_219191545));
	notech_ao4 i_117457005(.A(n_58637), .B(nbus_11271[11]), .C(n_58655), .D(n_58974
		), .Z(n_219291546));
	notech_ao4 i_117357006(.A(n_61665), .B(n_32676), .C(n_58673), .D(n_31814
		), .Z(n_219491548));
	notech_ao4 i_117157008(.A(n_58637), .B(nbus_11271[10]), .C(n_58655), .D(n_59023
		), .Z(n_219591549));
	notech_ao4 i_117057009(.A(n_61665), .B(n_32675), .C(n_58673), .D(n_31813
		), .Z(n_219791551));
	notech_ao4 i_116857011(.A(n_58637), .B(nbus_11271[9]), .C(n_58655), .D(n_59032
		), .Z(n_219891552));
	notech_ao4 i_116757012(.A(n_61669), .B(n_32674), .C(n_58673), .D(n_31812
		), .Z(n_220091554));
	notech_ao4 i_116557014(.A(n_58637), .B(nbus_11271[8]), .C(n_58655), .D(n_59014
		), .Z(n_220191555));
	notech_ao4 i_116457015(.A(n_61670), .B(n_32673), .C(n_58673), .D(n_31811
		), .Z(n_220391557));
	notech_ao4 i_116257017(.A(n_58637), .B(nbus_11271[7]), .C(n_58655), .D(\nbus_11290[7] 
		), .Z(n_220491558));
	notech_ao4 i_116157018(.A(n_61670), .B(n_32672), .C(n_58673), .D(n_31810
		), .Z(n_220691560));
	notech_ao4 i_115957020(.A(n_58637), .B(nbus_11271[6]), .C(n_58655), .D(\nbus_11290[6] 
		), .Z(n_220791561));
	notech_ao4 i_115857021(.A(n_61670), .B(n_32671), .C(n_58673), .D(n_31809
		), .Z(n_220991563));
	notech_ao4 i_115657023(.A(n_4461), .B(nbus_11271[5]), .C(n_4460), .D(\nbus_11290[5] 
		), .Z(n_221091564));
	notech_ao4 i_115557024(.A(n_61670), .B(n_32670), .C(n_390164432), .D(n_31808
		), .Z(n_221291566));
	notech_ao4 i_115357026(.A(n_58637), .B(nbus_11271[4]), .C(n_58655), .D(\nbus_11290[4] 
		), .Z(n_221391567));
	notech_ao4 i_115257027(.A(n_61670), .B(n_32669), .C(n_58673), .D(n_31807
		), .Z(n_221591569));
	notech_ao4 i_115057029(.A(n_58637), .B(nbus_11271[3]), .C(n_58655), .D(\nbus_11290[3] 
		), .Z(n_221691570));
	notech_ao4 i_114957030(.A(n_61670), .B(n_32668), .C(n_31806), .D(n_58673
		), .Z(n_221891572));
	notech_ao4 i_114757032(.A(n_58637), .B(nbus_11271[2]), .C(n_58655), .D(\nbus_11290[2] 
		), .Z(n_221991573));
	notech_ao4 i_114657033(.A(n_61675), .B(n_32667), .C(n_58673), .D(n_31805
		), .Z(n_222191575));
	notech_ao4 i_114457035(.A(n_58637), .B(nbus_11271[1]), .C(n_58655), .D(n_59005
		), .Z(n_222291576));
	notech_ao4 i_114357036(.A(n_61670), .B(n_32666), .C(n_58673), .D(n_31804
		), .Z(n_222491578));
	notech_ao4 i_114157038(.A(n_58637), .B(nbus_11271[0]), .C(n_58655), .D(\nbus_11290[0] 
		), .Z(n_222591579));
	notech_ao4 i_114057039(.A(n_61670), .B(n_32665), .C(n_58673), .D(n_31803
		), .Z(n_222791581));
	notech_nand3 i_80357360(.A(n_196291322), .B(n_196191321), .C(n_196391323
		), .Z(n_223091584));
	notech_ao4 i_80057363(.A(n_56235), .B(n_33761), .C(n_56215), .D(n_33760)
		, .Z(n_223191585));
	notech_ao4 i_79757366(.A(n_56268), .B(n_31932), .C(n_56257), .D(nbus_11271
		[1]), .Z(n_223491588));
	notech_ao4 i_79557368(.A(n_58619), .B(n_31329), .C(n_58646), .D(n_33759)
		, .Z(n_223691590));
	notech_or4 i_79957364(.A(n_195491314), .B(n_195791317), .C(n_30686), .D(n_30685
		), .Z(n_223891592));
	notech_or4 i_79555986(.A(n_61076), .B(n_61739), .C(n_60170), .D(n_230891662
		), .Z(n_223991593));
	notech_nand3 i_10655820(.A(n_284331524), .B(n_194984376), .C(n_295392296
		), .Z(n_224091594));
	notech_ao4 i_9855828(.A(n_224991603), .B(n_30687), .C(CFOF_mul), .D(n_284331524
		), .Z(n_224391597));
	notech_mux2 i_9955827(.S(n_61670), .A(n_27823), .B(n_316760795), .Z(n_224491598
		));
	notech_or4 i_10055826(.A(n_230491658), .B(n_230591659), .C(n_230391657),
		 .D(n_30699), .Z(n_224591599));
	notech_and4 i_10155825(.A(n_232191675), .B(n_231991673), .C(n_230091654)
		, .D(n_229791651), .Z(n_224691600));
	notech_and4 i_10255824(.A(n_235491708), .B(n_234791701), .C(n_233991693)
		, .D(n_233291686), .Z(n_224791601));
	notech_ao4 i_8455842(.A(n_30696), .B(n_32702), .C(n_27922), .D(n_96629667
		), .Z(n_224991603));
	notech_or4 i_98454999(.A(n_32574), .B(n_309960727), .C(n_61076), .D(n_61052
		), .Z(n_225391607));
	notech_nand3 i_48155478(.A(n_58532), .B(n_224591599), .C(n_61669), .Z(n_225791611
		));
	notech_or4 i_48255477(.A(n_61718), .B(n_61878), .C(n_58532), .D(n_224691600
		), .Z(n_225891612));
	notech_and3 i_47755482(.A(n_30687), .B(n_27826), .C(n_27827), .Z(n_226191615
		));
	notech_and4 i_47855481(.A(n_1839), .B(rep_en2), .C(nCF_shift4box), .D(n_61618
		), .Z(n_226291616));
	notech_or4 i_50055459(.A(n_32396), .B(n_61739), .C(n_60170), .D(n_32768)
		, .Z(n_229791651));
	notech_nao3 i_49755462(.A(nbus_133[32]), .B(n_32697), .C(n_27924), .Z(n_230091654
		));
	notech_and3 i_49055469(.A(nbus_134[16]), .B(n_32321), .C(n_27923), .Z(n_230391657
		));
	notech_and4 i_49155468(.A(nbus_143[16]), .B(n_61953), .C(n_63762), .D(n_27933
		), .Z(n_230491658));
	notech_and4 i_49255467(.A(n_27933), .B(nbus_137[16]), .C(n_61953), .D(n_61933
		), .Z(n_230591659));
	notech_ao3 i_22785(.A(n_316260790), .B(n_224091594), .C(n_61878), .Z(n_230691660
		));
	notech_or4 i_185454143(.A(n_61878), .B(n_61718), .C(n_61866), .D(n_4450)
		, .Z(n_230891662));
	notech_ao4 i_132154669(.A(n_224491598), .B(n_33763), .C(n_224391597), .D
		(n_61618), .Z(n_231291666));
	notech_ao4 i_135854632(.A(n_58523), .B(n_32837), .C(n_27920), .D(n_32820
		), .Z(n_231891672));
	notech_ao4 i_135654634(.A(n_27922), .B(n_30369), .C(n_27930), .D(n_32913
		), .Z(n_231991673));
	notech_ao4 i_135454636(.A(n_27920), .B(n_32752), .C(n_27932), .D(n_32735
		), .Z(n_232191675));
	notech_or4 i_2355903(.A(n_312460752), .B(n_2952), .C(n_60170), .D(n_27909
		), .Z(n_232591679));
	notech_ao4 i_135054640(.A(n_58465), .B(n_32056), .C(n_32057), .D(n_58474
		), .Z(n_232691680));
	notech_ao4 i_134954641(.A(n_58447), .B(n_32054), .C(n_58456), .D(n_32055
		), .Z(n_232791681));
	notech_ao4 i_134754643(.A(n_58225), .B(n_32029), .C(n_32028), .D(n_58238
		), .Z(n_232991683));
	notech_ao4 i_134654644(.A(n_58247), .B(n_32030), .C(n_58256), .D(n_32031
		), .Z(n_233091684));
	notech_and4 i_135254638(.A(n_233091684), .B(n_232991683), .C(n_232791681
		), .D(n_232691680), .Z(n_233291686));
	notech_ao4 i_134354647(.A(nbus_11273[4]), .B(n_32032), .C(nbus_11273[5])
		, .D(n_32033), .Z(n_233391687));
	notech_ao4 i_134254648(.A(n_58265), .B(n_32034), .C(n_58275), .D(n_32035
		), .Z(n_233491688));
	notech_ao4 i_134054650(.A(n_32036), .B(n_58285), .C(n_58294), .D(n_32037
		), .Z(n_233691690));
	notech_ao4 i_133954651(.A(n_32038), .B(n_58303), .C(n_58312), .D(n_32039
		), .Z(n_233791691));
	notech_and4 i_134554645(.A(n_233791691), .B(n_233691690), .C(n_233491688
		), .D(n_233391687), .Z(n_233991693));
	notech_ao4 i_133554655(.A(n_58321), .B(n_32040), .C(n_58330), .D(n_32041
		), .Z(n_234191695));
	notech_ao4 i_133454656(.A(n_32042), .B(n_58339), .C(n_32043), .D(n_58348
		), .Z(n_234291696));
	notech_ao4 i_133254658(.A(n_32044), .B(n_58357), .C(n_32045), .D(n_58366
		), .Z(n_234491698));
	notech_ao4 i_133154659(.A(n_32046), .B(n_58375), .C(n_32047), .D(n_58384
		), .Z(n_234591699));
	notech_and4 i_133754653(.A(n_234591699), .B(n_234491698), .C(n_234291696
		), .D(n_234191695), .Z(n_234791701));
	notech_ao4 i_132854662(.A(n_32048), .B(n_58393), .C(n_32049), .D(n_58402
		), .Z(n_234891702));
	notech_ao4 i_132754663(.A(n_32050), .B(n_58411), .C(n_32051), .D(n_58420
		), .Z(n_234991703));
	notech_ao4 i_132554665(.A(n_58429), .B(n_32052), .C(n_58438), .D(n_32053
		), .Z(n_235191705));
	notech_ao4 i_132454666(.A(n_32058), .B(n_58483), .C(n_60458), .D(n_32059
		), .Z(n_235291706));
	notech_and4 i_133054660(.A(n_235291706), .B(n_235191705), .C(n_234991703
		), .D(n_234891702), .Z(n_235491708));
	notech_ao4 i_131854672(.A(n_58215), .B(n_33762), .C(n_224791601), .D(n_232591679
		), .Z(n_235691710));
	notech_nand3 i_132054670(.A(n_225891612), .B(n_235691710), .C(n_225791611
		), .Z(n_235791711));
	notech_xor2 i_4753027(.A(vliw_pc[1]), .B(vliw_pc[0]), .Z(n_235891712));
	notech_xor2 i_4853026(.A(vliw_pc[2]), .B(n_32779), .Z(n_235991713));
	notech_xor2 i_4953025(.A(n_31257), .B(n_310892436), .Z(n_236091714));
	notech_ao4 i_5053024(.A(n_236491718), .B(n_31258), .C(n_32756), .D(n_310892436
		), .Z(n_236191715));
	notech_and4 i_1953051(.A(vliw_pc[1]), .B(vliw_pc[0]), .C(vliw_pc[2]), .D
		(vliw_pc[3]), .Z(n_236491718));
	notech_and2 i_2746385(.A(n_23847), .B(n_30701), .Z(n_236991723));
	notech_ao4 i_2846384(.A(n_32627), .B(n_29534), .C(n_4086), .D(n_25670), 
		.Z(n_237091724));
	notech_xor2 i_2546387(.A(opc[0]), .B(opc[1]), .Z(n_237191725));
	notech_ao3 i_2646386(.A(n_56929), .B(n_240891762), .C(n_4442), .Z(n_237291726
		));
	notech_and2 i_2346389(.A(n_4444), .B(n_237591729), .Z(n_237391727));
	notech_and2 i_2446388(.A(n_237691730), .B(n_4453), .Z(n_237491728));
	notech_nao3 i_10046312(.A(opc[0]), .B(opc[1]), .C(n_23847), .Z(n_237591729
		));
	notech_or2 i_10146311(.A(n_23847), .B(n_57222), .Z(n_237691730));
	notech_and3 i_2146390(.A(n_4028), .B(n_4453), .C(n_237891732), .Z(n_237791731
		));
	notech_nand2 i_11946295(.A(n_4445), .B(opc[2]), .Z(n_237891732));
	notech_nao3 i_8446328(.A(n_406282377), .B(n_3683), .C(n_57336), .Z(n_239391747
		));
	notech_or2 i_8546327(.A(n_23847), .B(n_60467), .Z(n_240891762));
	notech_nao3 i_11846296(.A(nbus_11271[3]), .B(nbus_11271[2]), .C(n_4444),
		 .Z(n_242391777));
	notech_or4 i_12946285(.A(n_61065), .B(n_58610), .C(n_61616), .D(nbus_11271
		[24]), .Z(n_244291796));
	notech_nao3 i_12646288(.A(n_30371), .B(n_3657), .C(n_24147), .Z(n_244591799
		));
	notech_or4 i_14146273(.A(n_61065), .B(n_58610), .C(n_61616), .D(nbus_11271
		[25]), .Z(n_245591808));
	notech_nao3 i_13846276(.A(n_30371), .B(n_3658), .C(n_24147), .Z(n_245891811
		));
	notech_or4 i_15346261(.A(n_61065), .B(n_58610), .C(n_61616), .D(n_60582)
		, .Z(n_247091820));
	notech_nao3 i_15046264(.A(n_30371), .B(n_3659), .C(n_24147), .Z(n_247391823
		));
	notech_or4 i_16546249(.A(n_61065), .B(n_58610), .C(n_61618), .D(n_60573)
		, .Z(n_248291832));
	notech_nao3 i_16246252(.A(n_30371), .B(n_3660), .C(n_24147), .Z(n_248591835
		));
	notech_or4 i_17746237(.A(n_61065), .B(n_58610), .C(n_61616), .D(n_60564)
		, .Z(n_249491844));
	notech_nao3 i_17446240(.A(n_30371), .B(n_3661), .C(n_24147), .Z(n_249791847
		));
	notech_or4 i_18946225(.A(n_61065), .B(n_340561033), .C(n_61616), .D(n_60620
		), .Z(n_250691856));
	notech_nao3 i_18646228(.A(n_30371), .B(n_3662), .C(n_24147), .Z(n_250991859
		));
	notech_or4 i_20146213(.A(n_61065), .B(n_58610), .C(n_61618), .D(nbus_11271
		[30]), .Z(n_251891868));
	notech_nao3 i_19846216(.A(n_30371), .B(n_3663), .C(n_24147), .Z(n_252191871
		));
	notech_nand2 i_21246202(.A(n_30422), .B(opb[16]), .Z(n_252691876));
	notech_or2 i_21146203(.A(n_24144), .B(nbus_11270[16]), .Z(n_252991879)
		);
	notech_nao3 i_20646208(.A(\opc_5[16] ), .B(n_30364), .C(n_4086), .Z(n_253491884
		));
	notech_nand2 i_22146193(.A(n_30422), .B(opb[17]), .Z(n_253591885));
	notech_or2 i_22046194(.A(n_24141), .B(nbus_11271[9]), .Z(n_253891888));
	notech_nand2 i_21546199(.A(opc_14[17]), .B(n_19698), .Z(n_254391893));
	notech_nand2 i_23046184(.A(n_30422), .B(opb[18]), .Z(n_254491894));
	notech_or2 i_22946185(.A(n_24141), .B(nbus_11271[10]), .Z(n_254791897)
		);
	notech_nand2 i_22446190(.A(opc_14[18]), .B(n_19698), .Z(n_255291902));
	notech_nand2 i_23946175(.A(n_30422), .B(opb[19]), .Z(n_255391903));
	notech_or2 i_23846176(.A(n_24141), .B(nbus_11271[11]), .Z(n_255691906)
		);
	notech_nand2 i_23346181(.A(opc_14[19]), .B(n_19698), .Z(n_256191911));
	notech_nand2 i_24946166(.A(n_30422), .B(opb[20]), .Z(n_256291912));
	notech_or2 i_24746167(.A(n_24141), .B(nbus_11271[12]), .Z(n_256591915)
		);
	notech_nand2 i_24246172(.A(opc_14[20]), .B(n_19698), .Z(n_257091920));
	notech_nand2 i_25946157(.A(n_30422), .B(opb[21]), .Z(n_257191921));
	notech_or2 i_25746158(.A(n_24141), .B(nbus_11271[13]), .Z(n_257491924)
		);
	notech_nand2 i_25246163(.A(opc_14[21]), .B(n_61119), .Z(n_257991929));
	notech_nand2 i_26946148(.A(n_30422), .B(opb[22]), .Z(n_258091930));
	notech_or2 i_26746149(.A(n_24141), .B(nbus_11271[14]), .Z(n_258391933)
		);
	notech_nand2 i_26246154(.A(opc_14[22]), .B(n_61119), .Z(n_258891938));
	notech_nand2 i_27946139(.A(n_30422), .B(opb[23]), .Z(n_258991939));
	notech_or2 i_27746140(.A(n_24141), .B(nbus_11271[15]), .Z(n_259291942)
		);
	notech_nand2 i_27246145(.A(opc_14[23]), .B(n_61119), .Z(n_259791947));
	notech_nand2 i_28846130(.A(n_30422), .B(opb[24]), .Z(n_259891948));
	notech_or2 i_28746131(.A(n_24141), .B(nbus_11271[0]), .Z(n_260191951));
	notech_nand2 i_28246136(.A(opc_14[24]), .B(n_61119), .Z(n_260691956));
	notech_nand2 i_29746121(.A(n_30422), .B(opb[25]), .Z(n_260791957));
	notech_or2 i_29646122(.A(n_24141), .B(nbus_11271[1]), .Z(n_261091960));
	notech_nand2 i_29146127(.A(opc_14[25]), .B(n_61119), .Z(n_261591965));
	notech_nand2 i_30646112(.A(n_30422), .B(opb[26]), .Z(n_261691966));
	notech_or2 i_30546113(.A(n_24141), .B(nbus_11271[2]), .Z(n_261991969));
	notech_nand2 i_30046118(.A(opc_14[26]), .B(n_61119), .Z(n_262491974));
	notech_nand2 i_31546103(.A(n_30422), .B(opb[27]), .Z(n_262591975));
	notech_or2 i_31446104(.A(n_24141), .B(nbus_11271[3]), .Z(n_262891978));
	notech_nand2 i_30946109(.A(opc_14[27]), .B(n_61119), .Z(n_263391983));
	notech_nand2 i_32446094(.A(n_30422), .B(opb[29]), .Z(n_263491984));
	notech_or2 i_32346095(.A(n_24141), .B(nbus_11271[5]), .Z(n_263791987));
	notech_nand2 i_31846100(.A(opc_14[29]), .B(n_19698), .Z(n_264291992));
	notech_nand2 i_33346085(.A(n_30422), .B(opb[30]), .Z(n_264391993));
	notech_or2 i_33246086(.A(n_24141), .B(nbus_11271[6]), .Z(n_264691996));
	notech_nand2 i_32746091(.A(opc_14[30]), .B(n_61119), .Z(n_265192001));
	notech_or2 i_34246076(.A(n_24141), .B(nbus_11271[7]), .Z(n_265292002));
	notech_nand3 i_34146077(.A(divr[31]), .B(n_30371), .C(n_24147), .Z(n_265592005
		));
	notech_or2 i_33646082(.A(n_4447), .B(n_31642), .Z(n_266092010));
	notech_ao4 i_139645100(.A(n_56929), .B(n_60591), .C(n_4446), .D(n_58983)
		, .Z(n_266192011));
	notech_ao4 i_139545101(.A(n_30712), .B(n_32931), .C(n_24134), .D(n_33810
		), .Z(n_266392013));
	notech_ao4 i_139245104(.A(n_24138), .B(n_33809), .C(n_218373551), .D(n_33689
		), .Z(n_266592015));
	notech_and4 i_139445102(.A(n_24127), .B(n_266592015), .C(n_265292002), .D
		(n_265592005), .Z(n_266892018));
	notech_ao4 i_138645108(.A(n_24134), .B(n_33808), .C(n_4447), .D(n_31641)
		, .Z(n_266992019));
	notech_ao4 i_138345109(.A(n_218373551), .B(n_33690), .C(n_56929), .D(n_60611
		), .Z(n_267192021));
	notech_ao4 i_138045112(.A(n_24144), .B(nbus_11270[30]), .C(n_24138), .D(n_33807
		), .Z(n_267392023));
	notech_and4 i_138245110(.A(n_24127), .B(n_267392023), .C(n_264391993), .D
		(n_264691996), .Z(n_267692026));
	notech_ao4 i_137645116(.A(n_24134), .B(n_33806), .C(n_4447), .D(n_31640)
		, .Z(n_267792027));
	notech_ao4 i_137545117(.A(n_218373551), .B(n_33691), .C(n_56929), .D(n_60620
		), .Z(n_267992029));
	notech_ao4 i_137245120(.A(n_24144), .B(nbus_11270[29]), .C(n_24138), .D(n_33805
		), .Z(n_268192031));
	notech_and4 i_137445118(.A(n_24127), .B(n_268192031), .C(n_263491984), .D
		(n_263791987), .Z(n_268492034));
	notech_ao4 i_136845124(.A(n_24134), .B(n_33804), .C(n_4447), .D(n_31638)
		, .Z(n_268592035));
	notech_ao4 i_136745125(.A(n_218373551), .B(n_33692), .C(n_56929), .D(n_60573
		), .Z(n_268792037));
	notech_ao4 i_136245128(.A(n_24144), .B(nbus_11270[27]), .C(n_24138), .D(n_33803
		), .Z(n_268992039));
	notech_and4 i_136645126(.A(n_24127), .B(n_268992039), .C(n_262591975), .D
		(n_262891978), .Z(n_269292042));
	notech_ao4 i_135745132(.A(n_24134), .B(n_33802), .C(n_4447), .D(n_31637)
		, .Z(n_269392043));
	notech_ao4 i_135645133(.A(n_218373551), .B(n_33693), .C(n_56929), .D(n_60582
		), .Z(n_269592045));
	notech_ao4 i_135345136(.A(n_24144), .B(nbus_11270[26]), .C(n_24138), .D(n_33801
		), .Z(n_269792047));
	notech_and4 i_135545134(.A(n_24127), .B(n_269792047), .C(n_261691966), .D
		(n_261991969), .Z(n_270092050));
	notech_ao4 i_134945140(.A(n_24134), .B(n_33800), .C(n_4447), .D(n_31636)
		, .Z(n_270192051));
	notech_ao4 i_134845141(.A(n_57978), .B(n_33694), .C(n_56929), .D(n_60510
		), .Z(n_270392053));
	notech_ao4 i_134545144(.A(n_24144), .B(nbus_11270[25]), .C(n_24138), .D(n_33799
		), .Z(n_270692055));
	notech_and4 i_134745142(.A(n_24127), .B(n_270692055), .C(n_260791957), .D
		(n_261091960), .Z(n_271092058));
	notech_ao4 i_134145148(.A(n_24134), .B(n_33798), .C(n_4447), .D(n_31635)
		, .Z(n_271192059));
	notech_ao4 i_134045149(.A(n_57974), .B(n_33695), .C(n_56929), .D(n_60519
		), .Z(n_271392061));
	notech_ao4 i_133745152(.A(n_24144), .B(nbus_11270[24]), .C(n_24138), .D(n_33797
		), .Z(n_271592063));
	notech_and4 i_133945150(.A(n_24127), .B(n_271592063), .C(n_259891948), .D
		(n_260191951), .Z(n_271892066));
	notech_ao4 i_133345156(.A(n_24134), .B(n_33796), .C(n_4447), .D(n_31634)
		, .Z(n_271992067));
	notech_ao4 i_133245157(.A(n_57974), .B(n_33696), .C(n_56923), .D(n_60528
		), .Z(n_272192069));
	notech_ao4 i_132945160(.A(n_24144), .B(nbus_11270[23]), .C(n_24138), .D(n_33795
		), .Z(n_272392071));
	notech_and4 i_133145158(.A(n_24127), .B(n_272392071), .C(n_258991939), .D
		(n_259291942), .Z(n_272692074));
	notech_ao4 i_132545164(.A(n_24134), .B(n_33794), .C(n_4447), .D(n_31633)
		, .Z(n_272792075));
	notech_ao4 i_132445165(.A(n_57974), .B(n_33697), .C(n_56923), .D(n_60537
		), .Z(n_272992077));
	notech_ao4 i_132145168(.A(n_24144), .B(nbus_11270[22]), .C(n_24138), .D(n_33793
		), .Z(n_273192079));
	notech_and4 i_132345166(.A(n_24127), .B(n_273192079), .C(n_258091930), .D
		(n_258391933), .Z(n_273492082));
	notech_ao4 i_131745172(.A(n_24134), .B(n_33792), .C(n_4447), .D(n_31632)
		, .Z(n_273592083));
	notech_ao4 i_131645173(.A(n_57978), .B(n_33698), .C(n_56923), .D(n_60546
		), .Z(n_273792085));
	notech_ao4 i_131345176(.A(n_24144), .B(nbus_11270[21]), .C(n_24138), .D(n_33791
		), .Z(n_273992087));
	notech_and4 i_131545174(.A(n_24127), .B(n_273992087), .C(n_257191921), .D
		(n_257491924), .Z(n_274292090));
	notech_ao4 i_130945180(.A(n_24134), .B(n_33790), .C(n_4447), .D(n_31631)
		, .Z(n_274392091));
	notech_ao4 i_130845181(.A(n_57974), .B(n_33699), .C(n_56923), .D(n_60555
		), .Z(n_274592093));
	notech_ao4 i_130545184(.A(n_24144), .B(nbus_11270[20]), .C(n_24138), .D(n_33789
		), .Z(n_274792095));
	notech_and4 i_130745182(.A(n_24127), .B(n_274792095), .C(n_256291912), .D
		(n_256591915), .Z(n_275092098));
	notech_ao4 i_130045188(.A(n_24134), .B(n_33788), .C(n_4447), .D(n_31630)
		, .Z(n_275192099));
	notech_ao4 i_129945189(.A(n_57974), .B(n_33700), .C(n_56923), .D(n_60483
		), .Z(n_275392101));
	notech_ao4 i_129645192(.A(n_24144), .B(nbus_11270[19]), .C(n_56728), .D(n_33787
		), .Z(n_275792103));
	notech_and4 i_129845190(.A(n_24127), .B(n_275792103), .C(n_255391903), .D
		(n_255691906), .Z(n_276092106));
	notech_ao4 i_129145196(.A(n_56774), .B(n_33786), .C(n_4447), .D(n_31629)
		, .Z(n_276192107));
	notech_ao4 i_129045197(.A(n_57974), .B(n_33701), .C(n_56923), .D(n_60492
		), .Z(n_276392109));
	notech_ao4 i_128745200(.A(n_24144), .B(nbus_11270[18]), .C(n_56728), .D(n_33785
		), .Z(n_276592111));
	notech_and4 i_128945198(.A(n_24127), .B(n_276592111), .C(n_254491894), .D
		(n_254791897), .Z(n_276892114));
	notech_ao4 i_128345204(.A(n_56774), .B(n_33784), .C(n_4447), .D(n_31628)
		, .Z(n_276992115));
	notech_ao4 i_128245205(.A(n_57974), .B(n_33702), .C(n_56923), .D(n_60501
		), .Z(n_277192117));
	notech_ao4 i_127945208(.A(n_24144), .B(nbus_11270[17]), .C(n_56728), .D(n_33783
		), .Z(n_277392119));
	notech_and4 i_128145206(.A(n_24127), .B(n_277392119), .C(n_253591885), .D
		(n_253891888), .Z(n_277692122));
	notech_ao4 i_127345212(.A(n_4447), .B(n_31627), .C(n_24141), .D(nbus_11271
		[8]), .Z(n_277792123));
	notech_ao4 i_127245213(.A(n_56923), .B(n_60474), .C(n_30712), .D(n_32930
		), .Z(n_277992125));
	notech_ao4 i_126745216(.A(n_56728), .B(n_33782), .C(n_57974), .D(n_33703
		), .Z(n_278192127));
	notech_and4 i_127145214(.A(n_24127), .B(n_278192127), .C(n_252691876), .D
		(n_252991879), .Z(n_278492130));
	notech_ao4 i_125945220(.A(n_56762), .B(n_31625), .C(n_4446), .D(n_59041)
		, .Z(n_278592131));
	notech_ao4 i_125845221(.A(n_30712), .B(n_32928), .C(n_56774), .D(n_33781
		), .Z(n_278692132));
	notech_ao4 i_125645223(.A(n_57974), .B(n_33704), .C(n_56923), .D(\nbus_11290[6] 
		), .Z(n_278892134));
	notech_and4 i_126145218(.A(n_278892134), .B(n_278692132), .C(n_278592131
		), .D(n_252191871), .Z(n_279092136));
	notech_ao4 i_125345226(.A(n_56707), .B(n_60537), .C(n_24144), .D(nbus_11270
		[14]), .Z(n_279192137));
	notech_ao4 i_125145228(.A(n_23989), .B(n_33412), .C(n_23988), .D(n_31538
		), .Z(n_279392139));
	notech_and4 i_125545224(.A(n_56750), .B(n_279392139), .C(n_279192137), .D
		(n_251891868), .Z(n_279592141));
	notech_ao4 i_124845231(.A(n_56762), .B(n_31624), .C(n_58965), .D(n_4446)
		, .Z(n_279692142));
	notech_ao4 i_124745232(.A(n_30712), .B(n_32927), .C(n_56774), .D(n_33780
		), .Z(n_279792143));
	notech_ao4 i_124545234(.A(n_57974), .B(n_33705), .C(n_56923), .D(\nbus_11290[5] 
		), .Z(n_279992145));
	notech_and4 i_125045229(.A(n_279992145), .B(n_279792143), .C(n_279692142
		), .D(n_250991859), .Z(n_280192147));
	notech_ao4 i_124045237(.A(n_56707), .B(n_60546), .C(n_56738), .D(nbus_11270
		[13]), .Z(n_280292148));
	notech_ao4 i_123645239(.A(n_23989), .B(n_33410), .C(n_23988), .D(n_31537
		), .Z(n_280492150));
	notech_and4 i_124245235(.A(n_56750), .B(n_280492150), .C(n_280292148), .D
		(n_250691856), .Z(n_280692152));
	notech_ao4 i_123345242(.A(n_56762), .B(n_31623), .C(n_4446), .D(n_59050)
		, .Z(n_280792153));
	notech_ao4 i_123245243(.A(n_30712), .B(n_32926), .C(n_56774), .D(n_33779
		), .Z(n_280892154));
	notech_ao4 i_123045245(.A(n_57978), .B(n_33706), .C(n_56923), .D(\nbus_11290[4] 
		), .Z(n_281092156));
	notech_and4 i_123545240(.A(n_281092156), .B(n_280892154), .C(n_280792153
		), .D(n_249791847), .Z(n_281292158));
	notech_ao4 i_122745248(.A(n_56707), .B(n_60555), .C(n_56738), .D(nbus_11270
		[12]), .Z(n_281392159));
	notech_ao4 i_122545250(.A(n_23989), .B(n_33408), .C(n_23988), .D(n_31536
		), .Z(n_281592161));
	notech_and4 i_122945246(.A(n_56750), .B(n_281592161), .C(n_281392159), .D
		(n_249491844), .Z(n_281792163));
	notech_ao4 i_122245253(.A(n_56762), .B(n_31622), .C(n_4446), .D(n_58974)
		, .Z(n_281892164));
	notech_ao4 i_122145254(.A(n_30712), .B(n_32925), .C(n_56774), .D(n_33778
		), .Z(n_281992165));
	notech_ao4 i_121945256(.A(n_57978), .B(n_33707), .C(n_56923), .D(\nbus_11290[3] 
		), .Z(n_282192167));
	notech_and4 i_122445251(.A(n_282192167), .B(n_281992165), .C(n_281892164
		), .D(n_248591835), .Z(n_282392169));
	notech_ao4 i_121645259(.A(n_56707), .B(n_60483), .C(n_56738), .D(nbus_11270
		[11]), .Z(n_282492170));
	notech_ao4 i_121445261(.A(n_23989), .B(n_33406), .C(n_23988), .D(n_31535
		), .Z(n_282692172));
	notech_and4 i_121845257(.A(n_56750), .B(n_282692172), .C(n_282492170), .D
		(n_248291832), .Z(n_282892174));
	notech_ao4 i_121145264(.A(n_56762), .B(n_31621), .C(n_4446), .D(n_59023)
		, .Z(n_282992175));
	notech_ao4 i_121045265(.A(n_30712), .B(n_32924), .C(n_56774), .D(n_33777
		), .Z(n_283092176));
	notech_ao4 i_120845267(.A(n_57978), .B(n_33708), .C(n_56929), .D(\nbus_11290[2] 
		), .Z(n_283292178));
	notech_and4 i_121345262(.A(n_283292178), .B(n_283092176), .C(n_282992175
		), .D(n_247391823), .Z(n_283492180));
	notech_ao4 i_120545270(.A(n_56707), .B(n_60492), .C(n_56738), .D(nbus_11270
		[10]), .Z(n_283592181));
	notech_ao4 i_120345272(.A(n_23989), .B(n_33404), .C(n_23988), .D(n_31534
		), .Z(n_283792183));
	notech_and4 i_120745268(.A(n_56750), .B(n_283792183), .C(n_283592181), .D
		(n_247091820), .Z(n_283992185));
	notech_ao4 i_120045275(.A(n_56923), .B(n_59005), .C(n_4446), .D(n_59032)
		, .Z(n_284092186));
	notech_ao4 i_119945276(.A(n_56774), .B(n_33776), .C(n_56762), .D(n_31620
		), .Z(n_284192187));
	notech_ao4 i_119745278(.A(n_57978), .B(n_33709), .C(n_61110), .D(n_32923
		), .Z(n_284392189));
	notech_and4 i_120245273(.A(n_284392189), .B(n_284192187), .C(n_284092186
		), .D(n_245891811), .Z(n_284592191));
	notech_ao4 i_119245281(.A(n_56707), .B(n_60501), .C(n_56738), .D(nbus_11270
		[9]), .Z(n_284692192));
	notech_ao4 i_119045283(.A(n_23989), .B(n_33402), .C(n_23988), .D(n_31533
		), .Z(n_284892194));
	notech_and4 i_119645279(.A(n_56750), .B(n_284892194), .C(n_284692192), .D
		(n_245591808), .Z(n_285092196));
	notech_ao4 i_118545286(.A(n_56923), .B(\nbus_11290[0] ), .C(n_4446), .D(n_59014
		), .Z(n_285192197));
	notech_ao4 i_118445287(.A(n_56774), .B(n_33775), .C(n_56762), .D(n_31619
		), .Z(n_285292198));
	notech_ao4 i_118245289(.A(n_57978), .B(n_33710), .C(n_61110), .D(n_32922
		), .Z(n_285492200));
	notech_and4 i_118945284(.A(n_285492200), .B(n_285292198), .C(n_285192197
		), .D(n_244591799), .Z(n_285692202));
	notech_ao4 i_117945292(.A(n_56707), .B(n_60474), .C(n_56738), .D(nbus_11270
		[8]), .Z(n_285792203));
	notech_ao4 i_117745294(.A(n_23989), .B(n_33400), .C(n_23988), .D(n_31532
		), .Z(n_285992205));
	notech_and4 i_118145290(.A(n_56750), .B(n_285992205), .C(n_285792203), .D
		(n_244291796), .Z(n_286192207));
	notech_ao4 i_117445297(.A(n_444982454), .B(n_317051260), .C(n_237791731)
		, .D(nbus_11271[3]), .Z(n_286292208));
	notech_ao4 i_117345298(.A(n_56762), .B(n_31614), .C(n_25433), .D(n_58974
		), .Z(n_286392209));
	notech_ao4 i_117145300(.A(n_57978), .B(n_33711), .C(n_61110), .D(n_32917
		), .Z(n_286592211));
	notech_ao4 i_117045301(.A(n_56738), .B(nbus_11270[3]), .C(n_56728), .D(n_33774
		), .Z(n_286692212));
	notech_and4 i_117645295(.A(n_286692212), .B(n_286592211), .C(n_286392209
		), .D(n_286292208), .Z(n_286892214));
	notech_ao4 i_116745304(.A(n_4446), .B(\nbus_11290[3] ), .C(n_56707), .D(n_60573
		), .Z(n_286992215));
	notech_ao4 i_116645305(.A(n_23989), .B(n_33390), .C(n_23988), .D(n_31527
		), .Z(n_287092216));
	notech_ao4 i_116445307(.A(n_23839), .B(n_33773), .C(n_23836), .D(n_33772
		), .Z(n_287292218));
	notech_and3 i_116545306(.A(n_56750), .B(n_287292218), .C(n_242391777), .Z
		(n_287592220));
	notech_mux2 i_116045311(.S(opc[2]), .A(n_237391727), .B(n_237491728), .Z
		(n_287792222));
	notech_ao4 i_115945312(.A(n_56762), .B(n_31613), .C(n_25433), .D(n_59023
		), .Z(n_287892223));
	notech_ao4 i_115745314(.A(n_57978), .B(n_33712), .C(n_61110), .D(n_32916
		), .Z(n_288092225));
	notech_ao4 i_115645315(.A(n_56738), .B(nbus_11270[2]), .C(n_56728), .D(n_33771
		), .Z(n_288192226));
	notech_and4 i_116245309(.A(n_288192226), .B(n_288092225), .C(n_287892223
		), .D(n_287792222), .Z(n_288392228));
	notech_ao4 i_115145318(.A(n_4446), .B(\nbus_11290[2] ), .C(n_56707), .D(n_60582
		), .Z(n_288492229));
	notech_ao4 i_114845319(.A(n_23989), .B(n_33388), .C(n_23988), .D(n_31526
		), .Z(n_288592230));
	notech_ao4 i_114645321(.A(n_23839), .B(n_33770), .C(n_23836), .D(n_33769
		), .Z(n_288792232));
	notech_and4 i_115545316(.A(n_56750), .B(n_288792232), .C(n_288592230), .D
		(n_288492229), .Z(n_288992234));
	notech_or2 i_114545322(.A(n_23847), .B(opc[1]), .Z(n_289092235));
	notech_ao4 i_113945326(.A(n_237191725), .B(n_30701), .C(n_289092235), .D
		(nbus_11271[0]), .Z(n_289192236));
	notech_ao4 i_113845327(.A(n_25433), .B(n_59032), .C(n_237291726), .D(nbus_11271
		[1]), .Z(n_289392238));
	notech_ao4 i_113645329(.A(n_56762), .B(n_31612), .C(n_4446), .D(n_59005)
		, .Z(n_289592240));
	notech_ao4 i_113545330(.A(n_57978), .B(n_33713), .C(n_61110), .D(n_32915
		), .Z(n_289692241));
	notech_and4 i_114145324(.A(n_289692241), .B(n_289592240), .C(n_289392238
		), .D(n_289192236), .Z(n_289992243));
	notech_ao4 i_113245333(.A(n_56738), .B(nbus_11270[1]), .C(n_56728), .D(n_33768
		), .Z(n_290092244));
	notech_ao4 i_113145334(.A(n_31525), .B(n_23988), .C(n_56707), .D(n_60510
		), .Z(n_290192245));
	notech_ao4 i_112945336(.A(n_23836), .B(n_33767), .C(n_23989), .D(n_33386
		), .Z(n_290392247));
	notech_and3 i_113045335(.A(n_56750), .B(n_290392247), .C(n_239391747), .Z
		(n_290592249));
	notech_mux2 i_112545340(.S(n_60467), .A(n_236991723), .B(n_237091724), .Z
		(n_290792251));
	notech_ao4 i_112445341(.A(n_4446), .B(n_58956), .C(n_25433), .D(n_59014)
		, .Z(n_290992252));
	notech_ao4 i_112245343(.A(n_61110), .B(n_32914), .C(n_56762), .D(n_31611
		), .Z(n_291192254));
	notech_ao4 i_112145344(.A(n_56728), .B(n_33766), .C(n_57978), .D(n_33714
		), .Z(n_291292255));
	notech_and4 i_112745338(.A(n_291292255), .B(n_291192254), .C(n_290992252
		), .D(n_290792251), .Z(n_291492257));
	notech_ao4 i_111745347(.A(n_56707), .B(n_60519), .C(n_56738), .D(nbus_11270
		[0]), .Z(n_291592258));
	notech_ao4 i_111645348(.A(n_23989), .B(n_33384), .C(n_23988), .D(n_31524
		), .Z(n_291692259));
	notech_ao4 i_111345350(.A(n_23839), .B(n_33765), .C(n_23836), .D(n_33764
		), .Z(n_291892261));
	notech_and4 i_112045345(.A(n_291892261), .B(n_291692259), .C(n_291592258
		), .D(n_56750), .Z(n_292092263));
	notech_or4 i_63743314(.A(n_32244), .B(n_32261), .C(n_32266), .D(n_32273)
		, .Z(n_292192264));
	notech_nand3 i_65143309(.A(n_57467), .B(n_293892281), .C(n_57429), .Z(n_292292265
		));
	notech_and2 i_106742273(.A(imm[30]), .B(n_57236), .Z(n_292392266));
	notech_or2 i_2743250(.A(n_56359), .B(n_60611), .Z(n_293292275));
	notech_nand2 i_38358(.A(n_32244), .B(n_57429), .Z(n_293792280));
	notech_nand2 i_114142199(.A(n_57500), .B(n_57512), .Z(n_293892281));
	notech_ao4 i_218641194(.A(n_55227), .B(n_5758), .C(n_55218), .D(n_31324)
		, .Z(n_294292285));
	notech_ao4 i_218541195(.A(n_57429), .B(n_31028), .C(n_55207), .D(n_31291
		), .Z(n_294392286));
	notech_ao4 i_116242178(.A(n_56350), .B(n_58483), .C(n_4351), .D(n_32911)
		, .Z(n_294492287));
	notech_ao4 i_116142179(.A(n_4348), .B(n_31538), .C(n_56341), .D(n_33814)
		, .Z(n_294692289));
	notech_and3 i_116442176(.A(n_294492287), .B(n_294692289), .C(n_293292275
		), .Z(n_294792290));
	notech_ao4 i_115942181(.A(n_56330), .B(n_33813), .C(n_33812), .D(n_111142552
		), .Z(n_294892291));
	notech_ao4 i_115842182(.A(n_56718), .B(n_33811), .C(n_112042561), .D(n_32344
		), .Z(n_294992292));
	notech_or4 i_152155997(.A(n_32574), .B(n_309960727), .C(n_61076), .D(n_60170
		), .Z(n_295192294));
	notech_nand2 i_8739989(.A(n_57340), .B(n_295592298), .Z(n_295292295));
	notech_and2 i_165155967(.A(n_295192294), .B(n_225391607), .Z(n_295392296
		));
	notech_or4 i_93339173(.A(n_61076), .B(n_61739), .C(n_60170), .D(n_56908)
		, .Z(n_295492297));
	notech_or4 i_107839029(.A(n_61076), .B(n_61739), .C(n_60170), .D(n_4450)
		, .Z(n_295592298));
	notech_or4 i_93139175(.A(n_32628), .B(n_32394), .C(n_60154), .D(n_33815)
		, .Z(n_295692299));
	notech_or4 i_93239174(.A(n_30368), .B(n_156269600), .C(n_27835), .D(n_295392296
		), .Z(n_295792300));
	notech_nao3 i_96139145(.A(mul64[37]), .B(n_61669), .C(n_1861), .Z(n_296692309
		));
	notech_nao3 i_97439132(.A(mul64[38]), .B(n_61669), .C(n_1861), .Z(n_297992322
		));
	notech_nao3 i_98739119(.A(mul64[39]), .B(n_61669), .C(n_1861), .Z(n_299292335
		));
	notech_nand2 i_100339103(.A(n_30422), .B(opb[15]), .Z(n_300192344));
	notech_or4 i_100039106(.A(n_58610), .B(n_32627), .C(n_61618), .D(\nbus_11290[7] 
		), .Z(n_300492347));
	notech_nand2 i_101739089(.A(opc_14[28]), .B(n_61119), .Z(n_301192352));
	notech_nand2 i_101639090(.A(n_30422), .B(opb[28]), .Z(n_301492355));
	notech_nao3 i_101139095(.A(n_30371), .B(n_3677), .C(n_24147), .Z(n_302292360
		));
	notech_and2 i_22666(.A(n_348378486), .B(n_295292295), .Z(n_302392361));
	notech_ao4 i_199838147(.A(n_56738), .B(nbus_11270[28]), .C(n_56707), .D(nbus_11271
		[4]), .Z(n_302492362));
	notech_ao4 i_199738148(.A(n_56774), .B(n_33827), .C(n_57978), .D(n_33715
		), .Z(n_302692364));
	notech_ao4 i_199438151(.A(n_56762), .B(n_31639), .C(n_56923), .D(n_60564
		), .Z(n_302892366));
	notech_and4 i_199638149(.A(n_56750), .B(n_302892366), .C(n_301492355), .D
		(n_301192352), .Z(n_303392369));
	notech_ao4 i_197438169(.A(n_56707), .B(n_60528), .C(n_23989), .D(n_33414
		), .Z(n_303492370));
	notech_ao4 i_197338170(.A(n_56728), .B(n_33826), .C(n_56738), .D(nbus_11270
		[15]), .Z(n_303592371));
	notech_ao4 i_197138172(.A(n_56774), .B(n_33825), .C(n_57978), .D(n_33716
		), .Z(n_303792373));
	notech_and4 i_197738167(.A(n_303792373), .B(n_303592371), .C(n_303492370
		), .D(n_300492347), .Z(n_303992375));
	notech_ao4 i_196838175(.A(n_56762), .B(n_31626), .C(n_25433), .D(n_60591
		), .Z(n_304092376));
	notech_ao4 i_196638177(.A(n_23988), .B(n_31539), .C(n_61110), .D(n_32929
		), .Z(n_304292378));
	notech_and4 i_197038173(.A(n_56750), .B(n_304292378), .C(n_304092376), .D
		(n_300192344), .Z(n_304492380));
	notech_nao3 i_206840060(.A(n_30364), .B(rep_en1), .C(n_4086), .Z(n_304792381
		));
	notech_nao3 i_197640062(.A(n_30364), .B(n_30937), .C(n_4086), .Z(n_304892382
		));
	notech_ao4 i_196238180(.A(n_304892382), .B(n_33824), .C(n_304792381), .D
		(n_33823), .Z(n_304992383));
	notech_ao4 i_196138181(.A(n_56707), .B(n_60591), .C(n_23989), .D(n_33398
		), .Z(n_305092384));
	notech_ao4 i_195938183(.A(n_56728), .B(n_33822), .C(n_56738), .D(nbus_11270
		[7]), .Z(n_305292386));
	notech_and4 i_196438178(.A(n_305292386), .B(n_305092384), .C(n_304992383
		), .D(n_299292335), .Z(n_305492388));
	notech_ao4 i_195638186(.A(n_25433), .B(n_59068), .C(n_56923), .D(nbus_11271
		[7]), .Z(n_305592389));
	notech_ao4 i_195538187(.A(n_4446), .B(\nbus_11290[7] ), .C(n_56762), .D(n_31618
		), .Z(n_305692390));
	notech_ao4 i_195338189(.A(n_23988), .B(n_31531), .C(n_61110), .D(n_32921
		), .Z(n_305892392));
	notech_and4 i_195838184(.A(n_56750), .B(n_305892392), .C(n_305692390), .D
		(n_305592389), .Z(n_306092394));
	notech_ao4 i_195038192(.A(n_304892382), .B(n_33821), .C(n_304792381), .D
		(n_33820), .Z(n_306392395));
	notech_ao4 i_194938193(.A(n_56707), .B(n_60611), .C(n_23989), .D(n_33396
		), .Z(n_306492396));
	notech_ao4 i_194738195(.A(n_56728), .B(n_33819), .C(n_56738), .D(nbus_11270
		[6]), .Z(n_306692398));
	notech_and4 i_195238190(.A(n_306692398), .B(n_306492396), .C(n_306392395
		), .D(n_297992322), .Z(n_306892400));
	notech_ao4 i_194338198(.A(n_25433), .B(n_59041), .C(n_56923), .D(nbus_11271
		[6]), .Z(n_306992401));
	notech_ao4 i_194238199(.A(n_4446), .B(\nbus_11290[6] ), .C(n_56762), .D(n_31617
		), .Z(n_307092402));
	notech_ao4 i_194038201(.A(n_23988), .B(n_31530), .C(n_61110), .D(n_32920
		), .Z(n_307292404));
	notech_and4 i_194638196(.A(n_56750), .B(n_307292404), .C(n_307092402), .D
		(n_306992401), .Z(n_307492406));
	notech_ao4 i_193738204(.A(n_304892382), .B(n_33818), .C(n_304792381), .D
		(n_33817), .Z(n_307592407));
	notech_ao4 i_193638205(.A(n_56707), .B(n_60620), .C(n_23989), .D(n_33394
		), .Z(n_307692408));
	notech_ao4 i_193438207(.A(n_56728), .B(n_33816), .C(n_56738), .D(nbus_11270
		[5]), .Z(n_308092410));
	notech_and4 i_193938202(.A(n_308092410), .B(n_307692408), .C(n_307592407
		), .D(n_296692309), .Z(n_308292412));
	notech_ao4 i_193138210(.A(n_25433), .B(n_58965), .C(n_56923), .D(nbus_11271
		[5]), .Z(n_308392413));
	notech_ao4 i_193038211(.A(n_4446), .B(\nbus_11290[5] ), .C(n_56762), .D(n_31616
		), .Z(n_308492414));
	notech_ao4 i_192838213(.A(n_23988), .B(n_31529), .C(n_61110), .D(n_32919
		), .Z(n_308692416));
	notech_and4 i_193338208(.A(n_56750), .B(n_308692416), .C(n_308492414), .D
		(n_308392413), .Z(n_308892418));
	notech_or4 i_101437773(.A(n_32589), .B(n_28008), .C(n_60154), .D(n_61618
		), .Z(n_309192421));
	notech_ao4 i_15137349(.A(n_35412112), .B(n_19620), .C(n_57001), .D(n_310792435
		), .Z(n_309392423));
	notech_ao4 i_56037729(.A(n_2111), .B(n_310492432), .C(n_2112), .D(n_61621
		), .Z(n_309892426));
	notech_or4 i_106836580(.A(n_61917), .B(n_61903), .C(n_61878), .D(n_60629
		), .Z(n_310492432));
	notech_ao4 i_85236774(.A(n_32952), .B(n_56380), .C(n_59104), .D(n_32950)
		, .Z(n_310592433));
	notech_ao4 i_85136775(.A(n_24298), .B(n_33828), .C(n_56368), .D(n_58974)
		, .Z(n_310692434));
	notech_or4 i_71336882(.A(n_61912), .B(n_61896), .C(n_301760646), .D(n_72112478
		), .Z(n_310792435));
	notech_nand3 i_86595675(.A(vliw_pc[1]), .B(vliw_pc[2]), .C(vliw_pc[0]), 
		.Z(n_310892436));
	notech_nand2 i_47107(.A(n_97890345), .B(n_57724), .Z(n_8771));
	notech_nand2 i_46952(.A(n_97790344), .B(n_57724), .Z(n_8589));
	notech_nand2 i_50842(.A(n_57724), .B(n_97690343), .Z(n_14525));
	notech_nand2 i_47894(.A(n_57724), .B(n_97590342), .Z(n_10088));
	notech_ao4 i_46883(.A(n_295192294), .B(n_230891662), .C(n_57672), .D(n_57041
		), .Z(n_8508));
	notech_nand2 i_50663(.A(n_442468008), .B(n_3456), .Z(n_14184));
	notech_ao4 i_52160(.A(n_33496), .B(n_113590502), .C(n_4402), .D(n_348689368
		), .Z(\nbus_11334[0] ));
	notech_or4 i_47032(.A(n_61669), .B(n_30715), .C(n_61866), .D(n_14216), .Z
		(\nbus_11286[0] ));
	notech_ao4 i_54977(.A(n_61841), .B(n_348271368), .C(n_311071092), .D(n_30364
		), .Z(\nbus_11355[0] ));
	notech_nand2 i_52649(.A(n_57678), .B(n_113490501), .Z(n_17446));
	notech_ao4 i_52263(.A(n_149390860), .B(n_60154), .C(n_311071092), .D(n_30364
		), .Z(n_16862));
	notech_nand2 i_46343(.A(n_57678), .B(n_97090337), .Z(n_7488));
	notech_and4 i_1611982(.A(n_115790524), .B(n_115690523), .C(n_115490521),
		 .D(n_115390520), .Z(to_acu101153[15]));
	notech_and4 i_1711983(.A(n_116390530), .B(n_116290529), .C(n_116090527),
		 .D(n_115990526), .Z(to_acu101153[16]));
	notech_and4 i_1911985(.A(n_116990536), .B(n_116890535), .C(n_116690533),
		 .D(n_116590532), .Z(to_acu101153[18]));
	notech_and4 i_2011986(.A(n_117590542), .B(n_117490541), .C(n_117290539),
		 .D(n_117190538), .Z(to_acu101153[19]));
	notech_and4 i_2111987(.A(n_118190548), .B(n_118090547), .C(n_117890545),
		 .D(n_117790544), .Z(to_acu101153[20]));
	notech_and4 i_2211988(.A(n_118790554), .B(n_118690553), .C(n_118490551),
		 .D(n_118390550), .Z(to_acu101153[21]));
	notech_nand2 i_117983(.A(n_119090557), .B(n_118990556), .Z(write_data_26
		[0]));
	notech_nand2 i_217984(.A(n_119290559), .B(n_119190558), .Z(write_data_26
		[1]));
	notech_nand2 i_317985(.A(n_119490561), .B(n_119390560), .Z(write_data_26
		[2]));
	notech_nand2 i_417986(.A(n_119690563), .B(n_119590562), .Z(write_data_26
		[3]));
	notech_nand2 i_517987(.A(n_119890565), .B(n_119790564), .Z(write_data_26
		[4]));
	notech_nand2 i_617988(.A(n_120090567), .B(n_119990566), .Z(write_data_26
		[5]));
	notech_nand2 i_717989(.A(n_120290569), .B(n_120190568), .Z(write_data_26
		[6]));
	notech_nand2 i_817990(.A(n_120490571), .B(n_120390570), .Z(write_data_26
		[7]));
	notech_nand2 i_917991(.A(n_120690573), .B(n_120590572), .Z(write_data_26
		[8]));
	notech_nand2 i_1017992(.A(n_120890575), .B(n_120790574), .Z(write_data_26
		[9]));
	notech_nand2 i_1517997(.A(n_121090577), .B(n_120990576), .Z(write_data_26
		[14]));
	notech_nand2 i_1717999(.A(n_121290579), .B(n_121190578), .Z(write_data_26
		[16]));
	notech_nand2 i_1818000(.A(n_121490581), .B(n_121390580), .Z(write_data_26
		[17]));
	notech_nand2 i_1918001(.A(n_121690583), .B(n_121590582), .Z(write_data_26
		[18]));
	notech_nand2 i_2018002(.A(n_121890585), .B(n_121790584), .Z(write_data_26
		[19]));
	notech_nand2 i_2118003(.A(n_122090587), .B(n_121990586), .Z(write_data_26
		[20]));
	notech_nand2 i_2218004(.A(n_122290589), .B(n_122190588), .Z(write_data_26
		[21]));
	notech_nand2 i_2318005(.A(n_122490591), .B(n_122390590), .Z(write_data_26
		[22]));
	notech_nand2 i_2418006(.A(n_122690593), .B(n_122590592), .Z(write_data_26
		[23]));
	notech_nand2 i_2518007(.A(n_122890595), .B(n_122790594), .Z(write_data_26
		[24]));
	notech_nand2 i_2618008(.A(n_123090597), .B(n_122990596), .Z(write_data_26
		[25]));
	notech_nand2 i_2718009(.A(n_123290599), .B(n_123190598), .Z(write_data_26
		[26]));
	notech_nand2 i_2818010(.A(n_123490601), .B(n_123390600), .Z(write_data_26
		[27]));
	notech_nand2 i_2918011(.A(n_123690603), .B(n_123590602), .Z(write_data_26
		[28]));
	notech_nand2 i_3218014(.A(n_123890605), .B(n_123790604), .Z(write_data_26
		[31]));
	notech_ao4 i_5969204(.A(n_288144316), .B(n_189162918), .C(n_323160859), 
		.D(n_33162), .Z(n_163262664));
	notech_or4 i_7069193(.A(instrc[127]), .B(instrc[125]), .C(n_163262664), 
		.D(n_33175), .Z(n_163162663));
	notech_or2 i_50692(.A(n_56734), .B(n_30722), .Z(n_14216));
	notech_and4 i_5869205(.A(n_322760855), .B(n_322860856), .C(n_188862915),
		 .D(n_162662658), .Z(n_163062662));
	notech_nao3 i_5669207(.A(n_323060858), .B(n_162762659), .C(n_322960857),
		 .Z(n_162962661));
	notech_nand3 i_5769206(.A(n_57595), .B(n_57081), .C(n_63762), .Z(n_162762659
		));
	notech_nand2 i_5569208(.A(n_57086), .B(n_57595), .Z(n_162662658));
	notech_nao3 i_4969214(.A(n_61953), .B(n_63762), .C(n_26957), .Z(n_162462656
		));
	notech_ao4 i_124969291(.A(n_63768), .B(n_61953), .C(n_26957), .D(n_61052
		), .Z(n_162262654));
	notech_and4 i_40571575(.A(n_161862650), .B(n_158762619), .C(n_158962621)
		, .D(n_158862620), .Z(n_161962651));
	notech_and4 i_40471576(.A(n_158562617), .B(n_161562647), .C(n_158662618)
		, .D(n_159062622), .Z(n_161862650));
	notech_ao4 i_39971581(.A(n_376464295), .B(n_61841), .C(n_57068), .D(n_114845640
		), .Z(n_161562647));
	notech_nao3 i_16994(.A(n_63718), .B(n_63762), .C(n_149390860), .Z(n_310992437
		));
	notech_ao3 i_16987(.A(calc_sz[1]), .B(n_57651), .C(n_348789369), .Z(n_311292438
		));
	notech_and4 i_17002(.A(n_25665), .B(n_63818), .C(n_61824), .D(n_30898), 
		.Z(n_311392439));
	notech_and2 i_17456(.A(n_125190618), .B(regs_10[0]), .Z(n_311492440));
	notech_and2 i_17457(.A(n_125190618), .B(regs_10[1]), .Z(n_311592441));
	notech_and2 i_17458(.A(n_125190618), .B(regs_10[2]), .Z(n_311692442));
	notech_and2 i_17459(.A(regs_10[3]), .B(n_125190618), .Z(n_311792443));
	notech_and2 i_17460(.A(n_125190618), .B(regs_10[4]), .Z(n_311892444));
	notech_and2 i_17461(.A(n_125190618), .B(regs_10[5]), .Z(n_311992445));
	notech_and2 i_17462(.A(n_125190618), .B(regs_10[6]), .Z(n_312092446));
	notech_and2 i_17463(.A(n_125190618), .B(regs_10[7]), .Z(n_312192447));
	notech_and2 i_17464(.A(n_125190618), .B(regs_10[8]), .Z(n_312292448));
	notech_and2 i_17465(.A(n_125190618), .B(regs_10[9]), .Z(n_312392449));
	notech_and2 i_17466(.A(n_125190618), .B(regs_10[10]), .Z(n_312492450));
	notech_and2 i_17467(.A(n_125190618), .B(regs_10[11]), .Z(n_312592451));
	notech_and2 i_17468(.A(n_125190618), .B(regs_10[12]), .Z(n_312792452));
	notech_and2 i_17469(.A(n_125190618), .B(regs_10[13]), .Z(n_312892453));
	notech_and2 i_17470(.A(n_125190618), .B(regs_10[14]), .Z(n_312992454));
	notech_and2 i_17471(.A(n_125190618), .B(regs_10[15]), .Z(n_313192455));
	notech_and2 i_17472(.A(n_54412), .B(regs_10[16]), .Z(n_313392456));
	notech_and2 i_17473(.A(n_54412), .B(regs_10[17]), .Z(n_313592457));
	notech_and2 i_17474(.A(n_54412), .B(regs_10[18]), .Z(n_313792458));
	notech_and2 i_17475(.A(n_54412), .B(regs_10[19]), .Z(n_313892459));
	notech_and2 i_17476(.A(n_54412), .B(regs_10[20]), .Z(n_313992460));
	notech_and2 i_17477(.A(n_54412), .B(regs_10[21]), .Z(n_314092461));
	notech_and2 i_17478(.A(n_54412), .B(regs_10[22]), .Z(n_314192462));
	notech_and2 i_17479(.A(n_54412), .B(regs_10[23]), .Z(n_314492463));
	notech_and2 i_17480(.A(n_54412), .B(regs_10[24]), .Z(n_314592464));
	notech_and2 i_17481(.A(n_54412), .B(regs_10[25]), .Z(n_314692465));
	notech_and2 i_17482(.A(n_54412), .B(regs_10[26]), .Z(n_314792466));
	notech_and2 i_17483(.A(n_54412), .B(regs_10[27]), .Z(n_314892467));
	notech_and2 i_17484(.A(n_54412), .B(regs_10[28]), .Z(n_314992468));
	notech_and2 i_17485(.A(n_54412), .B(regs_10[29]), .Z(n_315092469));
	notech_and2 i_17486(.A(n_54412), .B(regs_10[30]), .Z(n_315192470));
	notech_and2 i_17487(.A(n_54412), .B(regs_10[31]), .Z(n_315292471));
	notech_ao3 i_17932(.A(tcmp_arithbox), .B(n_61670), .C(n_27914), .Z(n_315392472
		));
	notech_and3 i_22830(.A(n_61670), .B(n_30935), .C(n_125290619), .Z(n_315492473
		));
	notech_ao3 i_22832(.A(n_128090647), .B(n_61670), .C(n_1849), .Z(n_315592474
		));
	notech_nor2 i_26417(.A(n_315892477), .B(n_61621), .Z(n_315692475));
	notech_or4 i_26423(.A(n_61797), .B(n_32628), .C(n_60170), .D(n_61841), .Z
		(n_315792476));
	notech_and2 i_3471930(.A(n_30560), .B(n_30341), .Z(n_315892477));
	notech_ao4 i_57669314(.A(n_2112), .B(n_61621), .C(n_60602), .D(n_56422),
		 .Z(n_315992478));
	notech_and4 i_121759(.A(n_192891288), .B(n_193091290), .C(n_190791267), 
		.D(n_192791287), .Z(n_15170));
	notech_ao4 i_8432(.A(n_193491294), .B(n_311371095), .C(n_61866), .D(n_61618
		), .Z(n_18354));
	notech_ao4 i_3015644(.A(n_55588), .B(n_31537), .C(n_55579), .D(n_31961),
		 .Z(n_14482));
	notech_nand2 i_323090(.A(n_213333664), .B(n_213091485), .Z(n_11287));
	notech_ao4 i_223089(.A(n_213333664), .B(n_59005), .C(n_213091485), .D(n_56956
		), .Z(n_11281));
	notech_ao4 i_123088(.A(n_213333664), .B(n_58956), .C(n_213091485), .D(n_56965
		), .Z(n_11275));
	notech_nand3 i_3218814(.A(n_213191486), .B(n_213391488), .C(n_212591483)
		, .Z(n_20999));
	notech_nand3 i_3118813(.A(n_213491489), .B(n_213691491), .C(n_212091478)
		, .Z(n_20994));
	notech_nand3 i_3018812(.A(n_213791492), .B(n_213991494), .C(n_211591473)
		, .Z(n_20989));
	notech_nand3 i_2918811(.A(n_214191495), .B(n_214391497), .C(n_211091468)
		, .Z(n_20984));
	notech_nand3 i_2818810(.A(n_214491498), .B(n_214691500), .C(n_210591463)
		, .Z(n_20979));
	notech_nand3 i_2718809(.A(n_214791501), .B(n_214991503), .C(n_210091458)
		, .Z(n_20974));
	notech_nao3 i_2618808(.A(n_215091504), .B(n_215291506), .C(n_209591453),
		 .Z(n_20969));
	notech_nao3 i_2518807(.A(n_215391507), .B(n_215591509), .C(n_208991448),
		 .Z(n_20964));
	notech_nand3 i_2418806(.A(n_215691510), .B(n_215891512), .C(n_208491443)
		, .Z(n_20959));
	notech_nao3 i_2318805(.A(n_215991513), .B(n_216191515), .C(n_207991438),
		 .Z(n_20954));
	notech_nand3 i_2218804(.A(n_216291516), .B(n_216491518), .C(n_207491433)
		, .Z(n_20949));
	notech_nao3 i_2118803(.A(n_216591519), .B(n_216791521), .C(n_206991428),
		 .Z(n_20944));
	notech_nand3 i_2018802(.A(n_216891522), .B(n_217091524), .C(n_206491423)
		, .Z(n_20939));
	notech_nand3 i_1918801(.A(n_217191525), .B(n_217391527), .C(n_205991418)
		, .Z(n_20934));
	notech_nand3 i_1818800(.A(n_217491528), .B(n_217691530), .C(n_205491413)
		, .Z(n_20929));
	notech_nand3 i_1718799(.A(n_217791531), .B(n_217991533), .C(n_204991408)
		, .Z(n_20924));
	notech_nand3 i_1618798(.A(n_218091534), .B(n_218291536), .C(n_204491403)
		, .Z(n_20919));
	notech_nand3 i_1518797(.A(n_218391537), .B(n_218591539), .C(n_203991398)
		, .Z(n_20914));
	notech_nand3 i_1418796(.A(n_218691540), .B(n_218891542), .C(n_203491393)
		, .Z(n_20909));
	notech_nand3 i_1318795(.A(n_218991543), .B(n_219191545), .C(n_202991388)
		, .Z(n_20904));
	notech_nand3 i_1218794(.A(n_219291546), .B(n_219491548), .C(n_202491383)
		, .Z(n_20899));
	notech_nand3 i_1118793(.A(n_219591549), .B(n_219791551), .C(n_201991378)
		, .Z(n_20894));
	notech_nand3 i_1018792(.A(n_219891552), .B(n_220091554), .C(n_201391373)
		, .Z(n_20889));
	notech_nand3 i_918791(.A(n_220191555), .B(n_220391557), .C(n_200891368),
		 .Z(n_20884));
	notech_nand3 i_818790(.A(n_220491558), .B(n_220691560), .C(n_200391363),
		 .Z(n_20879));
	notech_nand3 i_718789(.A(n_220791561), .B(n_220991563), .C(n_199891358),
		 .Z(n_20874));
	notech_nand3 i_618788(.A(n_221091564), .B(n_221291566), .C(n_199391353),
		 .Z(n_20869));
	notech_nand3 i_518787(.A(n_221391567), .B(n_221591569), .C(n_198891348),
		 .Z(n_20864));
	notech_nand3 i_418786(.A(n_221691570), .B(n_221891572), .C(n_198391343),
		 .Z(n_20859));
	notech_nand3 i_318785(.A(n_221991573), .B(n_222191575), .C(n_197891338),
		 .Z(n_20854));
	notech_nand3 i_218784(.A(n_222291576), .B(n_222491578), .C(n_197391333),
		 .Z(n_20849));
	notech_nand3 i_118783(.A(n_222591579), .B(n_222791581), .C(n_196891328),
		 .Z(n_20844));
	notech_or4 i_218944(.A(n_196091320), .B(n_223091584), .C(n_30684), .D(n_223891592
		), .Z(n_20634));
	notech_ao4 i_50702(.A(n_61841), .B(n_284331524), .C(n_295192294), .D(n_230891662
		), .Z(n_14229));
	notech_or4 i_202555926(.A(n_32574), .B(n_32184), .C(n_32396), .D(n_60170
		), .Z(n_284331524));
	notech_or4 i_6346(.A(n_226191615), .B(n_226291616), .C(n_235791711), .D(n_30692
		), .Z(n_7418));
	notech_ao4 i_6408(.A(n_447068054), .B(n_295192294), .C(CFOF_mul), .D(n_284331524
		), .Z(n_14232));
	notech_and2 i_17804(.A(n_235891712), .B(n_30654), .Z(n_316092479));
	notech_and2 i_17805(.A(n_235991713), .B(n_30654), .Z(n_316192480));
	notech_and2 i_17806(.A(n_236091714), .B(n_30654), .Z(n_316292481));
	notech_nor2 i_17807(.A(n_236191715), .B(n_353728636), .Z(n_316392482));
	notech_and4 i_3217182(.A(n_266192011), .B(n_266392013), .C(n_266892018),
		 .D(n_266092010), .Z(n_9971));
	notech_and4 i_3117181(.A(n_266992019), .B(n_267192021), .C(n_267692026),
		 .D(n_265192001), .Z(n_9966));
	notech_and4 i_3017180(.A(n_267792027), .B(n_267992029), .C(n_268492034),
		 .D(n_264291992), .Z(n_9961));
	notech_and4 i_2817178(.A(n_268592035), .B(n_268792037), .C(n_269292042),
		 .D(n_263391983), .Z(n_9951));
	notech_and4 i_2717177(.A(n_269392043), .B(n_269592045), .C(n_270092050),
		 .D(n_262491974), .Z(n_9946));
	notech_and4 i_2617176(.A(n_270192051), .B(n_270392053), .C(n_271092058),
		 .D(n_261591965), .Z(n_9941));
	notech_and4 i_2517175(.A(n_271192059), .B(n_271392061), .C(n_271892066),
		 .D(n_260691956), .Z(n_9936));
	notech_and4 i_2417174(.A(n_271992067), .B(n_272192069), .C(n_272692074),
		 .D(n_259791947), .Z(n_9931));
	notech_and4 i_2317173(.A(n_272792075), .B(n_272992077), .C(n_273492082),
		 .D(n_258891938), .Z(n_9926));
	notech_and4 i_2217172(.A(n_273592083), .B(n_273792085), .C(n_274292090),
		 .D(n_257991929), .Z(n_9921));
	notech_and4 i_2117171(.A(n_274392091), .B(n_274592093), .C(n_275092098),
		 .D(n_257091920), .Z(n_9916));
	notech_and4 i_2017170(.A(n_275192099), .B(n_275392101), .C(n_276092106),
		 .D(n_256191911), .Z(n_9911));
	notech_and4 i_1917169(.A(n_276192107), .B(n_276392109), .C(n_276892114),
		 .D(n_255291902), .Z(n_9906));
	notech_and4 i_1817168(.A(n_276992115), .B(n_277192117), .C(n_277692122),
		 .D(n_254391893), .Z(n_9901));
	notech_and4 i_1717167(.A(n_277792123), .B(n_277992125), .C(n_278492130),
		 .D(n_253491884), .Z(n_9896));
	notech_nand2 i_1517165(.A(n_279592141), .B(n_279092136), .Z(n_9886));
	notech_nand2 i_1417164(.A(n_280692152), .B(n_280192147), .Z(n_9881));
	notech_nand2 i_1317163(.A(n_281792163), .B(n_281292158), .Z(n_9876));
	notech_nand2 i_1217162(.A(n_282892174), .B(n_282392169), .Z(n_9871));
	notech_nand2 i_1117161(.A(n_283992185), .B(n_283492180), .Z(n_9866));
	notech_nand2 i_1017160(.A(n_285092196), .B(n_284592191), .Z(n_9861));
	notech_nand2 i_917159(.A(n_286192207), .B(n_285692202), .Z(n_9856));
	notech_and4 i_417154(.A(n_287092216), .B(n_286992215), .C(n_286892214), 
		.D(n_287592220), .Z(n_9831));
	notech_nand2 i_317153(.A(n_288992234), .B(n_288392228), .Z(n_9826));
	notech_and4 i_217152(.A(n_290192245), .B(n_290092244), .C(n_289992243), 
		.D(n_290592249), .Z(n_9821));
	notech_nand2 i_117151(.A(n_292092263), .B(n_291492257), .Z(n_9816));
	notech_nand2 i_3118013(.A(n_294392286), .B(n_294292285), .Z(write_data_26
		[30]));
	notech_or2 i_20243360(.A(n_57024), .B(n_292392266), .Z(\nbus_11309[30] )
		);
	notech_nand3 i_3112925(.A(n_294992292), .B(n_294892291), .C(n_294792290)
		, .Z(n_21457));
	notech_or2 i_73940115(.A(n_331960947), .B(n_336460992), .Z(n_57742));
	notech_nand3 i_7023(.A(n_295792300), .B(n_295692299), .C(n_295492297), .Z
		(n_16833));
	notech_and4 i_2917179(.A(n_302492362), .B(n_302692364), .C(n_303392369),
		 .D(n_302292360), .Z(n_9956));
	notech_nand2 i_1617166(.A(n_304492380), .B(n_303992375), .Z(n_9891));
	notech_nand2 i_817158(.A(n_306092394), .B(n_305492388), .Z(n_9851));
	notech_nand2 i_717157(.A(n_307492406), .B(n_306892400), .Z(n_9846));
	notech_nand2 i_617156(.A(n_308892418), .B(n_308292412), .Z(n_9841));
	notech_and4 i_25171728(.A(n_156862600), .B(n_159962631), .C(n_156562597)
		, .D(n_160362635), .Z(n_160662638));
	notech_nand2 i_35097(.A(n_19707), .B(n_61618), .Z(n_2140));
	notech_ao4 i_8449(.A(n_309392423), .B(n_19725), .C(n_61866), .D(n_61618)
		, .Z(n_9190));
	notech_nand2 i_1227479(.A(n_310692434), .B(n_310592433), .Z(n_7839));
	notech_and3 i_24771732(.A(n_160162633), .B(n_160062632), .C(n_156462596)
		, .Z(n_160362635));
	notech_ao4 i_24571734(.A(n_111445606), .B(n_57622), .C(n_57609), .D(n_114845640
		), .Z(n_160162633));
	notech_ao4 i_24471735(.A(n_61841), .B(n_32181), .C(n_375564286), .D(n_375664287
		), .Z(n_160062632));
	notech_ao4 i_24971730(.A(n_155862590), .B(n_30550), .C(n_155762589), .D(n_30551
		), .Z(n_159962631));
	notech_or4 i_22771752(.A(instrc[102]), .B(n_322060848), .C(n_30550), .D(instrc
		[101]), .Z(n_159862630));
	notech_or4 i_22171758(.A(instrc[125]), .B(n_376064291), .C(instrc[126]),
		 .D(n_33153), .Z(n_159762629));
	notech_nand2 i_6871896(.A(n_33179), .B(instrc[88]), .Z(n_159662628));
	notech_nand2 i_6771897(.A(n_33177), .B(instrc[92]), .Z(n_159562627));
	notech_nao3 i_4271922(.A(instrc[96]), .B(instrc[99]), .C(n_30617), .Z(n_159462626
		));
	notech_and4 i_49550(.A(n_159162623), .B(n_161962651), .C(n_159262624), .D
		(n_30881), .Z(n_159362625));
	notech_nand2 i_39071590(.A(n_157962611), .B(n_26063), .Z(n_159262624));
	notech_or2 i_38971591(.A(n_1460), .B(n_157862610), .Z(n_159162623));
	notech_nao3 i_38671594(.A(n_33157), .B(n_1464), .C(n_375664287), .Z(n_159062622
		));
	notech_nao3 i_38871592(.A(n_26063), .B(n_63762), .C(n_157762609), .Z(n_158962621
		));
	notech_or4 i_39471586(.A(n_1462), .B(n_30551), .C(instrc[103]), .D(n_29584
		), .Z(n_158862620));
	notech_or4 i_39371587(.A(n_322660854), .B(n_30551), .C(instrc[99]), .D(n_29572
		), .Z(n_158762619));
	notech_or4 i_38771593(.A(n_323160859), .B(n_30552), .C(n_33162), .D(instrc
		[127]), .Z(n_158662618));
	notech_or4 i_39271588(.A(instrc[123]), .B(n_111445606), .C(n_318060808),
		 .D(n_61757), .Z(n_158562617));
	notech_ao4 i_39171589(.A(n_241746909), .B(n_157662608), .C(n_376264293),
		 .D(n_30886), .Z(n_158062612));
	notech_nao3 i_38071600(.A(n_323060858), .B(n_157562607), .C(n_322960857)
		, .Z(n_157962611));
	notech_ao4 i_37771603(.A(n_159662628), .B(n_1466), .C(n_159562627), .D(n_1465
		), .Z(n_157862610));
	notech_ao4 i_37571605(.A(n_57633), .B(n_2810), .C(n_30798), .D(n_32210),
		 .Z(n_157762609));
	notech_ao4 i_38371597(.A(n_321860846), .B(n_30547), .C(n_58716), .D(n_2845
		), .Z(n_157662608));
	notech_nand3 i_38171599(.A(n_57595), .B(n_57072), .C(n_63762), .Z(n_157562607
		));
	notech_or4 i_37371607(.A(n_30552), .B(n_376364294), .C(instrc[127]), .D(n_30310
		), .Z(n_157162603));
	notech_ao3 i_52004(.A(n_160662638), .B(n_155962591), .C(n_156962601), .Z
		(n_157062602));
	notech_and2 i_23971740(.A(n_241746909), .B(n_30890), .Z(n_156962601));
	notech_nao3 i_23871741(.A(n_286063762), .B(n_241346905), .C(n_57696), .Z
		(n_156862600));
	notech_or4 i_24071739(.A(n_57696), .B(n_155662588), .C(n_61933), .D(n_30733
		), .Z(n_156562597));
	notech_or4 i_23771742(.A(n_323160859), .B(n_79112547), .C(n_33162), .D(n_33153
		), .Z(n_156462596));
	notech_ao4 i_23171748(.A(n_155562587), .B(n_114845640), .C(n_322560853),
		 .D(n_30319), .Z(n_156062592));
	notech_nand2 i_24371736(.A(n_57609), .B(n_30895), .Z(n_155962591));
	notech_ao4 i_22871751(.A(n_159562627), .B(n_375464285), .C(n_159662628),
		 .D(n_375364284), .Z(n_155862590));
	notech_ao4 i_22471755(.A(n_159862630), .B(n_33142), .C(n_375164282), .D(n_159462626
		), .Z(n_155762589));
	notech_ao4 i_22271757(.A(n_57633), .B(n_2810), .C(n_30798), .D(n_32227),
		 .Z(n_155662588));
	notech_ao4 i_2671938(.A(n_57622), .B(n_285763759), .C(n_159762629), .D(n_30310
		), .Z(n_155562587));
	notech_ao4 i_133373204(.A(n_375064281), .B(n_55227), .C(n_55218), .D(n_31307
		), .Z(n_154662578));
	notech_ao4 i_133473203(.A(n_55207), .B(n_31274), .C(n_57429), .D(n_30993
		), .Z(n_154562577));
	notech_ao4 i_133973198(.A(n_353164063), .B(n_55227), .C(n_55218), .D(n_31304
		), .Z(n_154462576));
	notech_ao4 i_134073197(.A(n_55207), .B(n_31271), .C(n_57429), .D(n_30987
		), .Z(n_154362575));
	notech_ao4 i_99074839(.A(n_56003), .B(n_30975), .C(n_30753), .D(n_31298)
		, .Z(n_153462566));
	notech_ao4 i_99174838(.A(n_20898), .B(n_31615), .C(n_20897), .D(n_31265)
		, .Z(n_153362565));
	notech_nand3 i_26427(.A(n_61775), .B(n_61815), .C(n_30898), .Z(n_32390)
		);
	notech_ao4 i_1754(.A(n_60170), .B(n_25485), .C(n_26637), .D(n_32627), .Z
		(n_23350));
	notech_and4 i_1558(.A(n_58532), .B(n_57662), .C(n_61670), .D(n_27923), .Z
		(n_22746));
	notech_nao3 i_1321(.A(n_58532), .B(n_61670), .C(n_58523), .Z(n_22968));
	notech_nand2 i_1006(.A(n_61775), .B(n_63800), .Z(n_32574));
	notech_nor2 i_1003(.A(n_32396), .B(n_59120), .Z(n_27933));
	notech_ao3 i_997(.A(fsm[3]), .B(fsm[2]), .C(fsm[4]), .Z(n_32536));
	notech_nand2 i_993(.A(n_63818), .B(n_61815), .Z(n_32628));
	notech_nao3 i_992(.A(n_32663), .B(n_30899), .C(n_61076), .Z(n_25681));
	notech_or4 i_961(.A(n_32663), .B(n_309860726), .C(n_312460752), .D(n_30900
		), .Z(n_32394));
	notech_nand2 i_940(.A(n_31258), .B(vliw_pc[3]), .Z(n_32756));
	notech_nor2 i_93975835(.A(n_61907), .B(n_31251), .Z(n_32520));
	notech_nor2 i_90975834(.A(n_32589), .B(n_61065), .Z(n_28097));
	notech_nand2 i_859(.A(n_2952), .B(n_30901), .Z(n_32396));
	notech_and3 i_551(.A(n_19707), .B(n_30307), .C(n_32487), .Z(n_32485));
	notech_or4 i_547(.A(n_32184), .B(n_61076), .C(\opcode[0] ), .D(n_61815),
		 .Z(n_25676));
	notech_or4 i_539(.A(n_312460752), .B(n_32574), .C(n_309960727), .D(n_30900
		), .Z(n_27924));
	notech_nao3 i_525(.A(n_63818), .B(n_61815), .C(n_309960727), .Z(n_32627)
		);
	notech_nao3 i_467(.A(n_61775), .B(n_61815), .C(n_309960727), .Z(n_28098)
		);
	notech_nand2 i_421(.A(n_61775), .B(n_61815), .Z(n_32391));
	notech_nand2 i_418(.A(n_32663), .B(n_30899), .Z(n_32184));
	notech_and3 i_209(.A(n_61775), .B(n_63800), .C(n_30898), .Z(n_32388));
	notech_or4 i_1613(.A(n_309960727), .B(n_32396), .C(n_63800), .D(1'b0), .Z
		(n_27914));
	notech_or2 i_51575(.A(n_301560644), .B(n_301960648), .Z(n_19707));
	notech_nao3 i_51584(.A(n_61907), .B(n_32536), .C(n_61896), .Z(n_19655)
		);
	notech_nor2 i_51587(.A(n_317460802), .B(n_30304), .Z(n_19637));
	notech_and4 i_51751(.A(fsm[4]), .B(fsm[2]), .C(n_31254), .D(n_32520), .Z
		(n_19620));
	notech_and2 i_51582(.A(n_32536), .B(n_61730), .Z(n_19663));
	notech_or4 i_36656(.A(n_61907), .B(n_61896), .C(n_61878), .D(n_1844), .Z
		(n_22742));
	notech_or4 i_36653(.A(n_61907), .B(n_61896), .C(n_61883), .D(n_1799), .Z
		(n_22745));
	notech_nand3 i_1168(.A(n_58532), .B(n_27826), .C(n_57662), .Z(n_22752)
		);
	notech_nand3 i_740(.A(n_58532), .B(n_27923), .C(n_32321), .Z(n_1799));
	notech_or2 i_36431(.A(n_23341), .B(n_30521), .Z(n_22967));
	notech_or4 i_36422(.A(n_61907), .B(n_61896), .C(n_61883), .D(n_1803), .Z
		(n_22976));
	notech_or4 i_36421(.A(n_61907), .B(n_61896), .C(n_61883), .D(n_1804), .Z
		(n_22977));
	notech_or4 i_36419(.A(n_32574), .B(n_25681), .C(n_60154), .D(n_61618), .Z
		(n_22979));
	notech_or4 i_36418(.A(n_61907), .B(n_61896), .C(n_61883), .D(n_1802), .Z
		(n_22980));
	notech_or4 i_36414(.A(n_61907), .B(n_61896), .C(n_61883), .D(n_1801), .Z
		(n_22984));
	notech_or4 i_36413(.A(n_61907), .B(n_61896), .C(n_61883), .D(n_1800), .Z
		(n_22985));
	notech_or4 i_692(.A(n_63698), .B(n_32390), .C(n_61933), .D(n_57662), .Z(n_1800
		));
	notech_or4 i_687(.A(n_32396), .B(n_59120), .C(n_60169), .D(n_58532), .Z(n_1801
		));
	notech_or2 i_686(.A(n_58523), .B(n_27843), .Z(n_1802));
	notech_or4 i_685(.A(n_63718), .B(n_32390), .C(n_61933), .D(n_58532), .Z(n_1803
		));
	notech_nand2 i_684(.A(n_30521), .B(n_27923), .Z(n_1804));
	notech_or4 i_1776(.A(n_32574), .B(n_25681), .C(n_63700), .D(n_63762), .Z
		(n_1805));
	notech_or4 i_1499(.A(n_32628), .B(n_61748), .C(n_61076), .D(n_61052), .Z
		(n_23326));
	notech_nand3 i_36069(.A(n_27823), .B(n_30364), .C(n_317260800), .Z(n_23329
		));
	notech_and4 i_36068(.A(sign_div), .B(n_315760785), .C(opd[31]), .D(n_61730
		), .Z(n_23330));
	notech_nao3 i_36064(.A(n_24147), .B(n_315760785), .C(n_61718), .Z(n_23334
		));
	notech_or4 i_36057(.A(n_61907), .B(n_61896), .C(n_61883), .D(n_27920), .Z
		(n_23341));
	notech_or4 i_36053(.A(n_61907), .B(n_61896), .C(n_61883), .D(n_2852), .Z
		(n_23345));
	notech_nand2 i_1411(.A(n_1823), .B(n_338861016), .Z(n_1806));
	notech_nor2 i_36047(.A(n_58501), .B(n_58561), .Z(n_23351));
	notech_or4 i_36045(.A(instrc[123]), .B(n_61964), .C(n_318160809), .D(n_58501
		), .Z(n_23353));
	notech_or4 i_36039(.A(n_58501), .B(n_32241), .C(n_32249), .D(n_58601), .Z
		(n_23359));
	notech_or4 i_36031(.A(n_32589), .B(n_59120), .C(n_60169), .D(n_61618), .Z
		(n_23367));
	notech_or4 i_1703(.A(n_32589), .B(n_59120), .C(n_63762), .D(n_61953), .Z
		(n_1807));
	notech_or4 i_1492(.A(n_25485), .B(n_63700), .C(n_61933), .D(n_61618), .Z
		(n_23371));
	notech_or4 i_1758(.A(n_32628), .B(n_25681), .C(n_63700), .D(n_61924), .Z
		(n_1808));
	notech_or4 i_1314(.A(n_32574), .B(n_25681), .C(n_61052), .D(n_61618), .Z
		(n_23373));
	notech_or4 i_1809(.A(n_32574), .B(n_25681), .C(n_61924), .D(n_61953), .Z
		(n_1809));
	notech_or4 i_694(.A(n_32589), .B(n_61739), .C(n_60189), .D(n_61614), .Z(n_23379
		));
	notech_or4 i_36015(.A(instrc[123]), .B(n_318060808), .C(n_58501), .D(instrc
		[120]), .Z(n_23383));
	notech_nand2 i_36009(.A(n_58570), .B(n_58561), .Z(n_23389));
	notech_nand2 i_1485(.A(sign_div), .B(opd[31]), .Z(n_24147));
	notech_ao4 i_558(.A(n_339661024), .B(n_32627), .C(n_61065), .D(n_26637),
		 .Z(n_25467));
	notech_ao4 i_1317(.A(n_32627), .B(n_25713), .C(n_61065), .D(n_339661024)
		, .Z(n_25468));
	notech_or4 i_543(.A(n_32184), .B(n_61076), .C(n_61775), .D(\opcode[3] ),
		 .Z(n_25485));
	notech_nand2 i_33749(.A(n_30691), .B(n_30364), .Z(n_25649));
	notech_nand3 i_33728(.A(n_1839), .B(rep_en2), .C(n_30364), .Z(n_25670)
		);
	notech_or4 i_538(.A(n_32184), .B(n_61076), .C(\opcode[0] ), .D(\opcode[3] 
		), .Z(n_25680));
	notech_or4 i_33685(.A(n_2952), .B(n_30901), .C(n_63762), .D(n_61953), .Z
		(n_25713));
	notech_or4 i_532(.A(n_2952), .B(n_30901), .C(n_61924), .D(n_61953), .Z(n_26637
		));
	notech_or4 i_31584(.A(n_61907), .B(n_61896), .C(n_61885), .D(n_27914), .Z
		(n_27814));
	notech_and2 i_210004(.A(n_1839), .B(rep_en2), .Z(n_27823));
	notech_nor2 i_31572(.A(n_27922), .B(n_61614), .Z(n_27826));
	notech_and2 i_1437(.A(n_58532), .B(n_57662), .Z(n_27842));
	notech_or4 i_531(.A(calc_sz[0]), .B(calc_sz[3]), .C(calc_sz[1]), .D(n_31374
		), .Z(n_27843));
	notech_or4 i_1650(.A(n_32574), .B(n_61748), .C(n_32396), .D(n_60169), .Z
		(n_27919));
	notech_or4 i_1637(.A(n_32383), .B(n_61748), .C(n_32396), .D(n_60169), .Z
		(n_27920));
	notech_or4 i_1717(.A(n_32391), .B(n_63700), .C(n_61924), .D(n_32394), .Z
		(n_27922));
	notech_ao3 i_1620(.A(n_61953), .B(n_61924), .C(n_27924), .Z(n_27923));
	notech_or4 i_31309(.A(n_61907), .B(n_61896), .C(n_61885), .D(n_1849), .Z
		(n_28089));
	notech_nand2 i_959(.A(n_1858), .B(n_1857), .Z(n_28092));
	notech_nand2 i_27148(.A(n_32161), .B(n_61757), .Z(n_32250));
	notech_ao3 i_51576(.A(n_61907), .B(n_61896), .C(n_301960648), .Z(n_19698
		));
	notech_or4 i_51578(.A(fsm[4]), .B(fsm[2]), .C(n_31254), .D(n_61718), .Z(n_19689
		));
	notech_ao3 i_51572(.A(n_61912), .B(n_61898), .C(n_61885), .Z(n_19725));
	notech_nor2 i_51570(.A(n_30304), .B(n_61885), .Z(n_19734));
	notech_ao4 i_26911(.A(n_30304), .B(n_61883), .C(n_301960648), .D(n_61718
		), .Z(n_32487));
	notech_ao3 i_51579(.A(n_61912), .B(n_315760785), .C(n_61898), .Z(n_19680
		));
	notech_nand3 i_51581(.A(n_61912), .B(n_61898), .C(n_315760785), .Z(n_19672
		));
	notech_and2 i_26890(.A(n_19672), .B(n_30524), .Z(n_32508));
	notech_nao3 i_51754(.A(n_61912), .B(n_61898), .C(n_301760646), .Z(n_19603
		));
	notech_and3 i_26877(.A(n_19612), .B(n_30636), .C(n_30714), .Z(n_32521)
		);
	notech_nor2 i_51585(.A(n_317460802), .B(n_61718), .Z(n_19645));
	notech_and3 i_51764(.A(n_61912), .B(n_61898), .C(n_32536), .Z(n_19548)
		);
	notech_or4 i_1453(.A(n_32628), .B(n_61748), .C(n_61076), .D(n_60154), .Z
		(n_32590));
	notech_and2 i_987(.A(vliw_pc[1]), .B(n_31256), .Z(n_1816));
	notech_and2 i_857(.A(vliw_pc[1]), .B(vliw_pc[0]), .Z(n_32779));
	notech_or4 i_2131(.A(n_312460752), .B(n_32663), .C(n_2952), .D(n_30899),
		 .Z(n_1817));
	notech_or4 i_1739(.A(n_32391), .B(n_25681), .C(n_63762), .D(n_61958), .Z
		(n_1820));
	notech_or4 i_9425(.A(n_61797), .B(n_60169), .C(\opcode[0] ), .D(n_61815)
		, .Z(n_1823));
	notech_or4 i_9223(.A(n_61748), .B(n_25713), .C(n_61775), .D(\opcode[3] )
		, .Z(n_1824));
	notech_mux2 i_577(.S(n_61665), .A(n_30324), .B(n_23326), .Z(n_1826));
	notech_ao4 i_1123(.A(n_25649), .B(n_30926), .C(n_316760795), .D(n_61614)
		, .Z(n_1827));
	notech_ao4 i_1124(.A(n_30364), .B(n_30926), .C(n_32590), .D(n_61614), .Z
		(n_1828));
	notech_or4 i_1625(.A(n_61912), .B(n_61898), .C(n_61883), .D(n_2974), .Z(n_1832
		));
	notech_or4 i_2040(.A(n_61748), .B(n_339661024), .C(\opcode[0] ), .D(\opcode[3] 
		), .Z(n_1834));
	notech_or4 i_1752(.A(n_32391), .B(n_25681), .C(n_63710), .D(n_61924), .Z
		(n_1838));
	notech_nand3 i_1936(.A(nbus_11271[3]), .B(nbus_11271[2]), .C(nbus_11271[
		4]), .Z(n_1839));
	notech_and2 i_681(.A(n_1859), .B(n_1860), .Z(n_1844));
	notech_ao3 i_584(.A(n_2968), .B(n_1861), .C(n_28092), .Z(n_1849));
	notech_and4 i_2149(.A(n_63818), .B(\opcode[3] ), .C(n_32697), .D(n_30898
		), .Z(n_1852));
	notech_ao3 i_2137(.A(n_63796), .B(n_63720), .C(n_32390), .Z(n_1854));
	notech_or4 i_1661(.A(n_61748), .B(n_315160779), .C(n_61775), .D(\opcode[3] 
		), .Z(n_1857));
	notech_or4 i_1678(.A(n_32628), .B(n_61748), .C(n_32589), .D(n_60189), .Z
		(n_1858));
	notech_or4 i_1725(.A(n_32391), .B(n_25681), .C(n_63720), .D(n_63762), .Z
		(n_1859));
	notech_or4 i_1732(.A(n_32628), .B(n_25681), .C(n_63700), .D(n_63784), .Z
		(n_1860));
	notech_or4 i_553(.A(n_312460752), .B(n_2952), .C(n_61065), .D(n_2967), .Z
		(n_1861));
	notech_and4 i_1416(.A(n_19672), .B(n_19655), .C(n_30524), .D(n_30324), .Z
		(n_32506));
	notech_and4 i_26884(.A(n_19603), .B(n_30374), .C(n_32521), .D(n_30358), 
		.Z(n_32514));
	notech_nand2 i_2045(.A(n_63818), .B(\opcode[3] ), .Z(n_32383));
	notech_and4 i_827955(.A(n_2922), .B(n_308360711), .C(n_291060622), .D(n_2923
		), .Z(n_32663));
	notech_and4 i_127948(.A(n_2894), .B(n_305960688), .C(n_2882), .D(n_2895)
		, .Z(n_32646));
	notech_and3 i_2157(.A(n_61958), .B(n_63760), .C(n_32388), .Z(n_1855));
	notech_and4 i_51588(.A(fsm[4]), .B(fsm[2]), .C(n_31254), .D(n_61730), .Z
		(n_19629));
	notech_nao3 i_459(.A(n_63818), .B(\opcode[3] ), .C(n_61748), .Z(n_28534)
		);
	notech_or4 i_104037503(.A(n_312460752), .B(n_32383), .C(n_61748), .D(n_2952
		), .Z(n_340661034));
	notech_nand2 i_26914(.A(n_32485), .B(n_61085), .Z(n_32484));
	notech_and2 i_26917(.A(n_19689), .B(n_61110), .Z(n_32481));
	notech_and4 i_51755(.A(fsm[4]), .B(n_31252), .C(fsm[3]), .D(n_61730), .Z
		(n_19595));
	notech_or4 i_53337544(.A(n_63720), .B(n_63784), .C(n_2952), .D(n_30901),
		 .Z(n_340561033));
	notech_nand2 i_137557(.A(n_60440), .B(n_32157), .Z(n_340461032));
	notech_or2 i_037558(.A(n_60440), .B(n_60431), .Z(n_340361031));
	notech_and2 i_51799(.A(n_30842), .B(n_33162), .Z(n_340261030));
	notech_and4 i_51805(.A(n_33163), .B(instrc[94]), .C(n_33155), .D(n_33141
		), .Z(n_340161029));
	notech_and4 i_51806(.A(n_33160), .B(instrc[90]), .C(n_33154), .D(n_33138
		), .Z(n_340061028));
	notech_ao3 i_105937502(.A(n_2850), .B(n_328160909), .C(n_276460613), .Z(n_26398
		));
	notech_or2 i_51752(.A(n_301560644), .B(n_301760646), .Z(n_19612));
	notech_or2 i_169737608(.A(n_19612), .B(n_72012477), .Z(n_71912476));
	notech_nao3 i_54037543(.A(n_312460752), .B(n_61806), .C(n_61739), .Z(n_28007
		));
	notech_or4 i_71837526(.A(n_80512561), .B(all_cnt[2]), .C(n_31370), .D(n_30788
		), .Z(n_30786));
	notech_and2 i_28608(.A(n_57705), .B(n_57686), .Z(n_339961027));
	notech_or4 i_28602(.A(tcmp), .B(n_61815), .C(n_30804), .D(n_336260990), 
		.Z(n_339861026));
	notech_or2 i_205137444(.A(n_61815), .B(tcmp), .Z(n_30800));
	notech_nand2 i_165937620(.A(n_33163), .B(instrc[94]), .Z(n_30815));
	notech_nand2 i_166037621(.A(n_33160), .B(instrc[90]), .Z(n_30822));
	notech_or2 i_71637527(.A(n_75912515), .B(n_32273), .Z(n_30823));
	notech_and4 i_71937525(.A(n_2814), .B(n_30739), .C(all_cnt[1]), .D(n_31371
		), .Z(n_30829));
	notech_and4 i_830574(.A(n_33174), .B(instrc[106]), .C(n_33156), .D(n_33157
		), .Z(n_339761025));
	notech_nand2 i_165837622(.A(n_33174), .B(instrc[106]), .Z(n_30835));
	notech_or4 i_71437528(.A(n_80512561), .B(all_cnt[1]), .C(all_cnt[2]), .D
		(n_340261030), .Z(n_30839));
	notech_ao3 i_137937494(.A(n_33153), .B(instrc[126]), .C(instrc[125]), .Z
		(n_30842));
	notech_or4 i_53437626(.A(n_63720), .B(n_61924), .C(n_61806), .D(n_30901)
		, .Z(n_339661024));
	notech_or2 i_189437461(.A(instrc[112]), .B(n_32158), .Z(n_32217));
	notech_nand2 i_154537483(.A(instrc[112]), .B(instrc[115]), .Z(n_339561023
		));
	notech_nand2 i_864(.A(n_30900), .B(n_312460752), .Z(n_32576));
	notech_or4 i_27082(.A(n_32663), .B(n_309860726), .C(n_61806), .D(n_30901
		), .Z(n_339461022));
	notech_or4 i_52637648(.A(calc_sz[3]), .B(calc_sz[1]), .C(calc_sz[2]), .D
		(n_31373), .Z(n_32319));
	notech_ao3 i_56237540(.A(n_32506), .B(n_32514), .C(n_30336), .Z(n_32353)
		);
	notech_and4 i_148637652(.A(n_61806), .B(n_32663), .C(\opcode[0] ), .D(n_63212389
		), .Z(n_63012387));
	notech_or4 i_1953(.A(n_32576), .B(n_61056), .C(n_32184), .D(n_32628), .Z
		(n_1847));
	notech_or4 i_7537423(.A(tcmp), .B(n_1850), .C(n_61866), .D(n_61614), .Z(n_339361021
		));
	notech_and2 i_4637429(.A(n_322860856), .B(n_322760855), .Z(n_339261020)
		);
	notech_or4 i_67837750(.A(tcmp), .B(n_61815), .C(n_30804), .D(n_57651), .Z
		(n_339161019));
	notech_and4 i_427951(.A(n_290860621), .B(n_307160700), .C(n_2896), .D(n_2909
		), .Z(n_32629));
	notech_and2 i_56837536(.A(n_331860946), .B(n_2817), .Z(n_339061018));
	notech_or4 i_208937785(.A(n_32383), .B(n_61797), .C(n_63784), .D(n_61958
		), .Z(n_338861016));
	notech_nao3 i_31390(.A(n_61775), .B(\opcode[3] ), .C(n_61748), .Z(n_28008
		));
	notech_nand2 i_850(.A(n_30901), .B(n_30900), .Z(n_32589));
	notech_nor2 i_930842(.A(n_32269), .B(instrc[120]), .Z(n_32268));
	notech_ao3 i_930839(.A(n_32161), .B(n_61786), .C(n_58583), .Z(n_32241)
		);
	notech_and4 i_23839(.A(n_61964), .B(n_61828), .C(n_32161), .D(n_61757), 
		.Z(n_32244));
	notech_and4 i_3643341(.A(n_61828), .B(n_32160), .C(n_61766), .D(n_61786)
		, .Z(n_32252));
	notech_and4 i_3943342(.A(n_61964), .B(n_61828), .C(n_61766), .D(n_61786)
		, .Z(n_32259));
	notech_nao3 i_1833(.A(n_61766), .B(n_61964), .C(n_61828), .Z(n_32269));
	notech_nor2 i_4143344(.A(n_32269), .B(n_61757), .Z(n_32263));
	notech_nand2 i_181443275(.A(n_61828), .B(n_32160), .Z(n_338661014));
	notech_ao3 i_4943346(.A(n_61786), .B(instrc[122]), .C(n_58583), .Z(n_32272
		));
	notech_nand3 i_161643279(.A(n_61828), .B(n_61757), .C(n_61944), .Z(n_32305
		));
	notech_and4 i_3243340(.A(n_61828), .B(n_61757), .C(n_61766), .D(n_32160)
		, .Z(n_32247));
	notech_or2 i_1450(.A(n_61828), .B(n_61964), .Z(n_32275));
	notech_and4 i_4243365(.A(n_61828), .B(n_61964), .C(n_61757), .D(n_61944)
		, .Z(n_32304));
	notech_and4 i_3743366(.A(n_61828), .B(n_61786), .C(n_61944), .D(n_61964)
		, .Z(n_32254));
	notech_nao3 i_61246442(.A(n_61928), .B(opa[1]), .C(n_63700), .Z(n_30891)
		);
	notech_or2 i_10279(.A(n_338061008), .B(n_329360921), .Z(n_338561013));
	notech_nao3 i_10278(.A(n_30903), .B(n_32273), .C(n_338061008), .Z(n_338461012
		));
	notech_and4 i_91429156(.A(n_2634), .B(n_2633), .C(n_2629), .D(n_2632), .Z
		(n_338361011));
	notech_and4 i_421762(.A(n_2289), .B(n_2288), .C(n_2283), .D(n_2287), .Z(n_338261010
		));
	notech_and4 i_142649749(.A(n_2272), .B(n_2271), .C(n_2267), .D(n_2270), 
		.Z(n_338161009));
	notech_ao4 i_30737716(.A(n_57672), .B(n_2848), .C(n_32288), .D(n_32215),
		 .Z(n_338061008));
	notech_and4 i_93643348(.A(n_275060599), .B(n_274960598), .C(n_274560594)
		, .D(n_274860597), .Z(n_101026337));
	notech_and4 i_93529168(.A(n_273660587), .B(n_273560586), .C(n_273060582)
		, .D(n_273460585), .Z(n_106826395));
	notech_and4 i_93429167(.A(n_272160573), .B(n_272060572), .C(n_271660568)
		, .D(n_271960571), .Z(n_109226419));
	notech_ao3 i_38349783(.A(n_331660944), .B(n_331760945), .C(n_333660964),
		 .Z(n_122226549));
	notech_and2 i_114049774(.A(n_335460982), .B(n_332960957), .Z(n_122626553
		));
	notech_ao4 i_114149773(.A(n_61841), .B(n_335360981), .C(n_330960937), .D
		(n_323260860), .Z(n_122726554));
	notech_ao3 i_118449756(.A(n_335560983), .B(n_329560923), .C(n_333060958)
		, .Z(n_122826555));
	notech_and3 i_118549755(.A(n_332860956), .B(n_329660924), .C(n_335760985
		), .Z(n_122926556));
	notech_ao3 i_38149785(.A(n_328760915), .B(n_328860916), .C(n_330360931),
		 .Z(n_124126568));
	notech_and2 i_113149781(.A(n_335460982), .B(n_330060928), .Z(n_124526572
		));
	notech_ao4 i_113249780(.A(n_61838), .B(n_335360981), .C(n_328360911), .D
		(n_329060918), .Z(n_124626573));
	notech_ao3 i_117649762(.A(n_328960917), .B(n_335560983), .C(n_329860926)
		, .Z(n_124726574));
	notech_and3 i_117749761(.A(n_329760925), .B(n_329160919), .C(n_335760985
		), .Z(n_124826575));
	notech_ao4 i_23037718(.A(n_61838), .B(n_30341), .C(n_71912476), .D(n_35412112
		), .Z(n_125926586));
	notech_ao4 i_24337719(.A(n_61838), .B(n_30560), .C(n_57001), .D(n_30714)
		, .Z(n_126126588));
	notech_and3 i_38249784(.A(n_331560943), .B(n_275360602), .C(n_26603), .Z
		(n_126226589));
	notech_ao4 i_113349779(.A(n_61838), .B(n_335360981), .C(n_2850), .D(n_329360921
		), .Z(n_126726594));
	notech_and3 i_113449778(.A(n_330160929), .B(n_331260940), .C(n_335460982
		), .Z(n_126826595));
	notech_and3 i_117849760(.A(n_329260920), .B(n_335560983), .C(n_338561013
		), .Z(n_126926596));
	notech_and3 i_117949759(.A(n_329460922), .B(n_335760985), .C(n_338461012
		), .Z(n_127026597));
	notech_or2 i_132749729(.A(n_2034), .B(n_56003), .Z(n_337961007));
	notech_or4 i_41537756(.A(instrc[115]), .B(instrc[112]), .C(n_2829), .D(n_32308
		), .Z(n_337861006));
	notech_nao3 i_32798(.A(n_19612), .B(n_30714), .C(n_57006), .Z(n_26600)
		);
	notech_nao3 i_1949706(.A(n_63770), .B(n_30788), .C(n_2850), .Z(n_337761005
		));
	notech_or4 i_41337546(.A(n_19629), .B(n_57006), .C(n_19612), .D(n_30331)
		, .Z(n_26585));
	notech_nand2 i_1549710(.A(n_203260403), .B(n_27378), .Z(n_337661004));
	notech_nand3 i_2149704(.A(n_63788), .B(n_27378), .C(n_30275), .Z(n_337561003
		));
	notech_nand2 i_132949727(.A(n_203360404), .B(n_28555), .Z(n_337461002)
		);
	notech_nand2 i_21837555(.A(n_61085), .B(n_61614), .Z(n_32196));
	notech_nand3 i_1849707(.A(n_63788), .B(n_28555), .C(n_30906), .Z(n_337361001
		));
	notech_nor2 i_837628(.A(n_340361031), .B(n_2845), .Z(n_32204));
	notech_nor2 i_2850(.A(n_340361031), .B(n_58707), .Z(n_32342));
	notech_nor2 i_3837646(.A(n_60422), .B(n_2821), .Z(n_32311));
	notech_nor2 i_4437630(.A(n_58716), .B(n_2845), .Z(n_32210));
	notech_nor2 i_4537631(.A(n_58716), .B(n_32217), .Z(n_32211));
	notech_nor2 i_2865(.A(n_2830), .B(n_2829), .Z(n_32215));
	notech_nor2 i_5037632(.A(n_340361031), .B(n_32217), .Z(n_32216));
	notech_nor2 i_5137633(.A(n_58716), .B(n_58707), .Z(n_32219));
	notech_and4 i_5337635(.A(n_60440), .B(n_60431), .C(instrc[115]), .D(n_60422
		), .Z(n_32223));
	notech_ao3 i_5437636(.A(instrc[115]), .B(n_60422), .C(n_58716), .Z(n_32224
		));
	notech_ao3 i_5537637(.A(instrc[115]), .B(n_60422), .C(n_340361031), .Z(n_32227
		));
	notech_and4 i_327950(.A(n_2880), .B(n_314660774), .C(n_2868), .D(n_2881)
		, .Z(n_1813));
	notech_nand2 i_1553081(.A(n_63788), .B(opc_10[24]), .Z(n_31942));
	notech_and4 i_144829769(.A(n_197895895), .B(n_197795896), .C(n_197395900
		), .D(n_197695897), .Z(n_363350926));
	notech_and4 i_144629746(.A(n_1994), .B(n_1993), .C(n_198860388), .D(n_1991
		), .Z(n_363450925));
	notech_and4 i_144729757(.A(n_196395907), .B(n_196295908), .C(n_1957), .D
		(n_196195909), .Z(n_364628688));
	notech_and4 i_142949751(.A(n_2244), .B(n_2243), .C(n_2239), .D(n_2242), 
		.Z(n_337261000));
	notech_ao4 i_5555871(.A(n_57566), .B(n_57662), .C(n_30721), .D(n_32220),
		 .Z(n_337160999));
	notech_nor2 i_99455935(.A(n_184660383), .B(n_57512), .Z(n_30725));
	notech_and2 i_97555959(.A(n_60154), .B(n_1862), .Z(n_337060998));
	notech_ao4 i_27955992(.A(n_57672), .B(n_57566), .C(n_57553), .D(n_32220)
		, .Z(n_336860996));
	notech_and4 i_142346451(.A(n_2351), .B(n_2350), .C(n_2346), .D(n_2349), 
		.Z(n_336760995));
	notech_and4 i_143246447(.A(n_2379), .B(n_2378), .C(n_2374), .D(n_2377), 
		.Z(n_336660994));
	notech_and4 i_147937777(.A(n_61806), .B(n_32663), .C(n_61775), .D(n_63212389
		), .Z(n_32368));
	notech_ao4 i_176558172(.A(n_1855), .B(n_30414), .C(n_32317), .D(n_30528)
		, .Z(n_336560993));
	notech_ao3 i_50337649(.A(calc_sz[1]), .B(calc_sz[0]), .C(n_317860806), .Z
		(n_32323));
	notech_nor2 i_830626(.A(n_317960807), .B(n_317860806), .Z(n_32321));
	notech_and2 i_137358180(.A(n_30287), .B(n_1850), .Z(n_336460992));
	notech_or4 i_2140(.A(n_32628), .B(n_61930), .C(n_61958), .D(n_32394), .Z
		(n_1850));
	notech_and2 i_107658190(.A(n_57651), .B(n_57662), .Z(n_336360991));
	notech_and2 i_104837647(.A(n_57672), .B(n_57662), .Z(n_336260990));
	notech_and4 i_142549793(.A(n_2191), .B(n_2190), .C(n_2186), .D(n_2189), 
		.Z(n_336160989));
	notech_and4 i_143049750(.A(n_2258), .B(n_225795868), .C(n_2253), .D(n_225695869
		), .Z(n_336060988));
	notech_nor2 i_51531(.A(n_61885), .B(n_61717), .Z(n_1974696898));
	notech_ao4 i_176760699(.A(n_1854), .B(n_1852), .C(n_32317), .D(n_30528),
		 .Z(n_335960987));
	notech_ao4 i_1163(.A(n_61056), .B(n_32390), .C(n_60189), .D(n_30305), .Z
		(n_32386));
	notech_and3 i_2374(.A(n_57672), .B(n_57662), .C(n_57651), .Z(n_32317));
	notech_or4 i_32160783(.A(n_61864), .B(n_61614), .C(n_1850), .D(n_32317),
		 .Z(n_335760985));
	notech_ao3 i_123060759(.A(n_30287), .B(n_30306), .C(n_1854), .Z(n_335660984
		));
	notech_or4 i_32060784(.A(n_335660984), .B(n_61866), .C(n_61614), .D(n_32317
		), .Z(n_335560983));
	notech_or4 i_31960785(.A(n_61885), .B(n_30694), .C(n_61717), .D(n_61866)
		, .Z(n_335460982));
	notech_nao3 i_21260791(.A(n_57651), .B(n_336260990), .C(n_176660368), .Z
		(n_335360981));
	notech_nao3 i_119346508(.A(n_32249), .B(n_23615), .C(n_365964190), .Z(n_335260980
		));
	notech_nao3 i_119446507(.A(n_23615), .B(n_58561), .C(n_365964190), .Z(n_335160979
		));
	notech_ao3 i_52860721(.A(n_381864349), .B(n_61660), .C(n_26028), .Z(n_335060978
		));
	notech_and4 i_142849752(.A(n_2230), .B(n_2229), .C(n_2225), .D(n_2228), 
		.Z(n_334960977));
	notech_and4 i_91629158(.A(n_266260517), .B(n_266160516), .C(n_265760512)
		, .D(n_266060515), .Z(n_334860976));
	notech_and4 i_142749753(.A(n_2216), .B(n_2215), .C(n_2211), .D(n_2214), 
		.Z(n_334760975));
	notech_and4 i_91529157(.A(n_264860503), .B(n_264760502), .C(n_264360498)
		, .D(n_264660501), .Z(n_334660974));
	notech_ao3 i_930778(.A(n_61766), .B(n_32159), .C(n_58583), .Z(n_32249)
		);
	notech_and3 i_106337760(.A(n_391064441), .B(n_23759), .C(n_23760), .Z(n_334560973
		));
	notech_and2 i_42837730(.A(n_390064431), .B(n_276760616), .Z(n_334460972)
		);
	notech_and4 i_91229154(.A(n_2620), .B(n_2619), .C(n_2615), .D(n_2618), .Z
		(n_334360971));
	notech_nand3 i_70246444(.A(n_63720), .B(n_61930), .C(opb[1]), .Z(n_334260970
		));
	notech_ao3 i_193737618(.A(n_339961027), .B(n_33152), .C(n_57714), .Z(n_30788
		));
	notech_and4 i_142446449(.A(n_2365), .B(n_2364), .C(n_2360), .D(n_2363), 
		.Z(n_334060968));
	notech_and4 i_217568(.A(n_175860360), .B(n_175760359), .C(n_175660358), 
		.D(n_176160363), .Z(n_333960967));
	notech_and4 i_516995(.A(n_174260346), .B(n_174160345), .C(n_174660350), 
		.D(n_174060344), .Z(n_333860966));
	notech_and4 i_616996(.A(n_172260326), .B(n_172160325), .C(n_173260336), 
		.D(n_172060324), .Z(n_333760965));
	notech_nand3 i_41063357(.A(n_176360365), .B(n_61085), .C(n_61660), .Z(n_28240
		));
	notech_and4 i_12185(.A(n_32310), .B(n_61094), .C(n_32321), .D(n_32548), 
		.Z(n_333660964));
	notech_nao3 i_30870(.A(n_171160315), .B(\eflags[10] ), .C(n_61841), .Z(n_333360961
		));
	notech_nao3 i_30868(.A(n_171160315), .B(n_33108), .C(n_61841), .Z(n_333260960
		));
	notech_or4 i_52437778(.A(instrc[115]), .B(n_60422), .C(n_2829), .D(n_32292
		), .Z(n_26603));
	notech_ao4 i_30937610(.A(n_2848), .B(n_57651), .C(n_32292), .D(n_32215),
		 .Z(n_26624));
	notech_ao3 i_194143362(.A(n_61757), .B(n_61944), .C(n_58583), .Z(n_32273
		));
	notech_or4 i_28594(.A(n_61883), .B(n_339461022), .C(n_61717), .D(n_61861
		), .Z(n_30804));
	notech_nor2 i_209163372(.A(n_28558), .B(n_323260860), .Z(n_333060958));
	notech_or4 i_205763374(.A(n_56792), .B(n_2383), .C(n_165695997), .D(n_330960937
		), .Z(n_332960957));
	notech_or4 i_197463375(.A(n_56792), .B(n_2383), .C(n_165695997), .D(n_28558
		), .Z(n_332860956));
	notech_xor2 i_137563378(.A(n_63720), .B(n_61930), .Z(n_332760955));
	notech_or4 i_41263359(.A(n_61880), .B(n_30380), .C(n_61717), .D(n_61861)
		, .Z(n_332660954));
	notech_nao3 i_10068(.A(n_30903), .B(n_32273), .C(n_26624), .Z(n_332560953
		));
	notech_and2 i_125963379(.A(n_332660954), .B(n_332560953), .Z(n_332460952
		));
	notech_or4 i_41163358(.A(n_61880), .B(n_2805), .C(n_61717), .D(n_61864),
		 .Z(n_332360951));
	notech_ao4 i_125863380(.A(n_61838), .B(n_2805), .C(n_26624), .D(n_329360921
		), .Z(n_332260950));
	notech_and2 i_107163388(.A(n_26398), .B(n_338061008), .Z(n_332160949));
	notech_ao4 i_5363304(.A(n_2848), .B(n_57662), .C(n_32290), .D(n_32548), 
		.Z(n_28552));
	notech_ao3 i_1143347(.A(n_61786), .B(n_61944), .C(n_2383), .Z(n_32544)
		);
	notech_ao3 i_137158181(.A(calc_sz[0]), .B(calc_sz[1]), .C(n_317860806), 
		.Z(n_331960947));
	notech_or2 i_56663401(.A(n_331960947), .B(n_176660368), .Z(n_331860946)
		);
	notech_or2 i_50463402(.A(n_32288), .B(n_59095), .Z(n_331760945));
	notech_or2 i_49863403(.A(n_32292), .B(n_59095), .Z(n_331660944));
	notech_or4 i_49937609(.A(instrc[115]), .B(n_60422), .C(n_2829), .D(n_32288
		), .Z(n_331560943));
	notech_and3 i_46263404(.A(n_337861006), .B(n_275360602), .C(n_331560943)
		, .Z(n_331460942));
	notech_nand3 i_24463352(.A(n_184060379), .B(n_61094), .C(n_61660), .Z(n_331360941
		));
	notech_or4 i_205937693(.A(n_61880), .B(n_1847), .C(n_61717), .D(n_61861)
		, .Z(n_331260940));
	notech_and2 i_42463408(.A(n_331360941), .B(n_331260940), .Z(n_331160939)
		);
	notech_or2 i_39463409(.A(n_32308), .B(n_59095), .Z(n_331060938));
	notech_ao4 i_30063411(.A(n_2848), .B(n_57651), .C(n_32292), .D(n_32548),
		 .Z(n_28551));
	notech_ao4 i_29663412(.A(n_2848), .B(n_57637), .C(n_32308), .D(n_32548),
		 .Z(n_330960937));
	notech_ao4 i_29263413(.A(n_57679), .B(n_2848), .C(n_32288), .D(n_32548),
		 .Z(n_28558));
	notech_ao3 i_737627(.A(n_60440), .B(n_60431), .C(n_58707), .Z(n_32203)
		);
	notech_ao3 i_1243339(.A(n_61757), .B(n_61944), .C(n_2383), .Z(n_32243)
		);
	notech_nao3 i_541(.A(n_312460752), .B(n_61806), .C(n_59120), .Z(n_28533)
		);
	notech_or4 i_40666157(.A(n_163296016), .B(n_61861), .C(n_61614), .D(\eflags[10] 
		), .Z(n_330560933));
	notech_or4 i_40566158(.A(n_163296016), .B(n_61861), .C(n_61614), .D(n_33108
		), .Z(n_330460932));
	notech_or4 i_866148(.A(n_2383), .B(n_61786), .C(n_61766), .D(n_163196017
		), .Z(n_27377));
	notech_and4 i_11146(.A(n_32310), .B(n_61094), .C(n_32321), .D(n_57236), 
		.Z(n_330360931));
	notech_or2 i_10284(.A(n_2850), .B(n_329360921), .Z(n_330260930));
	notech_nao3 i_10283(.A(n_30903), .B(n_32273), .C(n_2850), .Z(n_330160929
		));
	notech_nao3 i_208366164(.A(n_32243), .B(n_30275), .C(n_163196017), .Z(n_330060928
		));
	notech_nor2 i_204666166(.A(n_27379), .B(n_329060918), .Z(n_329860926));
	notech_nao3 i_198066168(.A(n_30911), .B(n_32243), .C(n_27379), .Z(n_329760925
		));
	notech_nao3 i_110466180(.A(n_163396015), .B(n_32544), .C(n_165695997), .Z
		(n_329660924));
	notech_nand2 i_110366181(.A(n_163396015), .B(n_30516), .Z(n_329560923)
		);
	notech_nand3 i_109266184(.A(n_30903), .B(n_32273), .C(n_30915), .Z(n_329460922
		));
	notech_and2 i_182437717(.A(n_60154), .B(n_2844), .Z(n_329360921));
	notech_nand2 i_109166185(.A(n_30915), .B(n_30389), .Z(n_329260920));
	notech_nao3 i_109066186(.A(n_220495876), .B(n_32243), .C(n_163196017), .Z
		(n_329160919));
	notech_and2 i_182666169(.A(n_60154), .B(n_164496008), .Z(n_329060918));
	notech_nand2 i_108966187(.A(n_220495876), .B(n_30912), .Z(n_328960917)
		);
	notech_or2 i_50566189(.A(n_32288), .B(n_57225), .Z(n_328860916));
	notech_or2 i_49766190(.A(n_32292), .B(n_57225), .Z(n_328760915));
	notech_or2 i_39566192(.A(n_32308), .B(n_57225), .Z(n_328660914));
	notech_nao3 i_23537781(.A(n_61094), .B(n_32323), .C(n_57566), .Z(n_328560913
		));
	notech_ao4 i_29966193(.A(n_2848), .B(n_57651), .C(n_32292), .D(n_57236),
		 .Z(n_27379));
	notech_ao4 i_29566194(.A(n_2848), .B(n_57637), .C(n_32308), .D(n_57236),
		 .Z(n_328360911));
	notech_ao4 i_29166195(.A(n_57672), .B(n_2848), .C(n_32288), .D(n_57236),
		 .Z(n_83739557));
	notech_or4 i_23837784(.A(calc_sz[3]), .B(calc_sz[2]), .C(n_317960807), .D
		(n_2848), .Z(n_328160909));
	notech_ao4 i_28766196(.A(n_2848), .B(n_57662), .C(n_32290), .D(n_57236),
		 .Z(n_83839558));
	notech_and3 i_11766197(.A(n_57705), .B(n_28557), .C(n_33152), .Z(n_27378
		));
	notech_ao4 i_26955994(.A(n_57566), .B(n_57651), .C(n_30723), .D(n_32220)
		, .Z(n_328060908));
	notech_and4 i_92043354(.A(n_270660559), .B(n_270560558), .C(n_270160554)
		, .D(n_270460557), .Z(n_99942440));
	notech_and4 i_91829159(.A(n_269260545), .B(n_269160544), .C(n_268560540)
		, .D(n_269060543), .Z(n_100242443));
	notech_and4 i_91743356(.A(n_267660531), .B(n_267560530), .C(n_267160526)
		, .D(n_267460529), .Z(n_100542446));
	notech_and4 i_91329155(.A(n_2606), .B(n_2605), .C(n_2601), .D(n_2604), .Z
		(n_100842449));
	notech_and4 i_91129153(.A(n_2592), .B(n_2591), .C(n_2587), .D(n_2590), .Z
		(n_101142452));
	notech_nand2 i_82558196(.A(n_30723), .B(n_30721), .Z(n_115442595));
	notech_or4 i_38855990(.A(n_61815), .B(n_57535), .C(n_57637), .D(n_57163)
		, .Z(n_327960907));
	notech_nand2 i_84158195(.A(n_57553), .B(n_30721), .Z(n_115942600));
	notech_nand3 i_22458211(.A(n_61815), .B(n_32315), .C(n_32323), .Z(n_116342604
		));
	notech_nao3 i_22358212(.A(n_57651), .B(n_336260990), .C(n_57566), .Z(n_116542606
		));
	notech_or4 i_22158214(.A(calc_sz[3]), .B(calc_sz[2]), .C(n_317960807), .D
		(n_57566), .Z(n_116742608));
	notech_and2 i_1038(.A(n_61958), .B(n_63784), .Z(n_32583));
	notech_nand2 i_1046(.A(n_63788), .B(n_63700), .Z(n_32397));
	notech_and3 i_48960678(.A(n_179595933), .B(n_179760373), .C(n_179195937)
		, .Z(n_327860906));
	notech_nand2 i_28627(.A(n_63788), .B(opc_10[0]), .Z(n_327760905));
	notech_nand2 i_28645(.A(n_63788), .B(n_60467), .Z(n_327660904));
	notech_nao3 i_47058137(.A(n_32310), .B(n_32323), .C(n_336760995), .Z(n_327560903
		));
	notech_and3 i_48360684(.A(n_1810), .B(n_1812), .C(n_178695942), .Z(n_327460902
		));
	notech_nao3 i_28077(.A(n_63788), .B(opa[9]), .C(n_63700), .Z(n_327360901
		));
	notech_nand2 i_28080(.A(n_63788), .B(opc_10[9]), .Z(n_327260900));
	notech_nand2 i_28078(.A(n_63788), .B(opc[9]), .Z(n_327160899));
	notech_nao3 i_28100(.A(n_61930), .B(opa[9]), .C(n_63700), .Z(n_327060898
		));
	notech_or2 i_28980(.A(n_336660994), .B(n_57553), .Z(n_326960897));
	notech_and3 i_49660674(.A(n_183160376), .B(n_183660378), .C(n_1771), .Z(n_326860896
		));
	notech_nand3 i_28428(.A(n_63720), .B(n_61930), .C(opb[2]), .Z(n_326760895
		));
	notech_nand3 i_28429(.A(n_63720), .B(n_61930), .C(n_60962), .Z(n_326660894
		));
	notech_nand3 i_28426(.A(n_63720), .B(n_63784), .C(opb[2]), .Z(n_326560893
		));
	notech_nand3 i_28425(.A(n_63720), .B(n_63784), .C(opa[2]), .Z(n_326460892
		));
	notech_nand2 i_28433(.A(n_63744), .B(opc[2]), .Z(n_326360891));
	notech_nand2 i_28432(.A(n_63744), .B(opc_10[2]), .Z(n_326260890));
	notech_nao3 i_34049788(.A(n_61930), .B(opa[2]), .C(n_63700), .Z(n_326160889
		));
	notech_or4 i_50160673(.A(n_61815), .B(n_57535), .C(n_336160989), .D(n_57651
		), .Z(n_326060888));
	notech_nao3 i_34449787(.A(n_63744), .B(opa[2]), .C(n_63700), .Z(n_325960887
		));
	notech_and3 i_49460676(.A(n_182560374), .B(n_183060375), .C(n_177695950)
		, .Z(n_325860886));
	notech_nand3 i_28225(.A(n_63720), .B(n_61930), .C(opb[6]), .Z(n_325760885
		));
	notech_nand3 i_28226(.A(n_63706), .B(n_61930), .C(opa[6]), .Z(n_325660884
		));
	notech_nand3 i_28223(.A(n_63706), .B(n_63760), .C(opb[6]), .Z(n_325560883
		));
	notech_nand3 i_28222(.A(n_63706), .B(n_63760), .C(opa[6]), .Z(n_325460882
		));
	notech_nand2 i_28230(.A(n_63774), .B(opc[6]), .Z(n_325360881));
	notech_nand2 i_28229(.A(n_63774), .B(opc_10[6]), .Z(n_325260880));
	notech_nao3 i_28250(.A(n_61933), .B(opa[6]), .C(n_63712), .Z(n_325160879
		));
	notech_or4 i_29044(.A(n_61815), .B(n_57535), .C(n_337261000), .D(n_57656
		), .Z(n_325060878));
	notech_nao3 i_28249(.A(n_63774), .B(opa[6]), .C(n_63712), .Z(n_324960877
		));
	notech_and3 i_49560675(.A(n_1814), .B(n_1821), .C(n_178195947), .Z(n_324860876
		));
	notech_nand3 i_28165(.A(n_63706), .B(n_63732), .C(opa[7]), .Z(n_324760875
		));
	notech_nand2 i_28177(.A(n_63772), .B(opc_10[7]), .Z(n_324660874));
	notech_nand2 i_28179(.A(n_63792), .B(opc[7]), .Z(n_324560873));
	notech_nand3 i_28171(.A(n_63706), .B(n_61930), .C(opb[7]), .Z(n_324460872
		));
	notech_nand3 i_28168(.A(n_63708), .B(n_63734), .C(opb[7]), .Z(n_324360871
		));
	notech_nand3 i_28173(.A(n_63718), .B(n_61930), .C(opa[7]), .Z(n_324260870
		));
	notech_nao3 i_28199(.A(n_63792), .B(opa[7]), .C(n_63712), .Z(n_324160869
		));
	notech_nao3 i_28200(.A(n_61930), .B(opa[7]), .C(n_63712), .Z(n_324060868
		));
	notech_or2 i_101755936(.A(n_337060998), .B(n_328060908), .Z(n_323960867)
		);
	notech_or4 i_101855976(.A(n_338661014), .B(n_56792), .C(n_184660383), .D
		(n_328060908), .Z(n_323860866));
	notech_or4 i_47560688(.A(n_61815), .B(n_57535), .C(n_336060988), .D(n_57656
		), .Z(n_323760865));
	notech_nor2 i_4337629(.A(n_2829), .B(n_2845), .Z(n_32208));
	notech_ao3 i_5237634(.A(instrc[115]), .B(n_60422), .C(n_2829), .Z(n_32220
		));
	notech_or4 i_21758215(.A(n_339461022), .B(n_61815), .C(n_57672), .D(n_61614
		), .Z(n_30719));
	notech_or4 i_21658142(.A(n_339461022), .B(n_61819), .C(n_61614), .D(n_57656
		), .Z(n_30723));
	notech_or4 i_21458144(.A(n_317960807), .B(n_317860806), .C(n_61819), .D(n_57535
		), .Z(n_30721));
	notech_and2 i_1047(.A(n_61958), .B(n_61930), .Z(n_32697));
	notech_nand2 i_174869261(.A(n_30395), .B(n_57512), .Z(n_30394));
	notech_nand3 i_174769262(.A(n_339961027), .B(n_30727), .C(n_30484), .Z(n_30393
		));
	notech_and4 i_205855964(.A(instrc[118]), .B(n_57714), .C(n_33173), .D(instrc
		[116]), .Z(n_323660864));
	notech_nao3 i_172969264(.A(n_339961027), .B(n_30727), .C(n_303944473), .Z
		(n_30391));
	notech_or4 i_169369270(.A(n_338661014), .B(n_303944473), .C(n_61757), .D
		(n_61766), .Z(n_30390));
	notech_and4 i_4743345(.A(n_61828), .B(n_32160), .C(n_61786), .D(n_61944)
		, .Z(n_32266));
	notech_or4 i_167969271(.A(n_55831), .B(n_303944473), .C(n_338661014), .D
		(n_56792), .Z(n_30387));
	notech_or2 i_167569273(.A(n_303944473), .B(n_32266), .Z(n_30386));
	notech_nor2 i_164269275(.A(n_303844472), .B(n_26957), .Z(n_26822));
	notech_nao3 i_158969278(.A(instrc[116]), .B(n_188662913), .C(n_26951), .Z
		(n_26821));
	notech_ao3 i_158069280(.A(instrc[116]), .B(n_188662913), .C(n_303844472)
		, .Z(n_26823));
	notech_nor2 i_130369287(.A(n_55831), .B(n_303944473), .Z(n_30395));
	notech_or4 i_94969298(.A(n_2577), .B(n_61964), .C(n_1532), .D(n_61766), 
		.Z(n_30002));
	notech_or2 i_94869299(.A(n_1532), .B(n_32261), .Z(n_30001));
	notech_nor2 i_4043343(.A(n_61964), .B(n_32305), .Z(n_32261));
	notech_or4 i_94469300(.A(n_2577), .B(n_61964), .C(n_61766), .D(n_30576),
		 .Z(n_29998));
	notech_nor2 i_13263227(.A(n_30212), .B(n_1532), .Z(n_323560863));
	notech_nand2 i_93869302(.A(n_57500), .B(n_323560863), .Z(n_29997));
	notech_nao3 i_89669303(.A(n_57714), .B(n_275560604), .C(n_1532), .Z(n_29994
		));
	notech_nand3 i_88469304(.A(n_57714), .B(n_275560604), .C(n_30483), .Z(n_29993
		));
	notech_nand2 i_1037(.A(n_61928), .B(n_63712), .Z(n_32401));
	notech_and4 i_196869322(.A(n_57705), .B(n_57714), .C(n_57686), .D(n_33152
		), .Z(n_30212));
	notech_or2 i_147369325(.A(n_288144316), .B(n_26951), .Z(n_26935));
	notech_or4 i_146869326(.A(n_32275), .B(n_56792), .C(n_26951), .D(n_162262654
		), .Z(n_26940));
	notech_and2 i_127169331(.A(n_303544469), .B(n_1492), .Z(n_303144465));
	notech_and2 i_127069332(.A(n_26942), .B(n_303644470), .Z(n_303244466));
	notech_nao3 i_120969335(.A(n_57401), .B(n_30662), .C(n_288444319), .Z(n_303544469
		));
	notech_or4 i_120869336(.A(n_58583), .B(n_56792), .C(n_288444319), .D(n_162262654
		), .Z(n_303644470));
	notech_and2 i_111369338(.A(n_288444319), .B(n_26949), .Z(n_303844472));
	notech_ao4 i_25955970(.A(n_57566), .B(n_57637), .C(n_32220), .D(n_30316)
		, .Z(n_323360861));
	notech_and4 i_107269339(.A(n_57544), .B(n_184360381), .C(n_323360861), .D
		(n_336860996), .Z(n_303944473));
	notech_nor2 i_103969342(.A(n_1481), .B(n_32261), .Z(n_304244476));
	notech_or4 i_87769348(.A(n_61964), .B(n_32305), .C(n_1481), .D(n_305844492
		), .Z(n_30196));
	notech_nor2 i_97469343(.A(n_304244476), .B(n_33214), .Z(n_304344477));
	notech_or2 i_86669350(.A(n_304344477), .B(n_305844492), .Z(n_30191));
	notech_nand3 i_81269354(.A(n_57544), .B(n_1486), .C(n_1484), .Z(n_30077)
		);
	notech_nand2 i_44569356(.A(n_305644490), .B(n_1491), .Z(n_305144485));
	notech_and2 i_43369357(.A(n_305744491), .B(n_1490), .Z(n_305244486));
	notech_and2 i_43269358(.A(n_327960907), .B(n_1489), .Z(n_305344487));
	notech_and3 i_21558143(.A(n_32310), .B(n_57656), .C(n_336260990), .Z(n_30729
		));
	notech_nor2 i_5637638(.A(n_32217), .B(n_2829), .Z(n_125342694));
	notech_or4 i_38969362(.A(n_61819), .B(n_57535), .C(n_57637), .D(n_57112)
		, .Z(n_305744491));
	notech_ao4 i_28069363(.A(n_57672), .B(n_57566), .C(n_57553), .D(n_125342694
		), .Z(n_30201));
	notech_ao4 i_27069365(.A(n_57566), .B(n_57656), .C(n_30723), .D(n_125342694
		), .Z(n_305844492));
	notech_ao4 i_25069368(.A(n_57566), .B(n_57662), .C(n_30721), .D(n_125342694
		), .Z(n_30200));
	notech_and2 i_96963369(.A(n_60154), .B(n_171360317), .Z(n_323260860));
	notech_ao4 i_107837661(.A(n_339061018), .B(n_76712523), .C(n_1460), .D(n_30839
		), .Z(n_323160859));
	notech_ao4 i_110537697(.A(n_1850), .B(n_76712523), .C(n_30823), .D(n_1460
		), .Z(n_111445606));
	notech_or4 i_141737663(.A(n_30786), .B(n_30618), .C(n_30343), .D(n_30550
		), .Z(n_323060858));
	notech_nor2 i_140537749(.A(n_339261020), .B(n_61928), .Z(n_322960857));
	notech_or2 i_28606(.A(n_336260990), .B(n_2810), .Z(n_322860856));
	notech_nao3 i_72937768(.A(n_336260990), .B(n_57656), .C(n_2810), .Z(n_116645658
		));
	notech_or2 i_73137662(.A(n_2810), .B(n_57656), .Z(n_322760855));
	notech_or4 i_96375832(.A(n_61912), .B(n_61898), .C(n_61880), .D(n_61861)
		, .Z(n_32789));
	notech_and2 i_178037694(.A(n_61861), .B(fecx), .Z(n_124545737));
	notech_ao3 i_1037655(.A(n_60440), .B(n_60431), .C(n_2845), .Z(n_32548)
		);
	notech_nand2 i_29128(.A(instrc[96]), .B(n_78412540), .Z(n_322660854));
	notech_and3 i_11863419(.A(n_57705), .B(n_28557), .C(instrc[116]), .Z(n_28555
		));
	notech_nand2 i_140637492(.A(n_57595), .B(n_63734), .Z(n_322560853));
	notech_or4 i_67737619(.A(tcmp), .B(n_61819), .C(n_30804), .D(n_57633), .Z
		(n_30798));
	notech_nand3 i_31266(.A(instrc[125]), .B(n_33153), .C(instrc[126]), .Z(n_322460852
		));
	notech_and2 i_29133(.A(n_63818), .B(instrc[124]), .Z(n_322360851));
	notech_nao3 i_5971905(.A(n_61786), .B(n_61944), .C(n_111445606), .Z(n_30257
		));
	notech_and4 i_72437523(.A(all_cnt[2]), .B(n_30737), .C(all_cnt[1]), .D(n_2814
		), .Z(n_322260850));
	notech_or4 i_29147(.A(n_79512551), .B(all_cnt[0]), .C(all_cnt[3]), .D(n_33143
		), .Z(n_322060848));
	notech_or2 i_3871926(.A(n_323160859), .B(n_33162), .Z(n_30240));
	notech_or4 i_72237524(.A(n_80512561), .B(n_31370), .C(n_31371), .D(n_340161029
		), .Z(n_321960847));
	notech_and2 i_56737537(.A(n_32353), .B(n_32481), .Z(n_30785));
	notech_nor2 i_69937529(.A(n_32484), .B(n_61656), .Z(n_30869));
	notech_nand2 i_1471950(.A(n_323060858), .B(n_30366), .Z(n_241346905));
	notech_nand3 i_971955(.A(n_322860856), .B(n_116645658), .C(n_322760855),
		 .Z(n_241746909));
	notech_nand2 i_2110(.A(n_339861026), .B(n_339161019), .Z(n_321860846));
	notech_nor2 i_371957(.A(n_57595), .B(n_30547), .Z(n_114845640));
	notech_nand2 i_179571969(.A(instrc[104]), .B(instrc[106]), .Z(n_30234)
		);
	notech_nand2 i_177771970(.A(instrc[98]), .B(instrc[97]), .Z(n_30858));
	notech_and4 i_1023(.A(n_321460842), .B(n_321360841), .C(n_301160640), .D
		(n_301360642), .Z(n_321760845));
	notech_ao4 i_1015(.A(n_22752), .B(n_2983), .C(n_57887), .D(n_32496), .Z(n_321460842
		));
	notech_and4 i_101475888(.A(n_321060838), .B(n_300260631), .C(n_300760636
		), .D(n_299960628), .Z(n_321360841));
	notech_ao4 i_996(.A(n_22968), .B(n_32826), .C(n_22967), .D(n_32809), .Z(n_321060838
		));
	notech_and4 i_1019(.A(n_320160829), .B(n_319160819), .C(n_320760835), .D
		(n_300560634), .Z(n_320860836));
	notech_and4 i_1017(.A(n_320460832), .B(n_300160630), .C(n_301060639), .D
		(n_300660635), .Z(n_320760835));
	notech_ao4 i_1000(.A(n_57917), .B(n_58330), .C(n_22977), .D(n_32774), .Z
		(n_320460832));
	notech_and4 i_1008(.A(n_2993), .B(n_319860826), .C(n_299660625), .D(n_300060629
		), .Z(n_320160829));
	notech_and4 i_991(.A(n_319660824), .B(n_2991), .C(n_2992), .D(n_319460822
		), .Z(n_319860826));
	notech_ao4 i_986(.A(n_58492), .B(n_31177), .C(n_31224), .D(n_23359), .Z(n_319660824
		));
	notech_ao3 i_985(.A(n_319260820), .B(n_2988), .C(n_2987), .Z(n_319460822
		));
	notech_ao4 i_982(.A(n_33137), .B(n_57987), .C(n_58007), .D(nbus_11271[5]
		), .Z(n_319260820));
	notech_ao4 i_1011(.A(n_30610), .B(n_32700), .C(n_22985), .D(n_33136), .Z
		(n_319160819));
	notech_and3 i_527(.A(n_58570), .B(n_58561), .C(n_58592), .Z(n_318760815)
		);
	notech_or4 i_65(.A(n_61880), .B(n_58610), .C(n_59120), .D(n_61717), .Z(n_318660814
		));
	notech_nand2 i_27145(.A(n_61766), .B(n_61786), .Z(n_318160809));
	notech_nand2 i_27128(.A(n_61766), .B(n_61964), .Z(n_318060808));
	notech_nand2 i_492(.A(calc_sz[1]), .B(n_31373), .Z(n_317960807));
	notech_or2 i_27071(.A(calc_sz[3]), .B(calc_sz[2]), .Z(n_317860806));
	notech_nand3 i_483(.A(fsm[4]), .B(n_31252), .C(n_31254), .Z(n_317460802)
		);
	notech_and3 i_1991(.A(n_19689), .B(n_61614), .C(n_30324), .Z(n_317260800
		));
	notech_and2 i_444(.A(n_2973), .B(n_1838), .Z(n_316860796));
	notech_or4 i_434(.A(n_312460752), .B(n_32184), .C(n_2970), .D(n_30900), 
		.Z(n_316760795));
	notech_nao3 i_1027(.A(n_31254), .B(n_31252), .C(fsm[4]), .Z(n_316460792)
		);
	notech_nor2 i_108(.A(n_61907), .B(n_61898), .Z(n_316260790));
	notech_nand3 i_1007(.A(fsm[4]), .B(n_31252), .C(fsm[3]), .Z(n_316160789)
		);
	notech_and2 i_92(.A(n_60189), .B(n_60154), .Z(n_315860786));
	notech_ao3 i_1026(.A(n_31252), .B(fsm[3]), .C(fsm[4]), .Z(n_315760785)
		);
	notech_nand2 i_958(.A(n_61907), .B(n_61898), .Z(n_315560783));
	notech_nao3 i_26485(.A(n_312460752), .B(n_61806), .C(n_32627), .Z(n_315460782
		));
	notech_or4 i_356(.A(n_61775), .B(n_61819), .C(n_63712), .D(n_63734), .Z(n_315360781
		));
	notech_or4 i_350(.A(n_312460752), .B(n_61806), .C(n_63712), .D(n_63764),
		 .Z(n_315160779));
	notech_nand2 i_860(.A(n_61806), .B(n_312460752), .Z(n_314960777));
	notech_and4 i_173(.A(n_313860766), .B(n_313760765), .C(n_314460772), .D(n_2879
		), .Z(n_314660774));
	notech_and3 i_171(.A(n_314260770), .B(n_314160769), .C(n_314060768), .Z(n_314460772
		));
	notech_ao4 i_165(.A(n_304260671), .B(n_32117), .C(n_304160670), .D(n_32125
		), .Z(n_314260770));
	notech_ao4 i_164(.A(n_30960), .B(n_32133), .C(n_33178), .D(n_30962), .Z(n_314160769
		));
	notech_ao4 i_168(.A(n_302660655), .B(n_32141), .C(n_302160650), .D(n_32149
		), .Z(n_314060768));
	notech_ao4 i_167(.A(n_303560664), .B(n_32093), .C(n_302860657), .D(n_33179
		), .Z(n_313860766));
	notech_ao4 i_166(.A(n_303760666), .B(n_32101), .C(n_303660665), .D(n_32109
		), .Z(n_313760765));
	notech_and4 i_143(.A(n_312660754), .B(n_312560753), .C(n_313260760), .D(n_2864
		), .Z(n_313460762));
	notech_and3 i_141(.A(n_313060758), .B(n_312960757), .C(n_312860756), .Z(n_313260760
		));
	notech_ao4 i_135(.A(n_304260671), .B(n_32116), .C(n_304160670), .D(n_32124
		), .Z(n_313060758));
	notech_ao4 i_134(.A(n_30960), .B(n_32132), .C(n_33159), .D(n_30962), .Z(n_312960757
		));
	notech_ao4 i_138(.A(n_302660655), .B(n_32140), .C(n_302160650), .D(n_32148
		), .Z(n_312860756));
	notech_ao4 i_137(.A(n_303560664), .B(n_32092), .C(n_302860657), .D(n_33154
		), .Z(n_312660754));
	notech_ao4 i_136(.A(n_303760666), .B(n_32100), .C(n_303660665), .D(n_32108
		), .Z(n_312560753));
	notech_and4 i_527952(.A(n_2965), .B(n_312160749), .C(n_2953), .D(n_2966)
		, .Z(n_312460752));
	notech_and4 i_337(.A(n_311360741), .B(n_311260740), .C(n_311960747), .D(n_2964
		), .Z(n_312160749));
	notech_and3 i_335(.A(n_311760745), .B(n_311660744), .C(n_311560743), .Z(n_311960747
		));
	notech_ao4 i_329(.A(n_32119), .B(n_304260671), .C(n_304160670), .D(n_32127
		), .Z(n_311760745));
	notech_ao4 i_328(.A(n_32135), .B(n_30960), .C(n_33143), .D(n_30962), .Z(n_311660744
		));
	notech_ao4 i_332(.A(n_302660655), .B(n_32143), .C(n_302160650), .D(n_32151
		), .Z(n_311560743));
	notech_ao4 i_331(.A(n_303560664), .B(n_32095), .C(n_302860657), .D(n_33163
		), .Z(n_311360741));
	notech_ao4 i_330(.A(n_303760666), .B(n_32103), .C(n_303660665), .D(n_32111
		), .Z(n_311260740));
	notech_and4 i_310(.A(n_310160729), .B(n_310060728), .C(n_310760735), .D(n_2949
		), .Z(n_310960737));
	notech_and3 i_308(.A(n_310560733), .B(n_310460732), .C(n_310360731), .Z(n_310760735
		));
	notech_ao4 i_302(.A(n_304260671), .B(n_32121), .C(n_304160670), .D(n_32129
		), .Z(n_310560733));
	notech_ao4 i_301(.A(n_30960), .B(n_32137), .C(n_30962), .D(n_33176), .Z(n_310460732
		));
	notech_ao4 i_305(.A(n_302660655), .B(n_32145), .C(n_302160650), .D(n_32153
		), .Z(n_310360731));
	notech_ao4 i_304(.A(n_303560664), .B(n_32097), .C(n_302860657), .D(n_33177
		), .Z(n_310160729));
	notech_ao4 i_303(.A(n_303760666), .B(n_32105), .C(n_303660665), .D(n_32113
		), .Z(n_310060728));
	notech_nand2 i_94775836(.A(n_32663), .B(n_309860726), .Z(n_309960727));
	notech_and4 i_627953(.A(n_2936), .B(n_309560723), .C(n_2924), .D(n_2937)
		, .Z(n_309860726));
	notech_and4 i_284(.A(n_308760715), .B(n_308660714), .C(n_309360721), .D(n_2935
		), .Z(n_309560723));
	notech_and3 i_282(.A(n_309160719), .B(n_309060718), .C(n_308960717), .Z(n_309360721
		));
	notech_ao4 i_276(.A(n_304260671), .B(n_32120), .C(n_304160670), .D(n_32128
		), .Z(n_309160719));
	notech_ao4 i_275(.A(n_30960), .B(n_32136), .C(n_33161), .D(n_30962), .Z(n_309060718
		));
	notech_ao4 i_279(.A(n_302660655), .B(n_32144), .C(n_302160650), .D(n_32152
		), .Z(n_308960717));
	notech_ao4 i_278(.A(n_303560664), .B(n_32096), .C(n_302860657), .D(n_33155
		), .Z(n_308760715));
	notech_ao4 i_277(.A(n_303760666), .B(n_32104), .C(n_303660665), .D(n_32112
		), .Z(n_308660714));
	notech_and4 i_257(.A(n_307560704), .B(n_307460703), .C(n_308160709), .D(n_2921
		), .Z(n_308360711));
	notech_and3 i_255(.A(n_307960707), .B(n_307860706), .C(n_307760705), .Z(n_308160709
		));
	notech_ao4 i_249(.A(n_304260671), .B(n_32122), .C(n_304160670), .D(n_32130
		), .Z(n_307960707));
	notech_ao4 i_248(.A(n_30960), .B(n_32138), .C(n_30962), .D(n_33142), .Z(n_307860706
		));
	notech_ao4 i_252(.A(n_302660655), .B(n_32146), .C(n_302160650), .D(n_32154
		), .Z(n_307760705));
	notech_ao4 i_251(.A(n_303560664), .B(n_32098), .C(n_302860657), .D(n_33141
		), .Z(n_307560704));
	notech_ao4 i_250(.A(n_303760666), .B(n_32106), .C(n_303660665), .D(n_32114
		), .Z(n_307460703));
	notech_and4 i_230(.A(n_306360692), .B(n_306260691), .C(n_306960698), .D(n_2907
		), .Z(n_307160700));
	notech_and3 i_228(.A(n_306760696), .B(n_306660695), .C(n_306560694), .Z(n_306960698
		));
	notech_ao4 i_222(.A(n_304260671), .B(n_32118), .C(n_304160670), .D(n_32126
		), .Z(n_306760696));
	notech_ao4 i_221(.A(n_30960), .B(n_32134), .C(n_30962), .D(n_33139), .Z(n_306660695
		));
	notech_ao4 i_225(.A(n_302660655), .B(n_32142), .C(n_302160650), .D(n_32150
		), .Z(n_306560694));
	notech_ao4 i_224(.A(n_303560664), .B(n_32094), .C(n_302860657), .D(n_33138
		), .Z(n_306360692));
	notech_ao4 i_223(.A(n_303760666), .B(n_32102), .C(n_303660665), .D(n_32110
		), .Z(n_306260691));
	notech_and4 i_201(.A(n_305160680), .B(n_305060679), .C(n_305760686), .D(n_2893
		), .Z(n_305960688));
	notech_and3 i_199(.A(n_305560684), .B(n_305460683), .C(n_305360682), .Z(n_305760686
		));
	notech_ao4 i_193(.A(n_304260671), .B(n_32115), .C(n_304160670), .D(n_32123
		), .Z(n_305560684));
	notech_ao4 i_192(.A(n_30960), .B(n_32131), .C(n_30962), .D(n_33140), .Z(n_305460683
		));
	notech_ao4 i_196(.A(n_302660655), .B(n_32139), .C(n_302160650), .D(n_32147
		), .Z(n_305360682));
	notech_ao4 i_195(.A(n_303560664), .B(n_32091), .C(n_302860657), .D(n_33160
		), .Z(n_305160680));
	notech_ao4 i_194(.A(n_303760666), .B(n_32099), .C(n_303660665), .D(n_32107
		), .Z(n_305060679));
	notech_ao3 i_43(.A(n_304460673), .B(n_304660675), .C(n_304560674), .Z(n_304860677
		));
	notech_nand3 i_1282679(.A(vliw_pc[2]), .B(n_302460653), .C(n_1816), .Z(n_304660675
		));
	notech_ao3 i_51543(.A(vliw_pc[0]), .B(n_304060669), .C(vliw_pc[1]), .Z(n_304560674
		));
	notech_and4 i_1288(.A(n_303760666), .B(n_303660665), .C(n_303560664), .D
		(n_304360672), .Z(n_304460673));
	notech_and2 i_20(.A(n_304260671), .B(n_304160670), .Z(n_304360672));
	notech_nao3 i_51546(.A(n_32779), .B(n_302460653), .C(vliw_pc[2]), .Z(n_304260671
		));
	notech_nand3 i_51545(.A(vliw_pc[2]), .B(n_302460653), .C(n_302560654), .Z
		(n_304160670));
	notech_and3 i_1024(.A(vliw_pc[2]), .B(n_31258), .C(n_31257), .Z(n_304060669
		));
	notech_or4 i_51549(.A(vliw_pc[2]), .B(vliw_pc[1]), .C(n_31256), .D(n_30963
		), .Z(n_303760666));
	notech_or4 i_51548(.A(vliw_pc[2]), .B(vliw_pc[4]), .C(vliw_pc[3]), .D(n_30653
		), .Z(n_303660665));
	notech_or4 i_51551(.A(vliw_pc[2]), .B(vliw_pc[4]), .C(vliw_pc[3]), .D(n_30964
		), .Z(n_303560664));
	notech_and4 i_51533(.A(vliw_pc[2]), .B(n_31258), .C(vliw_pc[3]), .D(n_302560654
		), .Z(n_303260661));
	notech_and4 i_1870(.A(n_302760656), .B(n_302260651), .C(n_302160650), .D
		(n_302860657), .Z(n_303060659));
	notech_nao3 i_51534(.A(vliw_pc[1]), .B(vliw_pc[0]), .C(n_302060649), .Z(n_302860657
		));
	notech_ao4 i_1459(.A(n_30964), .B(n_302060649), .C(vliw_pc[4]), .D(vliw_pc
		[3]), .Z(n_302760656));
	notech_or4 i_51539(.A(vliw_pc[1]), .B(vliw_pc[0]), .C(vliw_pc[2]), .D(n_32756
		), .Z(n_302660655));
	notech_nor2 i_995(.A(vliw_pc[1]), .B(vliw_pc[0]), .Z(n_302560654));
	notech_and2 i_885(.A(n_31258), .B(n_31257), .Z(n_302460653));
	notech_or4 i_1182677(.A(vliw_pc[2]), .B(vliw_pc[4]), .C(n_31257), .D(n_30653
		), .Z(n_302260651));
	notech_or4 i_51537(.A(vliw_pc[1]), .B(vliw_pc[2]), .C(n_32756), .D(n_31256
		), .Z(n_302160650));
	notech_nao3 i_1002(.A(n_31258), .B(vliw_pc[3]), .C(vliw_pc[2]), .Z(n_302060649
		));
	notech_nao3 i_1028(.A(n_31254), .B(fsm[2]), .C(fsm[4]), .Z(n_301960648)
		);
	notech_nand3 i_990(.A(fsm[4]), .B(fsm[2]), .C(n_31254), .Z(n_301760646)
		);
	notech_nand2 i_962(.A(n_61907), .B(n_31251), .Z(n_301560644));
	notech_nand3 i_617732(.A(n_320860836), .B(n_321760845), .C(n_301260641),
		 .Z(n_301460643));
	notech_or2 i_981(.A(n_2984), .B(nbus_11273[5]), .Z(n_301360642));
	notech_or2 i_971(.A(n_57867), .B(n_33135), .Z(n_301260641));
	notech_nand2 i_972(.A(resa_shiftbox[5]), .B(n_30273), .Z(n_301160640));
	notech_or2 i_952(.A(n_58512), .B(\nbus_11290[5] ), .Z(n_301060639));
	notech_nand3 i_94575884(.A(mul64[5]), .B(n_30648), .C(n_61656), .Z(n_300760636
		));
	notech_nao3 i_969(.A(nbus_134[5]), .B(n_61660), .C(n_1799), .Z(n_300660635
		));
	notech_nao3 i_96775886(.A(opa_0[5]), .B(n_61660), .C(n_1803), .Z(n_300560634
		));
	notech_or2 i_970(.A(n_22742), .B(n_56983), .Z(n_300260631));
	notech_nao3 i_960(.A(nbus_140[5]), .B(n_61660), .C(n_1801), .Z(n_300160630
		));
	notech_or4 i_977(.A(n_60189), .B(n_25485), .C(n_61616), .D(n_58965), .Z(n_300060629
		));
	notech_nao3 i_946(.A(resa_arithbox[5]), .B(n_61660), .C(n_27914), .Z(n_299960628
		));
	notech_nao3 i_96475885(.A(nbus_138[5]), .B(n_61660), .C(n_1802), .Z(n_299660625
		));
	notech_or2 i_965(.A(n_22979), .B(n_58884), .Z(n_2993));
	notech_or2 i_974(.A(n_57998), .B(n_32033), .Z(n_2992));
	notech_nand2 i_951(.A(\nbus_14542[5] ), .B(n_23351), .Z(n_2991));
	notech_nao3 i_948(.A(cr2_reg[5]), .B(n_58601), .C(n_58501), .Z(n_2988)
		);
	notech_and4 i_956(.A(resa_shift4box[5]), .B(n_27823), .C(n_30364), .D(n_317260800
		), .Z(n_2987));
	notech_ao4 i_943(.A(n_57896), .B(nbus_11291[5]), .C(n_2974), .D(n_61616)
		, .Z(n_2984));
	notech_xor2 i_938(.A(n_27831), .B(opa[5]), .Z(n_2983));
	notech_and4 i_445(.A(n_1820), .B(n_316860796), .C(n_58541), .D(n_25468),
		 .Z(n_2974));
	notech_or4 i_1708(.A(n_32589), .B(n_61739), .C(n_63712), .D(n_61928), .Z
		(n_2973));
	notech_and2 i_431(.A(n_63800), .B(n_60154), .Z(n_2970));
	notech_or4 i_362(.A(n_312460752), .B(n_61806), .C(n_61065), .D(n_315860786
		), .Z(n_2968));
	notech_and2 i_340(.A(n_61056), .B(n_60169), .Z(n_2967));
	notech_nand3 i_315(.A(n_304860677), .B(instrc[60]), .C(n_302460653), .Z(n_2966
		));
	notech_or2 i_326(.A(n_302260651), .B(n_33149), .Z(n_2965));
	notech_nand3 i_327(.A(instrc[52]), .B(n_304060669), .C(n_1816), .Z(n_2964
		));
	notech_nao3 i_314(.A(n_303060659), .B(instrc[124]), .C(n_303260661), .Z(n_2953
		));
	notech_and4 i_727954(.A(n_2950), .B(n_310960737), .C(n_2938), .D(n_2951)
		, .Z(n_2952));
	notech_nand3 i_288(.A(n_302460653), .B(n_304860677), .C(instrc[62]), .Z(n_2951
		));
	notech_or2 i_299(.A(n_302260651), .B(n_33148), .Z(n_2950));
	notech_nand3 i_300(.A(n_304060669), .B(n_1816), .C(instrc[54]), .Z(n_2949
		));
	notech_nao3 i_287(.A(n_303060659), .B(instrc[126]), .C(n_303260661), .Z(n_2938
		));
	notech_nand3 i_262(.A(n_302460653), .B(n_304860677), .C(instrc[61]), .Z(n_2937
		));
	notech_or2 i_273(.A(n_302260651), .B(n_33147), .Z(n_2936));
	notech_nand3 i_274(.A(n_304060669), .B(n_1816), .C(instrc[53]), .Z(n_2935
		));
	notech_ao4 i_575812(.A(n_33179), .B(n_91093393), .C(n_33154), .D(n_163094113
		), .Z(n_90793390));
	notech_and2 i_375814(.A(instrc[89]), .B(n_30743), .Z(n_91093393));
	notech_ao4 i_475813(.A(n_33177), .B(n_91593398), .C(n_33155), .D(n_156594048
		), .Z(n_91293395));
	notech_and2 i_275815(.A(n_156594048), .B(instrc[93]), .Z(n_91593398));
	notech_nao3 i_53075289(.A(n_375664287), .B(instrc[107]), .C(n_148993972)
		, .Z(n_91693399));
	notech_and2 i_26975550(.A(n_30822), .B(n_30922), .Z(n_104593528));
	notech_and2 i_39875421(.A(n_30815), .B(n_30921), .Z(n_117493657));
	notech_and2 i_53175288(.A(n_30835), .B(n_30234), .Z(n_130393786));
	notech_ao4 i_99974830(.A(n_20898), .B(n_31611), .C(n_31261), .D(n_20897)
		, .Z(n_142693909));
	notech_ao4 i_99874831(.A(n_56003), .B(n_30967), .C(n_30753), .D(n_31294)
		, .Z(n_142793910));
	notech_ao4 i_99774832(.A(n_20898), .B(n_31612), .C(n_20897), .D(n_31262)
		, .Z(n_142893911));
	notech_ao4 i_99674833(.A(n_56003), .B(n_30969), .C(n_30753), .D(n_31295)
		, .Z(n_142993912));
	notech_ao4 i_99574834(.A(n_20898), .B(n_31613), .C(n_20897), .D(n_31263)
		, .Z(n_143093913));
	notech_ao4 i_99474835(.A(n_56003), .B(n_30971), .C(n_30753), .D(n_31296)
		, .Z(n_143193914));
	notech_ao4 i_99374836(.A(n_20898), .B(n_31614), .C(n_20897), .D(n_31264)
		, .Z(n_143293915));
	notech_ao4 i_99274837(.A(n_56003), .B(n_30973), .C(n_30753), .D(n_31297)
		, .Z(n_143393916));
	notech_ao4 i_98974840(.A(n_20898), .B(n_31616), .C(n_20897), .D(n_31266)
		, .Z(n_143493917));
	notech_ao4 i_98874841(.A(n_56003), .B(n_30977), .C(n_30753), .D(n_31299)
		, .Z(n_143593918));
	notech_ao4 i_98774842(.A(n_20898), .B(n_31617), .C(n_20897), .D(n_31267)
		, .Z(n_143693919));
	notech_ao4 i_98674843(.A(n_56003), .B(n_30979), .C(n_30753), .D(n_31300)
		, .Z(n_143793920));
	notech_ao4 i_98574844(.A(n_20898), .B(n_31618), .C(n_20897), .D(n_31268)
		, .Z(n_143893921));
	notech_ao4 i_98474845(.A(n_56003), .B(n_30981), .C(n_30753), .D(n_31301)
		, .Z(n_143993922));
	notech_ao4 i_98374846(.A(n_20898), .B(n_31619), .C(n_20897), .D(n_31269)
		, .Z(n_144093923));
	notech_ao4 i_98274847(.A(n_56003), .B(n_30983), .C(n_30753), .D(n_31302)
		, .Z(n_144193924));
	notech_ao4 i_98174848(.A(n_20898), .B(n_31620), .C(n_20897), .D(n_31270)
		, .Z(n_144293925));
	notech_ao4 i_98074849(.A(n_56003), .B(n_30985), .C(n_30753), .D(n_31303)
		, .Z(n_144393926));
	notech_ao4 i_97974850(.A(n_20898), .B(n_31621), .C(n_20897), .D(n_31271)
		, .Z(n_144493927));
	notech_ao4 i_97874851(.A(n_56003), .B(n_30987), .C(n_30753), .D(n_31304)
		, .Z(n_144593928));
	notech_ao4 i_97774852(.A(n_20898), .B(n_31622), .C(n_20897), .D(n_31272)
		, .Z(n_144693929));
	notech_ao4 i_97674853(.A(n_56002), .B(n_30989), .C(n_30753), .D(n_31305)
		, .Z(n_144793930));
	notech_ao4 i_97574854(.A(n_20898), .B(n_31623), .C(n_20897), .D(n_31273)
		, .Z(n_144893931));
	notech_ao4 i_97474855(.A(n_55997), .B(n_30991), .C(n_30753), .D(n_31306)
		, .Z(n_144993932));
	notech_ao4 i_97374856(.A(n_20898), .B(n_31624), .C(n_20897), .D(n_31274)
		, .Z(n_145093933));
	notech_ao4 i_97274857(.A(n_55997), .B(n_30993), .C(n_30753), .D(n_31307)
		, .Z(n_145193934));
	notech_ao4 i_97174858(.A(n_20898), .B(n_31625), .C(n_20897), .D(n_31275)
		, .Z(n_145293935));
	notech_ao4 i_97074859(.A(n_55997), .B(n_30995), .C(n_30753), .D(n_31308)
		, .Z(n_145393936));
	notech_ao4 i_96974860(.A(n_20898), .B(n_31626), .C(n_20897), .D(n_31276)
		, .Z(n_145493937));
	notech_ao4 i_96874861(.A(n_55997), .B(n_30997), .C(n_30753), .D(n_31309)
		, .Z(n_145593938));
	notech_ao4 i_96774862(.A(n_55187), .B(n_31627), .C(n_55178), .D(n_31277)
		, .Z(n_145693939));
	notech_ao4 i_96674863(.A(n_55997), .B(n_30999), .C(n_55198), .D(n_31310)
		, .Z(n_145793940));
	notech_ao4 i_96574864(.A(n_55187), .B(n_31629), .C(n_55178), .D(n_31279)
		, .Z(n_145893941));
	notech_ao4 i_96474865(.A(n_55997), .B(n_31004), .C(n_55198), .D(n_31312)
		, .Z(n_145993942));
	notech_ao4 i_96374866(.A(n_55187), .B(n_31630), .C(n_55178), .D(n_31280)
		, .Z(n_146093943));
	notech_ao4 i_96274867(.A(n_55997), .B(n_31006), .C(n_55198), .D(n_31313)
		, .Z(n_146193944));
	notech_ao4 i_96174868(.A(n_55187), .B(n_31631), .C(n_55178), .D(n_31281)
		, .Z(n_146293945));
	notech_ao4 i_96074869(.A(n_55997), .B(n_31008), .C(n_55198), .D(n_31314)
		, .Z(n_146393946));
	notech_ao4 i_95974870(.A(n_55187), .B(n_31632), .C(n_55178), .D(n_31282)
		, .Z(n_146493947));
	notech_ao4 i_95874871(.A(n_55997), .B(n_31010), .C(n_55198), .D(n_31315)
		, .Z(n_146593948));
	notech_ao4 i_95774872(.A(n_55187), .B(n_31633), .C(n_55178), .D(n_31283)
		, .Z(n_146693949));
	notech_ao4 i_95574873(.A(n_55997), .B(n_31012), .C(n_55198), .D(n_31316)
		, .Z(n_146793950));
	notech_ao4 i_95474874(.A(n_55187), .B(n_31634), .C(n_55178), .D(n_31284)
		, .Z(n_146893951));
	notech_ao4 i_95374875(.A(n_55997), .B(n_31014), .C(n_55198), .D(n_31317)
		, .Z(n_146993952));
	notech_ao4 i_95274876(.A(n_55187), .B(n_31635), .C(n_55178), .D(n_31285)
		, .Z(n_147093953));
	notech_ao4 i_95174877(.A(n_56002), .B(n_31016), .C(n_31318), .D(n_55198)
		, .Z(n_147193954));
	notech_ao4 i_95074878(.A(n_55187), .B(n_31636), .C(n_55178), .D(n_31286)
		, .Z(n_147293955));
	notech_ao4 i_94974879(.A(n_56002), .B(n_31018), .C(n_55198), .D(n_31319)
		, .Z(n_147393956));
	notech_ao4 i_94874880(.A(n_55187), .B(n_31637), .C(n_55178), .D(n_31287)
		, .Z(n_147493957));
	notech_ao4 i_94774881(.A(n_56002), .B(n_31020), .C(n_55198), .D(n_31320)
		, .Z(n_147593958));
	notech_ao4 i_94674882(.A(n_55187), .B(n_31638), .C(n_20897), .D(n_31288)
		, .Z(n_147693959));
	notech_ao4 i_94574883(.A(n_56002), .B(n_31022), .C(n_30753), .D(n_31321)
		, .Z(n_147793960));
	notech_ao4 i_94474884(.A(n_55187), .B(n_31639), .C(n_55178), .D(n_31289)
		, .Z(n_147893961));
	notech_ao4 i_94374885(.A(n_56002), .B(n_31024), .C(n_55198), .D(n_31322)
		, .Z(n_147993962));
	notech_ao4 i_94274886(.A(n_55187), .B(n_31640), .C(n_55178), .D(n_31290)
		, .Z(n_148093963));
	notech_ao4 i_94174887(.A(n_56002), .B(n_31026), .C(n_55198), .D(n_31323)
		, .Z(n_148193964));
	notech_ao4 i_94074888(.A(n_55187), .B(n_31641), .C(n_55178), .D(n_31291)
		, .Z(n_148293965));
	notech_ao4 i_93974889(.A(n_56002), .B(n_31028), .C(n_55198), .D(n_31324)
		, .Z(n_148393966));
	notech_ao4 i_93874890(.A(n_55187), .B(n_31642), .C(n_55178), .D(n_31292)
		, .Z(n_148493967));
	notech_ao4 i_93774891(.A(n_56002), .B(n_31030), .C(n_55198), .D(n_31325)
		, .Z(n_148593968));
	notech_or4 i_65975820(.A(instrc[104]), .B(instrc[106]), .C(n_33156), .D(n_33157
		), .Z(n_148793970));
	notech_mux2 i_93474894(.S(instrc[105]), .A(n_33164), .B(n_29232), .Z(n_148993972
		));
	notech_nand2 i_65575823(.A(n_30739), .B(n_91693399), .Z(n_149093973));
	notech_ao4 i_93174897(.A(n_149093973), .B(n_33925), .C(n_31261), .D(n_148793970
		), .Z(n_149193974));
	notech_or4 i_65475824(.A(n_33157), .B(instrc[105]), .C(n_130393786), .D(n_339761025
		), .Z(n_149493977));
	notech_ao4 i_93074898(.A(n_30739), .B(n_30967), .C(n_31294), .D(n_149493977
		), .Z(n_149593978));
	notech_ao4 i_92974899(.A(n_149093973), .B(n_33924), .C(n_31262), .D(n_148793970
		), .Z(n_149693979));
	notech_ao4 i_92874900(.A(n_30739), .B(n_30969), .C(n_31295), .D(n_149493977
		), .Z(n_149793980));
	notech_ao4 i_92774901(.A(n_149093973), .B(n_33923), .C(n_31263), .D(n_148793970
		), .Z(n_149893981));
	notech_ao4 i_92674902(.A(n_30739), .B(n_30971), .C(n_31296), .D(n_149493977
		), .Z(n_149993982));
	notech_ao4 i_92574903(.A(n_149093973), .B(n_33922), .C(n_31264), .D(n_148793970
		), .Z(n_150093983));
	notech_ao4 i_92474904(.A(n_30739), .B(n_30973), .C(n_31297), .D(n_149493977
		), .Z(n_150193984));
	notech_ao4 i_92374905(.A(n_149093973), .B(n_33921), .C(n_31265), .D(n_148793970
		), .Z(n_150293985));
	notech_ao4 i_92274906(.A(n_30739), .B(n_30975), .C(n_31298), .D(n_149493977
		), .Z(n_150393986));
	notech_ao4 i_92174907(.A(n_149093973), .B(n_33920), .C(n_31266), .D(n_148793970
		), .Z(n_150493987));
	notech_ao4 i_92074908(.A(n_30739), .B(n_30977), .C(n_31299), .D(n_149493977
		), .Z(n_150593988));
	notech_ao4 i_91974909(.A(n_149093973), .B(n_33919), .C(n_31267), .D(n_148793970
		), .Z(n_150693989));
	notech_ao4 i_91874910(.A(n_30739), .B(n_30979), .C(n_31300), .D(n_149493977
		), .Z(n_150793990));
	notech_ao4 i_91774911(.A(n_149093973), .B(n_33918), .C(n_31268), .D(n_148793970
		), .Z(n_150893991));
	notech_ao4 i_91674912(.A(n_30739), .B(n_30981), .C(n_31301), .D(n_149493977
		), .Z(n_150993992));
	notech_ao4 i_91574913(.A(n_149093973), .B(n_33917), .C(n_31269), .D(n_148793970
		), .Z(n_151093993));
	notech_ao4 i_91474914(.A(n_30739), .B(n_30983), .C(n_31302), .D(n_149493977
		), .Z(n_151193994));
	notech_ao4 i_91374915(.A(n_149093973), .B(n_33916), .C(n_31270), .D(n_148793970
		), .Z(n_151293995));
	notech_ao4 i_91274916(.A(n_30739), .B(n_30985), .C(n_31303), .D(n_149493977
		), .Z(n_151393996));
	notech_ao4 i_91174917(.A(n_149093973), .B(n_33915), .C(n_31271), .D(n_148793970
		), .Z(n_151493997));
	notech_ao4 i_91074918(.A(n_30739), .B(n_30987), .C(n_31304), .D(n_149493977
		), .Z(n_151593998));
	notech_ao4 i_90974919(.A(n_149093973), .B(n_33914), .C(n_31272), .D(n_148793970
		), .Z(n_151693999));
	notech_ao4 i_90874920(.A(n_30739), .B(n_30989), .C(n_31305), .D(n_149493977
		), .Z(n_151794000));
	notech_ao4 i_90774921(.A(n_149093973), .B(n_33913), .C(n_31273), .D(n_148793970
		), .Z(n_151894001));
	notech_ao4 i_90674922(.A(n_30739), .B(n_30991), .C(n_31306), .D(n_149493977
		), .Z(n_151994002));
	notech_ao4 i_90574923(.A(n_149093973), .B(n_33912), .C(n_31274), .D(n_148793970
		), .Z(n_152094003));
	notech_ao4 i_90474924(.A(n_30739), .B(n_30993), .C(n_31307), .D(n_149493977
		), .Z(n_152194004));
	notech_ao4 i_90374925(.A(n_149093973), .B(n_33911), .C(n_31275), .D(n_148793970
		), .Z(n_152294005));
	notech_ao4 i_90274926(.A(n_30739), .B(n_30995), .C(n_31308), .D(n_149493977
		), .Z(n_152394006));
	notech_ao4 i_90174927(.A(n_149093973), .B(n_33910), .C(n_31276), .D(n_148793970
		), .Z(n_152494007));
	notech_ao4 i_90074928(.A(n_57586), .B(n_30997), .C(n_31309), .D(n_149493977
		), .Z(n_152594008));
	notech_ao4 i_89974929(.A(n_55158), .B(n_33909), .C(n_31277), .D(n_55039)
		, .Z(n_152694009));
	notech_ao4 i_89874930(.A(n_57586), .B(n_30999), .C(n_31310), .D(n_55169)
		, .Z(n_152794010));
	notech_ao4 i_89774931(.A(n_55158), .B(n_33908), .C(n_31278), .D(n_55039)
		, .Z(n_152894011));
	notech_ao4 i_89674932(.A(n_57586), .B(n_31002), .C(n_31311), .D(n_55169)
		, .Z(n_152994012));
	notech_ao4 i_89574933(.A(n_55158), .B(n_33907), .C(n_31279), .D(n_55039)
		, .Z(n_153094013));
	notech_ao4 i_89474934(.A(n_57586), .B(n_31004), .C(n_31312), .D(n_55169)
		, .Z(n_153194014));
	notech_ao4 i_89374935(.A(n_55158), .B(n_33906), .C(n_31280), .D(n_55039)
		, .Z(n_153294015));
	notech_ao4 i_89274936(.A(n_57586), .B(n_31006), .C(n_31313), .D(n_55169)
		, .Z(n_153394016));
	notech_ao4 i_89174937(.A(n_55158), .B(n_33905), .C(n_31281), .D(n_55039)
		, .Z(n_153494017));
	notech_ao4 i_89074938(.A(n_57586), .B(n_31008), .C(n_31314), .D(n_55169)
		, .Z(n_153594018));
	notech_ao4 i_88974939(.A(n_55158), .B(n_33904), .C(n_31282), .D(n_55039)
		, .Z(n_153694019));
	notech_ao4 i_88874940(.A(n_57586), .B(n_31010), .C(n_31315), .D(n_55169)
		, .Z(n_153794020));
	notech_ao4 i_88774941(.A(n_55158), .B(n_33903), .C(n_31283), .D(n_55039)
		, .Z(n_153894021));
	notech_ao4 i_88674942(.A(n_57586), .B(n_31012), .C(n_31316), .D(n_55169)
		, .Z(n_153994022));
	notech_ao4 i_88574943(.A(n_55158), .B(n_33902), .C(n_31284), .D(n_55039)
		, .Z(n_154094023));
	notech_ao4 i_88474944(.A(n_57586), .B(n_31014), .C(n_31317), .D(n_55169)
		, .Z(n_154194024));
	notech_ao4 i_88374945(.A(n_55158), .B(n_33901), .C(n_31285), .D(n_55039)
		, .Z(n_154294025));
	notech_ao4 i_88274946(.A(n_57586), .B(n_31016), .C(n_31318), .D(n_55169)
		, .Z(n_154394026));
	notech_ao4 i_88174947(.A(n_55158), .B(n_33900), .C(n_31286), .D(n_55039)
		, .Z(n_154494027));
	notech_ao4 i_88074948(.A(n_57586), .B(n_31018), .C(n_31319), .D(n_55169)
		, .Z(n_154594028));
	notech_ao4 i_87974949(.A(n_55158), .B(n_33899), .C(n_31287), .D(n_148793970
		), .Z(n_154694029));
	notech_ao4 i_87874950(.A(n_57586), .B(n_31020), .C(n_31320), .D(n_149493977
		), .Z(n_154794030));
	notech_ao4 i_87774951(.A(n_55158), .B(n_33898), .C(n_31288), .D(n_55039)
		, .Z(n_154894031));
	notech_ao4 i_87674952(.A(n_57586), .B(n_31022), .C(n_31321), .D(n_55169)
		, .Z(n_154994032));
	notech_ao4 i_87574953(.A(n_55158), .B(n_33897), .C(n_31289), .D(n_55039)
		, .Z(n_155094033));
	notech_ao4 i_87474954(.A(n_57586), .B(n_31024), .C(n_31322), .D(n_55169)
		, .Z(n_155194034));
	notech_ao4 i_87374955(.A(n_55158), .B(n_33896), .C(n_31290), .D(n_55039)
		, .Z(n_155294035));
	notech_ao4 i_87274956(.A(n_57586), .B(n_31026), .C(n_31323), .D(n_55169)
		, .Z(n_155394036));
	notech_ao4 i_87174957(.A(n_55158), .B(n_33895), .C(n_31291), .D(n_55039)
		, .Z(n_155494037));
	notech_ao4 i_87074958(.A(n_57586), .B(n_31028), .C(n_31324), .D(n_55169)
		, .Z(n_155594038));
	notech_ao4 i_86974959(.A(n_55158), .B(n_33894), .C(n_31292), .D(n_55039)
		, .Z(n_155694039));
	notech_ao4 i_86874960(.A(n_57586), .B(n_31030), .C(n_31325), .D(n_55169)
		, .Z(n_155794040));
	notech_or4 i_66975818(.A(instrc[93]), .B(n_340161029), .C(n_33141), .D(n_117493657
		), .Z(n_156094043));
	notech_or4 i_65775821(.A(n_156594048), .B(n_33141), .C(n_340161029), .D(n_33155
		), .Z(n_156394046));
	notech_ao4 i_86274966(.A(n_31261), .B(n_156394046), .C(n_31294), .D(n_156094043
		), .Z(n_156494047));
	notech_nand2 i_86374965(.A(n_33163), .B(n_33177), .Z(n_156594048));
	notech_ao4 i_64675826(.A(n_30815), .B(n_77812534), .C(n_91293395), .D(n_33141
		), .Z(n_156694049));
	notech_ao4 i_86174967(.A(n_30738), .B(n_30967), .C(n_30741), .D(n_33893)
		, .Z(n_156794050));
	notech_ao4 i_86074968(.A(n_31262), .B(n_156394046), .C(n_31295), .D(n_156094043
		), .Z(n_156894051));
	notech_ao4 i_85974969(.A(n_30738), .B(n_30969), .C(n_30741), .D(n_33892)
		, .Z(n_156994052));
	notech_ao4 i_85874970(.A(n_31263), .B(n_156394046), .C(n_156094043), .D(n_31296
		), .Z(n_157094053));
	notech_ao4 i_85774971(.A(n_30738), .B(n_30971), .C(n_30741), .D(n_33891)
		, .Z(n_157194054));
	notech_ao4 i_85674972(.A(n_31264), .B(n_156394046), .C(n_31297), .D(n_156094043
		), .Z(n_157294055));
	notech_ao4 i_85574973(.A(n_30738), .B(n_30973), .C(n_30741), .D(n_33890)
		, .Z(n_157394056));
	notech_ao4 i_85474974(.A(n_31265), .B(n_156394046), .C(n_156094043), .D(n_31298
		), .Z(n_157494057));
	notech_ao4 i_85374975(.A(n_30738), .B(n_30975), .C(n_30741), .D(n_33889)
		, .Z(n_157594058));
	notech_ao4 i_85274976(.A(n_31266), .B(n_156394046), .C(n_156094043), .D(n_31299
		), .Z(n_157694059));
	notech_ao4 i_85174977(.A(n_30738), .B(n_30977), .C(n_30741), .D(n_33888)
		, .Z(n_157794060));
	notech_ao4 i_85074978(.A(n_31267), .B(n_156394046), .C(n_156094043), .D(n_31300
		), .Z(n_157894061));
	notech_ao4 i_84974979(.A(n_30738), .B(n_30979), .C(n_30741), .D(n_33887)
		, .Z(n_157994062));
	notech_ao4 i_84874980(.A(n_31268), .B(n_156394046), .C(n_156094043), .D(n_31301
		), .Z(n_158094063));
	notech_ao4 i_84774981(.A(n_30981), .B(n_30738), .C(n_30741), .D(n_33886)
		, .Z(n_158194064));
	notech_ao4 i_84674982(.A(n_31269), .B(n_156394046), .C(n_31302), .D(n_156094043
		), .Z(n_158294065));
	notech_ao4 i_84574983(.A(n_30738), .B(n_30983), .C(n_30741), .D(n_33885)
		, .Z(n_158394066));
	notech_ao4 i_84474984(.A(n_31270), .B(n_156394046), .C(n_156094043), .D(n_31303
		), .Z(n_158494067));
	notech_ao4 i_84374985(.A(n_30738), .B(n_30985), .C(n_30741), .D(n_33884)
		, .Z(n_158594068));
	notech_ao4 i_84274986(.A(n_31271), .B(n_156394046), .C(n_31304), .D(n_156094043
		), .Z(n_158694069));
	notech_ao4 i_84174987(.A(n_30738), .B(n_30987), .C(n_30741), .D(n_33883)
		, .Z(n_158794070));
	notech_ao4 i_84074988(.A(n_31272), .B(n_156394046), .C(n_31305), .D(n_156094043
		), .Z(n_158894071));
	notech_ao4 i_83974989(.A(n_30738), .B(n_30989), .C(n_30741), .D(n_33882)
		, .Z(n_158994072));
	notech_ao4 i_83874990(.A(n_31273), .B(n_156394046), .C(n_31306), .D(n_156094043
		), .Z(n_159094073));
	notech_ao4 i_83774991(.A(n_30738), .B(n_30991), .C(n_30741), .D(n_33881)
		, .Z(n_159194074));
	notech_ao4 i_83674992(.A(n_31274), .B(n_156394046), .C(n_31307), .D(n_156094043
		), .Z(n_159294075));
	notech_ao4 i_83574993(.A(n_30738), .B(n_30993), .C(n_30741), .D(n_33880)
		, .Z(n_159394076));
	notech_ao4 i_83474994(.A(n_31275), .B(n_156394046), .C(n_31308), .D(n_156094043
		), .Z(n_159494077));
	notech_ao4 i_83374995(.A(n_30738), .B(n_30995), .C(n_30741), .D(n_33879)
		, .Z(n_159594078));
	notech_ao4 i_83274996(.A(n_31276), .B(n_156394046), .C(n_31309), .D(n_156094043
		), .Z(n_159694079));
	notech_ao4 i_83174997(.A(n_30738), .B(n_30997), .C(n_30741), .D(n_33878)
		, .Z(n_159794080));
	notech_ao4 i_83074998(.A(n_31277), .B(n_54582), .C(n_54573), .D(n_31310)
		, .Z(n_159894081));
	notech_ao4 i_82974999(.A(n_55637), .B(n_30999), .C(n_54701), .D(n_33877)
		, .Z(n_159994082));
	notech_ao4 i_82875000(.A(n_31278), .B(n_54582), .C(n_31311), .D(n_54573)
		, .Z(n_160094083));
	notech_ao4 i_82775001(.A(n_55637), .B(n_31002), .C(n_54701), .D(n_33876)
		, .Z(n_160194084));
	notech_ao4 i_82675002(.A(n_31279), .B(n_54582), .C(n_31312), .D(n_54573)
		, .Z(n_160294085));
	notech_ao4 i_82575003(.A(n_55637), .B(n_31004), .C(n_54701), .D(n_33875)
		, .Z(n_160394086));
	notech_ao4 i_82475004(.A(n_31280), .B(n_54582), .C(n_31313), .D(n_54573)
		, .Z(n_160494087));
	notech_ao4 i_82375005(.A(n_55637), .B(n_31006), .C(n_54701), .D(n_33874)
		, .Z(n_160594088));
	notech_ao4 i_82275006(.A(n_31281), .B(n_54582), .C(n_31314), .D(n_54573)
		, .Z(n_160694089));
	notech_ao4 i_82175007(.A(n_55637), .B(n_31008), .C(n_54701), .D(n_33873)
		, .Z(n_160794090));
	notech_ao4 i_82075008(.A(n_31282), .B(n_54582), .C(n_31315), .D(n_54573)
		, .Z(n_160894091));
	notech_ao4 i_81975009(.A(n_55637), .B(n_31010), .C(n_54701), .D(n_33872)
		, .Z(n_160994092));
	notech_ao4 i_81875010(.A(n_31283), .B(n_54582), .C(n_31316), .D(n_54573)
		, .Z(n_161094093));
	notech_ao4 i_81775011(.A(n_55637), .B(n_31012), .C(n_54701), .D(n_33871)
		, .Z(n_161194094));
	notech_ao4 i_81675012(.A(n_31284), .B(n_54582), .C(n_31317), .D(n_54573)
		, .Z(n_161294095));
	notech_ao4 i_81575013(.A(n_55637), .B(n_31014), .C(n_54701), .D(n_33870)
		, .Z(n_161394096));
	notech_ao4 i_81475014(.A(n_31285), .B(n_54582), .C(n_31318), .D(n_54573)
		, .Z(n_161494097));
	notech_ao4 i_81375015(.A(n_55637), .B(n_31016), .C(n_33869), .D(n_54701)
		, .Z(n_161594098));
	notech_ao4 i_81275016(.A(n_31286), .B(n_54582), .C(n_31319), .D(n_54573)
		, .Z(n_161694099));
	notech_ao4 i_81175017(.A(n_55637), .B(n_31018), .C(n_54701), .D(n_33868)
		, .Z(n_161794100));
	notech_ao4 i_81075018(.A(n_31287), .B(n_156394046), .C(n_31320), .D(n_156094043
		), .Z(n_161894101));
	notech_ao4 i_80975019(.A(n_30738), .B(n_31020), .C(n_30741), .D(n_33867)
		, .Z(n_161994102));
	notech_ao4 i_80875020(.A(n_31288), .B(n_54582), .C(n_31321), .D(n_54573)
		, .Z(n_162094103));
	notech_ao4 i_80775021(.A(n_55637), .B(n_31022), .C(n_54701), .D(n_33866)
		, .Z(n_162194104));
	notech_ao4 i_80675022(.A(n_31289), .B(n_54582), .C(n_31322), .D(n_54573)
		, .Z(n_162294105));
	notech_ao4 i_80575023(.A(n_55637), .B(n_31024), .C(n_54701), .D(n_33865)
		, .Z(n_162394106));
	notech_ao4 i_80475024(.A(n_31290), .B(n_54582), .C(n_54573), .D(n_31323)
		, .Z(n_162494107));
	notech_ao4 i_80375025(.A(n_55637), .B(n_31026), .C(n_54701), .D(n_33864)
		, .Z(n_162594108));
	notech_ao4 i_80275026(.A(n_31291), .B(n_54582), .C(n_31324), .D(n_54573)
		, .Z(n_162694109));
	notech_ao4 i_80175027(.A(n_55637), .B(n_31028), .C(n_54701), .D(n_33863)
		, .Z(n_162794110));
	notech_ao4 i_80075028(.A(n_31292), .B(n_54582), .C(n_31325), .D(n_54573)
		, .Z(n_162894111));
	notech_ao4 i_79975029(.A(n_55637), .B(n_31030), .C(n_54701), .D(n_33862)
		, .Z(n_162994112));
	notech_nand2 i_79875030(.A(n_33160), .B(n_33179), .Z(n_163094113));
	notech_ao4 i_66575819(.A(n_30822), .B(n_78212538), .C(n_90793390), .D(n_33138
		), .Z(n_163194114));
	notech_or4 i_65675822(.A(instrc[88]), .B(instrc[90]), .C(n_33154), .D(n_33138
		), .Z(n_163394116));
	notech_ao4 i_79475034(.A(n_31261), .B(n_163394116), .C(n_33861), .D(n_30742
		), .Z(n_163494117));
	notech_or4 i_65275825(.A(instrc[89]), .B(n_33138), .C(n_104593528), .D(n_340061028
		), .Z(n_163794120));
	notech_ao4 i_79375035(.A(n_30737), .B(n_30967), .C(n_31294), .D(n_163794120
		), .Z(n_163894121));
	notech_ao4 i_79275036(.A(n_163394116), .B(n_31262), .C(n_30742), .D(n_33860
		), .Z(n_163994122));
	notech_ao4 i_79175037(.A(n_30737), .B(n_30969), .C(n_31295), .D(n_163794120
		), .Z(n_164094123));
	notech_ao4 i_79075038(.A(n_163394116), .B(n_31263), .C(n_30742), .D(n_33859
		), .Z(n_164194124));
	notech_ao4 i_78975039(.A(n_30737), .B(n_30971), .C(n_31296), .D(n_163794120
		), .Z(n_164294125));
	notech_ao4 i_78875040(.A(n_163394116), .B(n_31264), .C(n_30742), .D(n_33858
		), .Z(n_164394126));
	notech_ao4 i_78775041(.A(n_30737), .B(n_30973), .C(n_31297), .D(n_163794120
		), .Z(n_164494127));
	notech_ao4 i_78675042(.A(n_163394116), .B(n_31265), .C(n_30742), .D(n_33857
		), .Z(n_164594128));
	notech_ao4 i_78575043(.A(n_30737), .B(n_30975), .C(n_31298), .D(n_163794120
		), .Z(n_164694129));
	notech_ao4 i_78475044(.A(n_163394116), .B(n_31266), .C(n_30742), .D(n_33856
		), .Z(n_164794130));
	notech_ao4 i_78375045(.A(n_30737), .B(n_30977), .C(n_31299), .D(n_163794120
		), .Z(n_164894131));
	notech_ao4 i_78275046(.A(n_163394116), .B(n_31267), .C(n_30742), .D(n_33855
		), .Z(n_164994132));
	notech_ao4 i_78175047(.A(n_30737), .B(n_30979), .C(n_31300), .D(n_163794120
		), .Z(n_165094133));
	notech_ao4 i_78075048(.A(n_163394116), .B(n_31268), .C(n_30742), .D(n_33854
		), .Z(n_165194134));
	notech_ao4 i_77975049(.A(n_30737), .B(n_30981), .C(n_31301), .D(n_163794120
		), .Z(n_165294135));
	notech_ao4 i_77875050(.A(n_163394116), .B(n_31269), .C(n_30742), .D(n_33853
		), .Z(n_165394136));
	notech_ao4 i_77775051(.A(n_30737), .B(n_30983), .C(n_31302), .D(n_163794120
		), .Z(n_165494137));
	notech_ao4 i_77675052(.A(n_163394116), .B(n_31270), .C(n_30742), .D(n_33852
		), .Z(n_165594138));
	notech_ao4 i_77575053(.A(n_30737), .B(n_30985), .C(n_31303), .D(n_163794120
		), .Z(n_165694139));
	notech_ao4 i_77475054(.A(n_163394116), .B(n_31271), .C(n_30742), .D(n_33851
		), .Z(n_165794140));
	notech_ao4 i_77375055(.A(n_30737), .B(n_30987), .C(n_31304), .D(n_163794120
		), .Z(n_165894141));
	notech_ao4 i_77275056(.A(n_163394116), .B(n_31272), .C(n_30742), .D(n_33850
		), .Z(n_165994142));
	notech_ao4 i_77175057(.A(n_30737), .B(n_30989), .C(n_31305), .D(n_163794120
		), .Z(n_166094143));
	notech_ao4 i_77075058(.A(n_163394116), .B(n_31273), .C(n_30742), .D(n_33849
		), .Z(n_166194144));
	notech_ao4 i_76975059(.A(n_30737), .B(n_30991), .C(n_31306), .D(n_163794120
		), .Z(n_166294145));
	notech_ao4 i_76875060(.A(n_163394116), .B(n_31274), .C(n_30742), .D(n_33848
		), .Z(n_166394146));
	notech_ao4 i_76775061(.A(n_30737), .B(n_30993), .C(n_31307), .D(n_163794120
		), .Z(n_166494147));
	notech_ao4 i_76675062(.A(n_163394116), .B(n_31275), .C(n_30742), .D(n_33847
		), .Z(n_166594148));
	notech_ao4 i_76575063(.A(n_30737), .B(n_30995), .C(n_31308), .D(n_163794120
		), .Z(n_166694149));
	notech_ao4 i_76475064(.A(n_163394116), .B(n_31276), .C(n_30742), .D(n_33846
		), .Z(n_166794150));
	notech_ao4 i_76375065(.A(n_57642), .B(n_30997), .C(n_31309), .D(n_163794120
		), .Z(n_166894151));
	notech_ao4 i_76275066(.A(n_54553), .B(n_31277), .C(n_54544), .D(n_33845)
		, .Z(n_166994152));
	notech_ao4 i_76175067(.A(n_57642), .B(n_30999), .C(n_31310), .D(n_54564)
		, .Z(n_167094153));
	notech_ao4 i_76075068(.A(n_54553), .B(n_31278), .C(n_54544), .D(n_33844)
		, .Z(n_167194154));
	notech_ao4 i_75975069(.A(n_57642), .B(n_31002), .C(n_31311), .D(n_54564)
		, .Z(n_167294155));
	notech_ao4 i_75875070(.A(n_54553), .B(n_31279), .C(n_54544), .D(n_33843)
		, .Z(n_167394156));
	notech_ao4 i_75775071(.A(n_57642), .B(n_31004), .C(n_31312), .D(n_54564)
		, .Z(n_167494157));
	notech_ao4 i_75675072(.A(n_54553), .B(n_31280), .C(n_54544), .D(n_33842)
		, .Z(n_167594158));
	notech_ao4 i_75575073(.A(n_57642), .B(n_31006), .C(n_31313), .D(n_54564)
		, .Z(n_167694159));
	notech_ao4 i_75475074(.A(n_54553), .B(n_31281), .C(n_54544), .D(n_33841)
		, .Z(n_167794160));
	notech_ao4 i_75375075(.A(n_57642), .B(n_31008), .C(n_31314), .D(n_54564)
		, .Z(n_167894161));
	notech_ao4 i_75275076(.A(n_54553), .B(n_31282), .C(n_54544), .D(n_33840)
		, .Z(n_167994162));
	notech_ao4 i_75175077(.A(n_57642), .B(n_31010), .C(n_31315), .D(n_54564)
		, .Z(n_168094163));
	notech_ao4 i_75075078(.A(n_54553), .B(n_31283), .C(n_54544), .D(n_33839)
		, .Z(n_168194164));
	notech_ao4 i_74975079(.A(n_57642), .B(n_31012), .C(n_31316), .D(n_54564)
		, .Z(n_168294165));
	notech_ao4 i_74875080(.A(n_54553), .B(n_31284), .C(n_54544), .D(n_33838)
		, .Z(n_168394166));
	notech_ao4 i_74775081(.A(n_57642), .B(n_31014), .C(n_31317), .D(n_54564)
		, .Z(n_168494167));
	notech_ao4 i_74675082(.A(n_54553), .B(n_31285), .C(n_54544), .D(n_33837)
		, .Z(n_168594168));
	notech_ao4 i_74575083(.A(n_57642), .B(n_31016), .C(n_31318), .D(n_54564)
		, .Z(n_168694169));
	notech_ao4 i_74475084(.A(n_54553), .B(n_31286), .C(n_54544), .D(n_33836)
		, .Z(n_168794170));
	notech_ao4 i_74375085(.A(n_57642), .B(n_31018), .C(n_31319), .D(n_54564)
		, .Z(n_168894171));
	notech_ao4 i_74275086(.A(n_54553), .B(n_31287), .C(n_30742), .D(n_33835)
		, .Z(n_168994172));
	notech_ao4 i_74175087(.A(n_30737), .B(n_31020), .C(n_31320), .D(n_163794120
		), .Z(n_169094173));
	notech_ao4 i_74075088(.A(n_54553), .B(n_31288), .C(n_54544), .D(n_33834)
		, .Z(n_169194174));
	notech_ao4 i_73975089(.A(n_57642), .B(n_31022), .C(n_31321), .D(n_54564)
		, .Z(n_169294175));
	notech_ao4 i_73875090(.A(n_54553), .B(n_31289), .C(n_54544), .D(n_33833)
		, .Z(n_169394176));
	notech_ao4 i_73775091(.A(n_57642), .B(n_31024), .C(n_31322), .D(n_54564)
		, .Z(n_169494177));
	notech_ao4 i_73675092(.A(n_54553), .B(n_31290), .C(n_54544), .D(n_33832)
		, .Z(n_169594178));
	notech_ao4 i_73575093(.A(n_57642), .B(n_31026), .C(n_31323), .D(n_54564)
		, .Z(n_169694179));
	notech_ao4 i_73475094(.A(n_54553), .B(n_31291), .C(n_54544), .D(n_33831)
		, .Z(n_169794180));
	notech_ao4 i_73375095(.A(n_57642), .B(n_31028), .C(n_31324), .D(n_54564)
		, .Z(n_169894181));
	notech_ao4 i_73275096(.A(n_54553), .B(n_31292), .C(n_54544), .D(n_33830)
		, .Z(n_169994182));
	notech_ao4 i_73175097(.A(n_57642), .B(n_31030), .C(n_31325), .D(n_54564)
		, .Z(n_170094183));
	notech_xor2 i_774495(.A(all_cnt[2]), .B(n_325695672), .Z(n_170194184));
	notech_xor2 i_874494(.A(n_31372), .B(n_325795673), .Z(n_170294185));
	notech_nand3 i_21674300(.A(n_318095601), .B(n_30858), .C(instrc[99]), .Z
		(n_176794250));
	notech_nand3 i_34574171(.A(instrc[103]), .B(n_203294515), .C(n_308895531
		), .Z(n_176894251));
	notech_nor2 i_19583(.A(n_59104), .B(n_33002), .Z(n_176994252));
	notech_and2 i_26413(.A(n_61616), .B(n_170194184), .Z(n_177094253));
	notech_and2 i_26414(.A(n_61616), .B(n_170294185), .Z(n_177194254));
	notech_nand2 i_074501(.A(n_33176), .B(n_33161), .Z(n_203294515));
	notech_ao4 i_181172726(.A(n_54270), .B(n_31867), .C(n_54152), .D(n_31643
		), .Z(n_262395104));
	notech_ao4 i_181072727(.A(n_54290), .B(n_31803), .C(n_54280), .D(n_31931
		), .Z(n_262495105));
	notech_ao4 i_180872729(.A(n_54310), .B(n_31408), .C(n_54300), .D(n_31996
		), .Z(n_262695107));
	notech_ao4 i_180772730(.A(n_54329), .B(n_31964), .C(n_54320), .D(n_31899
		), .Z(n_262795108));
	notech_ao4 i_180572732(.A(n_54270), .B(n_31868), .C(n_54152), .D(n_31644
		), .Z(n_262995110));
	notech_ao4 i_180472733(.A(n_54290), .B(n_31804), .C(n_54280), .D(n_31932
		), .Z(n_263095111));
	notech_ao4 i_180272735(.A(n_54310), .B(n_31409), .C(n_54300), .D(n_31997
		), .Z(n_263295113));
	notech_ao4 i_180172736(.A(n_54329), .B(n_31965), .C(n_54320), .D(n_31900
		), .Z(n_263395114));
	notech_ao4 i_179972738(.A(n_54273), .B(n_31869), .C(n_54154), .D(n_31645
		), .Z(n_263595116));
	notech_ao4 i_179872739(.A(n_54293), .B(n_31805), .C(n_54282), .D(n_31933
		), .Z(n_263695117));
	notech_ao4 i_179672741(.A(n_54313), .B(n_31410), .C(n_54302), .D(n_31998
		), .Z(n_263895119));
	notech_ao4 i_179572742(.A(n_54331), .B(n_31966), .C(n_54322), .D(n_31901
		), .Z(n_263995120));
	notech_ao4 i_179372744(.A(n_54273), .B(n_31870), .C(n_54154), .D(n_31646
		), .Z(n_264195122));
	notech_ao4 i_179272745(.A(n_54293), .B(n_31806), .C(n_54282), .D(n_31934
		), .Z(n_264295123));
	notech_ao4 i_179072747(.A(n_54313), .B(n_31411), .C(n_54302), .D(n_31999
		), .Z(n_264495125));
	notech_ao4 i_178972748(.A(n_54331), .B(n_31967), .C(n_31902), .D(n_54322
		), .Z(n_264595126));
	notech_ao4 i_178772750(.A(n_54273), .B(n_31871), .C(n_54154), .D(n_31647
		), .Z(n_264795128));
	notech_ao4 i_178672751(.A(n_54293), .B(n_31807), .C(n_54282), .D(n_31935
		), .Z(n_264895129));
	notech_ao4 i_178472753(.A(n_54313), .B(n_31412), .C(n_54302), .D(n_32000
		), .Z(n_265095131));
	notech_ao4 i_178372754(.A(n_54331), .B(n_31968), .C(n_54322), .D(n_31903
		), .Z(n_265195132));
	notech_ao4 i_178172756(.A(n_54273), .B(n_31872), .C(n_54154), .D(n_31648
		), .Z(n_265395134));
	notech_ao4 i_178072757(.A(n_54293), .B(n_31808), .C(n_54282), .D(n_31936
		), .Z(n_265495135));
	notech_ao4 i_177872759(.A(n_54313), .B(n_31413), .C(n_54302), .D(n_32001
		), .Z(n_265695137));
	notech_ao4 i_177772760(.A(n_54331), .B(n_31969), .C(n_54322), .D(n_31904
		), .Z(n_265795138));
	notech_ao4 i_177572762(.A(n_54272), .B(n_31873), .C(n_54153), .D(n_31649
		), .Z(n_265995140));
	notech_ao4 i_177472763(.A(n_54292), .B(n_31809), .C(n_54281), .D(n_31937
		), .Z(n_266095141));
	notech_ao4 i_177272765(.A(n_54312), .B(n_31414), .C(n_54301), .D(n_32002
		), .Z(n_266295143));
	notech_ao4 i_177172766(.A(n_54330), .B(n_31970), .C(n_54321), .D(n_31905
		), .Z(n_266395144));
	notech_ao4 i_176972768(.A(n_54272), .B(n_31874), .C(n_54153), .D(n_31650
		), .Z(n_266595146));
	notech_ao4 i_176872769(.A(n_54292), .B(n_31810), .C(n_54281), .D(n_31938
		), .Z(n_266695147));
	notech_ao4 i_176672771(.A(n_54312), .B(n_31415), .C(n_54301), .D(n_32003
		), .Z(n_266895149));
	notech_ao4 i_176572772(.A(n_54330), .B(n_31971), .C(n_54321), .D(n_31906
		), .Z(n_266995150));
	notech_ao4 i_176372774(.A(n_54272), .B(n_31875), .C(n_54154), .D(n_31651
		), .Z(n_267195152));
	notech_ao4 i_176272775(.A(n_54292), .B(n_31811), .C(n_54282), .D(n_31939
		), .Z(n_267295153));
	notech_ao4 i_176072777(.A(n_54312), .B(n_31416), .C(n_54302), .D(n_32004
		), .Z(n_267495155));
	notech_ao4 i_175972778(.A(n_54331), .B(n_31972), .C(n_54322), .D(n_31907
		), .Z(n_267595156));
	notech_ao4 i_175772780(.A(n_54272), .B(n_31876), .C(n_54154), .D(n_31652
		), .Z(n_267795158));
	notech_ao4 i_175672781(.A(n_54292), .B(n_31812), .C(n_54282), .D(n_31940
		), .Z(n_267895159));
	notech_ao4 i_175472783(.A(n_54312), .B(n_31417), .C(n_54302), .D(n_32005
		), .Z(n_268095161));
	notech_ao4 i_175372784(.A(n_54331), .B(n_31973), .C(n_54322), .D(n_31908
		), .Z(n_268195162));
	notech_ao4 i_175172786(.A(n_54266), .B(n_31877), .C(n_54149), .D(n_31653
		), .Z(n_268395164));
	notech_ao4 i_175072787(.A(n_54286), .B(n_31813), .C(n_54277), .D(n_31941
		), .Z(n_268495165));
	notech_ao4 i_174872789(.A(n_54306), .B(n_31418), .C(n_54297), .D(n_32006
		), .Z(n_268695167));
	notech_ao4 i_174772790(.A(n_54329), .B(n_31974), .C(n_54317), .D(n_31909
		), .Z(n_268795168));
	notech_ao4 i_174572792(.A(n_54266), .B(n_31878), .C(n_54148), .D(n_31654
		), .Z(n_268995170));
	notech_ao4 i_174472793(.A(n_54286), .B(n_31814), .C(n_54276), .D(n_31943
		), .Z(n_269095171));
	notech_ao4 i_174272795(.A(n_54306), .B(n_31419), .C(n_54296), .D(n_32007
		), .Z(n_269295173));
	notech_ao4 i_174172796(.A(n_54326), .B(n_31975), .C(n_54316), .D(n_31910
		), .Z(n_269395174));
	notech_ao4 i_173972798(.A(n_54266), .B(n_31879), .C(n_54149), .D(n_31655
		), .Z(n_269595176));
	notech_ao4 i_173872799(.A(n_54286), .B(n_31815), .C(n_54277), .D(n_31944
		), .Z(n_269695177));
	notech_ao4 i_173672801(.A(n_54306), .B(n_31420), .C(n_54297), .D(n_32008
		), .Z(n_269895179));
	notech_ao4 i_173572802(.A(n_54325), .B(n_31976), .C(n_54317), .D(n_31911
		), .Z(n_269995180));
	notech_ao4 i_173372804(.A(n_54266), .B(n_31880), .C(n_54149), .D(n_31656
		), .Z(n_270195182));
	notech_ao4 i_173272805(.A(n_54286), .B(n_31816), .C(n_54277), .D(n_31945
		), .Z(n_270295183));
	notech_ao4 i_173072807(.A(n_54306), .B(n_31421), .C(n_54297), .D(n_32009
		), .Z(n_270495185));
	notech_ao4 i_172972808(.A(n_54326), .B(n_31977), .C(n_54317), .D(n_31912
		), .Z(n_270595186));
	notech_ao4 i_172772810(.A(n_54265), .B(n_31881), .C(n_54148), .D(n_31657
		), .Z(n_270895188));
	notech_ao4 i_172672811(.A(n_54285), .B(n_31817), .C(n_54276), .D(n_31946
		), .Z(n_270995189));
	notech_ao4 i_172472813(.A(n_54305), .B(n_31422), .C(n_54296), .D(n_32010
		), .Z(n_271195191));
	notech_ao4 i_172372814(.A(n_54326), .B(n_31978), .C(n_54316), .D(n_31913
		), .Z(n_271295192));
	notech_ao4 i_170972828(.A(n_54265), .B(n_31884), .C(n_54148), .D(n_31660
		), .Z(n_271495194));
	notech_ao4 i_170872829(.A(n_54285), .B(n_31820), .C(n_54276), .D(n_31949
		), .Z(n_271595195));
	notech_ao4 i_170672831(.A(n_54305), .B(n_31425), .C(n_54296), .D(n_32013
		), .Z(n_271795197));
	notech_ao4 i_170572832(.A(n_54325), .B(n_31981), .C(n_54316), .D(n_31916
		), .Z(n_271895198));
	notech_ao4 i_167972858(.A(n_54265), .B(n_31889), .C(n_54148), .D(n_31665
		), .Z(n_272095200));
	notech_ao4 i_167872859(.A(n_54285), .B(n_31825), .C(n_54276), .D(n_31954
		), .Z(n_272195201));
	notech_ao4 i_167672861(.A(n_54305), .B(n_31430), .C(n_54296), .D(n_32018
		), .Z(n_272395203));
	notech_ao4 i_167572862(.A(n_54325), .B(n_31986), .C(n_54316), .D(n_31921
		), .Z(n_272495204));
	notech_ao4 i_167372864(.A(n_54265), .B(n_31890), .C(n_54148), .D(n_31666
		), .Z(n_272695206));
	notech_ao4 i_167272865(.A(n_54285), .B(n_31826), .C(n_54276), .D(n_31955
		), .Z(n_272795207));
	notech_ao4 i_167072867(.A(n_54305), .B(n_31431), .C(n_54296), .D(n_32019
		), .Z(n_272995209));
	notech_ao4 i_166972868(.A(n_54325), .B(n_31987), .C(n_54316), .D(n_31922
		), .Z(n_273095210));
	notech_ao4 i_166772870(.A(n_54268), .B(n_31891), .C(n_54150), .D(n_31667
		), .Z(n_273295212));
	notech_ao4 i_166672871(.A(n_54288), .B(n_31827), .C(n_54278), .D(n_31956
		), .Z(n_273395213));
	notech_ao4 i_166472873(.A(n_54308), .B(n_31432), .C(n_54298), .D(n_32020
		), .Z(n_273595215));
	notech_ao4 i_166372874(.A(n_54325), .B(n_31988), .C(n_54318), .D(n_31923
		), .Z(n_273695216));
	notech_ao4 i_166172876(.A(n_54268), .B(n_31892), .C(n_54150), .D(n_31668
		), .Z(n_273895218));
	notech_ao4 i_166072877(.A(n_54288), .B(n_31828), .C(n_54278), .D(n_31957
		), .Z(n_273995219));
	notech_ao4 i_165872879(.A(n_54308), .B(n_31433), .C(n_54298), .D(n_32021
		), .Z(n_274195221));
	notech_ao4 i_165772880(.A(n_54327), .B(n_31989), .C(n_54318), .D(n_31924
		), .Z(n_274295222));
	notech_ao4 i_165572882(.A(n_54268), .B(n_31893), .C(n_54152), .D(n_31669
		), .Z(n_274495224));
	notech_ao4 i_165472883(.A(n_54288), .B(n_31829), .C(n_54280), .D(n_31958
		), .Z(n_274595225));
	notech_ao4 i_165272885(.A(n_54308), .B(n_31434), .C(n_54300), .D(n_32022
		), .Z(n_274795227));
	notech_ao4 i_165172886(.A(n_54327), .B(n_31990), .C(n_54320), .D(n_31925
		), .Z(n_274895228));
	notech_ao4 i_164972888(.A(n_54268), .B(n_31894), .C(n_54150), .D(n_31670
		), .Z(n_275195230));
	notech_ao4 i_164872889(.A(n_54288), .B(n_31830), .C(n_54278), .D(n_31959
		), .Z(n_275395231));
	notech_ao4 i_164672891(.A(n_54308), .B(n_31435), .C(n_54298), .D(n_32023
		), .Z(n_275595233));
	notech_ao4 i_164572892(.A(n_54329), .B(n_31991), .C(n_54318), .D(n_31926
		), .Z(n_275695234));
	notech_ao4 i_164372894(.A(n_54267), .B(n_31895), .C(n_54149), .D(n_31671
		), .Z(n_276195236));
	notech_ao4 i_164272895(.A(n_54287), .B(n_31831), .C(n_54277), .D(n_31960
		), .Z(n_276395237));
	notech_ao4 i_164072897(.A(n_54307), .B(n_31436), .C(n_54297), .D(n_32024
		), .Z(n_276595239));
	notech_ao4 i_163972898(.A(n_54327), .B(n_31992), .C(n_54317), .D(n_31927
		), .Z(n_276695240));
	notech_ao4 i_163772900(.A(n_54267), .B(n_31896), .C(n_54149), .D(n_31672
		), .Z(n_276895242));
	notech_ao4 i_163672901(.A(n_54287), .B(n_31832), .C(n_54277), .D(n_31961
		), .Z(n_276995243));
	notech_ao4 i_163472903(.A(n_54307), .B(n_31437), .C(n_54297), .D(n_32025
		), .Z(n_277195245));
	notech_ao4 i_163372904(.A(n_54326), .B(n_31993), .C(n_54317), .D(n_31928
		), .Z(n_277295246));
	notech_ao4 i_163172906(.A(n_54267), .B(n_31897), .C(n_54150), .D(n_31673
		), .Z(n_277495248));
	notech_ao4 i_163072907(.A(n_54287), .B(n_31833), .C(n_54278), .D(n_31962
		), .Z(n_277595249));
	notech_ao4 i_162872909(.A(n_54307), .B(n_31438), .C(n_54298), .D(n_32026
		), .Z(n_277795251));
	notech_ao4 i_162772910(.A(n_54326), .B(n_31994), .C(n_54318), .D(n_31929
		), .Z(n_277895252));
	notech_ao4 i_162572912(.A(n_54267), .B(n_31898), .C(n_54150), .D(n_31674
		), .Z(n_278095254));
	notech_ao4 i_162472913(.A(n_54287), .B(n_31834), .C(n_54278), .D(n_31963
		), .Z(n_278195255));
	notech_ao4 i_162272915(.A(n_54307), .B(n_31439), .C(n_54298), .D(n_32027
		), .Z(n_278395257));
	notech_ao4 i_162172916(.A(n_54327), .B(n_31995), .C(n_54318), .D(n_31930
		), .Z(n_278495258));
	notech_or4 i_7074524(.A(from_acu[4]), .B(from_acu[7]), .C(n_32938), .D(n_32937
		), .Z(n_278895262));
	notech_or4 i_831081(.A(from_acu[7]), .B(from_acu[6]), .C(from_acu[5]), .D
		(from_acu[4]), .Z(n_279195265));
	notech_or4 i_6974525(.A(from_acu[5]), .B(from_acu[4]), .C(from_acu[7]), 
		.D(n_30748), .Z(n_279395267));
	notech_ao4 i_161872919(.A(n_54349), .B(n_31931), .C(n_54339), .D(n_31643
		), .Z(n_279595268));
	notech_or4 i_6874526(.A(from_acu[7]), .B(from_acu[6]), .C(n_32937), .D(n_32936
		), .Z(n_279795270));
	notech_or4 i_6774527(.A(from_acu[7]), .B(from_acu[6]), .C(n_32937), .D(from_acu
		[4]), .Z(n_279895271));
	notech_ao4 i_161772920(.A(n_54369), .B(n_31996), .C(n_54359), .D(n_31803
		), .Z(n_279995272));
	notech_or4 i_6674528(.A(from_acu[7]), .B(from_acu[6]), .C(n_32936), .D(from_acu
		[5]), .Z(n_280295275));
	notech_or4 i_6174533(.A(n_32938), .B(from_acu[7]), .C(from_acu[5]), .D(n_32936
		), .Z(n_280395276));
	notech_ao4 i_161572922(.A(n_54389), .B(n_31867), .C(n_54379), .D(n_31408
		), .Z(n_280495277));
	notech_and4 i_5874536(.A(from_acu[5]), .B(from_acu[4]), .C(from_acu[6]),
		 .D(n_32939), .Z(n_280595278));
	notech_ao4 i_161472923(.A(n_54408), .B(n_31964), .C(n_31899), .D(n_54399
		), .Z(n_280695279));
	notech_ao4 i_161272925(.A(n_54349), .B(n_31932), .C(n_54339), .D(n_31644
		), .Z(n_280895281));
	notech_ao4 i_161172926(.A(n_54369), .B(n_31997), .C(n_54359), .D(n_31804
		), .Z(n_280995282));
	notech_ao4 i_160972928(.A(n_54389), .B(n_31868), .C(n_54379), .D(n_31409
		), .Z(n_281195284));
	notech_ao4 i_160872929(.A(n_54408), .B(n_31965), .C(n_31900), .D(n_54399
		), .Z(n_281295285));
	notech_ao4 i_160672931(.A(n_54349), .B(n_31933), .C(n_54339), .D(n_31645
		), .Z(n_281495287));
	notech_ao4 i_160572932(.A(n_54369), .B(n_31998), .C(n_54359), .D(n_31805
		), .Z(n_281595288));
	notech_ao4 i_160372934(.A(n_54389), .B(n_31869), .C(n_54379), .D(n_31410
		), .Z(n_281795290));
	notech_ao4 i_160272935(.A(n_54408), .B(n_31966), .C(n_31901), .D(n_54399
		), .Z(n_281895291));
	notech_ao4 i_160072937(.A(n_54349), .B(n_31934), .C(n_31646), .D(n_54339
		), .Z(n_282095293));
	notech_ao4 i_159972938(.A(n_54369), .B(n_31999), .C(n_54359), .D(n_31806
		), .Z(n_282195294));
	notech_ao4 i_159772940(.A(n_31870), .B(n_54389), .C(n_54379), .D(n_31411
		), .Z(n_282395296));
	notech_ao4 i_159672941(.A(n_54408), .B(n_31967), .C(n_31902), .D(n_54399
		), .Z(n_282495297));
	notech_ao4 i_159472943(.A(n_54348), .B(n_31935), .C(n_54338), .D(n_31647
		), .Z(n_282695299));
	notech_ao4 i_159372944(.A(n_54368), .B(n_32000), .C(n_54358), .D(n_31807
		), .Z(n_282795300));
	notech_ao4 i_159172946(.A(n_54388), .B(n_31871), .C(n_54378), .D(n_31412
		), .Z(n_282995302));
	notech_ao4 i_159072947(.A(n_54407), .B(n_31968), .C(n_31903), .D(n_54398
		), .Z(n_283095303));
	notech_ao4 i_158872949(.A(n_54348), .B(n_31936), .C(n_54338), .D(n_31648
		), .Z(n_283295305));
	notech_ao4 i_158772950(.A(n_54368), .B(n_32001), .C(n_54358), .D(n_31808
		), .Z(n_283395306));
	notech_ao4 i_158572952(.A(n_54388), .B(n_31872), .C(n_54378), .D(n_31413
		), .Z(n_283595308));
	notech_ao4 i_158472953(.A(n_54407), .B(n_31969), .C(n_31904), .D(n_54398
		), .Z(n_283695309));
	notech_ao4 i_158272955(.A(n_54348), .B(n_31937), .C(n_54338), .D(n_31649
		), .Z(n_283895311));
	notech_ao4 i_158172956(.A(n_54368), .B(n_32002), .C(n_54358), .D(n_31809
		), .Z(n_283995312));
	notech_ao4 i_157972958(.A(n_54388), .B(n_31873), .C(n_54378), .D(n_31414
		), .Z(n_284195314));
	notech_ao4 i_157872959(.A(n_54407), .B(n_31970), .C(n_31905), .D(n_54398
		), .Z(n_284295315));
	notech_ao4 i_157672961(.A(n_54348), .B(n_31938), .C(n_54338), .D(n_31650
		), .Z(n_284495317));
	notech_ao4 i_157572962(.A(n_54368), .B(n_32003), .C(n_54358), .D(n_31810
		), .Z(n_284595318));
	notech_ao4 i_157372964(.A(n_54388), .B(n_31874), .C(n_54378), .D(n_31415
		), .Z(n_284795320));
	notech_ao4 i_157272965(.A(n_54407), .B(n_31971), .C(n_31906), .D(n_54398
		), .Z(n_284895321));
	notech_ao4 i_157072967(.A(n_54351), .B(n_31939), .C(n_54340), .D(n_31651
		), .Z(n_285095323));
	notech_ao4 i_156972968(.A(n_54371), .B(n_32004), .C(n_54360), .D(n_31811
		), .Z(n_285195324));
	notech_ao4 i_156772970(.A(n_54391), .B(n_31875), .C(n_54380), .D(n_31416
		), .Z(n_285395326));
	notech_ao4 i_156672971(.A(n_54409), .B(n_31972), .C(n_31907), .D(n_54400
		), .Z(n_285495327));
	notech_ao4 i_156472973(.A(n_54351), .B(n_31940), .C(n_54340), .D(n_31652
		), .Z(n_285695329));
	notech_ao4 i_156372974(.A(n_54371), .B(n_32005), .C(n_54360), .D(n_31812
		), .Z(n_285795330));
	notech_ao4 i_156172976(.A(n_54391), .B(n_31876), .C(n_54380), .D(n_31417
		), .Z(n_285995332));
	notech_ao4 i_156072977(.A(n_54409), .B(n_31973), .C(n_31908), .D(n_54400
		), .Z(n_286095333));
	notech_ao4 i_155872979(.A(n_54351), .B(n_31941), .C(n_54340), .D(n_31653
		), .Z(n_286295335));
	notech_ao4 i_155772980(.A(n_54371), .B(n_32006), .C(n_54360), .D(n_31813
		), .Z(n_286395336));
	notech_ao4 i_155572982(.A(n_54391), .B(n_31877), .C(n_54380), .D(n_31418
		), .Z(n_286595338));
	notech_ao4 i_155472983(.A(n_54409), .B(n_31974), .C(n_31909), .D(n_54400
		), .Z(n_286695339));
	notech_ao4 i_155272985(.A(n_54351), .B(n_31943), .C(n_54340), .D(n_31654
		), .Z(n_286895341));
	notech_ao4 i_155172986(.A(n_54371), .B(n_32007), .C(n_54360), .D(n_31814
		), .Z(n_286995342));
	notech_ao4 i_154972988(.A(n_54391), .B(n_31878), .C(n_54380), .D(n_31419
		), .Z(n_287195344));
	notech_ao4 i_154872989(.A(n_54409), .B(n_31975), .C(n_31910), .D(n_54400
		), .Z(n_287295345));
	notech_ao4 i_154672991(.A(n_54350), .B(n_31944), .C(n_54339), .D(n_31655
		), .Z(n_287495347));
	notech_ao4 i_154572992(.A(n_54370), .B(n_32008), .C(n_54359), .D(n_31815
		), .Z(n_287595348));
	notech_ao4 i_154372994(.A(n_54390), .B(n_31879), .C(n_54379), .D(n_31420
		), .Z(n_287795350));
	notech_ao4 i_154272995(.A(n_54408), .B(n_31976), .C(n_31911), .D(n_54399
		), .Z(n_287895351));
	notech_ao4 i_154072997(.A(n_54350), .B(n_31945), .C(n_54339), .D(n_31656
		), .Z(n_288095353));
	notech_ao4 i_153972998(.A(n_54370), .B(n_32009), .C(n_54359), .D(n_31816
		), .Z(n_288195354));
	notech_ao4 i_153773000(.A(n_54390), .B(n_31880), .C(n_54379), .D(n_31421
		), .Z(n_288395356));
	notech_ao4 i_153673001(.A(n_54408), .B(n_31977), .C(n_31912), .D(n_54399
		), .Z(n_288495357));
	notech_ao4 i_153473003(.A(n_54350), .B(n_31946), .C(n_54340), .D(n_31657
		), .Z(n_288695359));
	notech_ao4 i_153373004(.A(n_54370), .B(n_32010), .C(n_54360), .D(n_31817
		), .Z(n_288795360));
	notech_ao4 i_153173006(.A(n_54390), .B(n_31881), .C(n_54380), .D(n_31422
		), .Z(n_288995362));
	notech_ao4 i_153073007(.A(n_54409), .B(n_31978), .C(n_31913), .D(n_54400
		), .Z(n_289095363));
	notech_ao4 i_152873009(.A(n_54350), .B(n_31947), .C(n_54340), .D(n_31658
		), .Z(n_289295365));
	notech_ao4 i_152773010(.A(n_54370), .B(n_32011), .C(n_54360), .D(n_31818
		), .Z(n_289395366));
	notech_ao4 i_152573012(.A(n_54390), .B(n_31882), .C(n_54380), .D(n_31423
		), .Z(n_289595368));
	notech_ao4 i_152473013(.A(n_54409), .B(n_31979), .C(n_31914), .D(n_54400
		), .Z(n_289695369));
	notech_ao4 i_152273015(.A(n_54344), .B(n_31948), .C(n_54335), .D(n_31659
		), .Z(n_289895371));
	notech_ao4 i_152173016(.A(n_54364), .B(n_32012), .C(n_54355), .D(n_31819
		), .Z(n_289995372));
	notech_ao4 i_151973018(.A(n_54384), .B(n_31883), .C(n_54375), .D(n_31424
		), .Z(n_290195374));
	notech_ao4 i_151873019(.A(n_54407), .B(n_31980), .C(n_31915), .D(n_54395
		), .Z(n_290295375));
	notech_ao4 i_151673021(.A(n_54344), .B(n_31949), .C(n_54334), .D(n_31660
		), .Z(n_290495377));
	notech_ao4 i_151573022(.A(n_54364), .B(n_32013), .C(n_54354), .D(n_31820
		), .Z(n_290595378));
	notech_ao4 i_151373024(.A(n_54384), .B(n_31884), .C(n_54374), .D(n_31425
		), .Z(n_290795380));
	notech_ao4 i_151273025(.A(n_54404), .B(n_31981), .C(n_31916), .D(n_54394
		), .Z(n_290895381));
	notech_ao4 i_151073027(.A(n_54344), .B(n_31950), .C(n_54335), .D(n_31661
		), .Z(n_291195383));
	notech_ao4 i_150973028(.A(n_54364), .B(n_32014), .C(n_54355), .D(n_31821
		), .Z(n_291295384));
	notech_ao4 i_150773030(.A(n_54384), .B(n_31885), .C(n_54375), .D(n_31426
		), .Z(n_291495386));
	notech_ao4 i_150673031(.A(n_54403), .B(n_31982), .C(n_31917), .D(n_54395
		), .Z(n_291595387));
	notech_ao4 i_150473033(.A(n_54344), .B(n_31951), .C(n_54335), .D(n_31662
		), .Z(n_291795389));
	notech_ao4 i_150373034(.A(n_54364), .B(n_32015), .C(n_54355), .D(n_31822
		), .Z(n_291895390));
	notech_ao4 i_150173036(.A(n_54384), .B(n_31886), .C(n_54375), .D(n_31427
		), .Z(n_292095392));
	notech_ao4 i_150073037(.A(n_54404), .B(n_31983), .C(n_31918), .D(n_54395
		), .Z(n_292195393));
	notech_ao4 i_149873039(.A(n_54343), .B(n_31952), .C(n_54334), .D(n_31663
		), .Z(n_292395395));
	notech_ao4 i_149773040(.A(n_54363), .B(n_32016), .C(n_31823), .D(n_54354
		), .Z(n_292495396));
	notech_ao4 i_149573042(.A(n_54383), .B(n_31887), .C(n_54374), .D(n_31428
		), .Z(n_292695398));
	notech_ao4 i_149473043(.A(n_54404), .B(n_31984), .C(n_31919), .D(n_54394
		), .Z(n_292795399));
	notech_ao4 i_149273045(.A(n_54343), .B(n_31953), .C(n_54334), .D(n_31664
		), .Z(n_292995401));
	notech_ao4 i_149173046(.A(n_54363), .B(n_32017), .C(n_54354), .D(n_31824
		), .Z(n_293095402));
	notech_ao4 i_148973048(.A(n_54383), .B(n_31888), .C(n_54374), .D(n_31429
		), .Z(n_293295404));
	notech_ao4 i_148873049(.A(n_54403), .B(n_31985), .C(n_31920), .D(n_54394
		), .Z(n_293395405));
	notech_ao4 i_148673051(.A(n_54343), .B(n_31954), .C(n_54334), .D(n_31665
		), .Z(n_293595407));
	notech_ao4 i_148573052(.A(n_54363), .B(n_32018), .C(n_54354), .D(n_31825
		), .Z(n_293695408));
	notech_ao4 i_148373054(.A(n_54383), .B(n_31889), .C(n_54374), .D(n_31430
		), .Z(n_293895410));
	notech_ao4 i_148273055(.A(n_54403), .B(n_31986), .C(n_31921), .D(n_54394
		), .Z(n_293995411));
	notech_ao4 i_148073057(.A(n_54343), .B(n_31955), .C(n_54334), .D(n_31666
		), .Z(n_294195413));
	notech_ao4 i_147973058(.A(n_54363), .B(n_32019), .C(n_54354), .D(n_31826
		), .Z(n_294295414));
	notech_ao4 i_147773060(.A(n_54383), .B(n_31890), .C(n_54374), .D(n_31431
		), .Z(n_294495416));
	notech_ao4 i_147673061(.A(n_54403), .B(n_31987), .C(n_31922), .D(n_54394
		), .Z(n_294595417));
	notech_ao4 i_147473063(.A(n_54346), .B(n_31956), .C(n_54336), .D(n_31667
		), .Z(n_294795419));
	notech_ao4 i_147373064(.A(n_54366), .B(n_32020), .C(n_54356), .D(n_31827
		), .Z(n_294895420));
	notech_ao4 i_147173066(.A(n_54386), .B(n_31891), .C(n_54376), .D(n_31432
		), .Z(n_295095422));
	notech_ao4 i_147073067(.A(n_54403), .B(n_31988), .C(n_31923), .D(n_54396
		), .Z(n_295195423));
	notech_ao4 i_146873069(.A(n_54346), .B(n_31957), .C(n_54336), .D(n_31668
		), .Z(n_295395425));
	notech_ao4 i_146773070(.A(n_54366), .B(n_32021), .C(n_54356), .D(n_31828
		), .Z(n_295495426));
	notech_ao4 i_146573072(.A(n_54386), .B(n_31892), .C(n_54376), .D(n_31433
		), .Z(n_295695428));
	notech_ao4 i_146473073(.A(n_54405), .B(n_31989), .C(n_31924), .D(n_54396
		), .Z(n_295795429));
	notech_ao4 i_146273075(.A(n_54346), .B(n_31958), .C(n_54338), .D(n_31669
		), .Z(n_295995431));
	notech_ao4 i_146173076(.A(n_54366), .B(n_32022), .C(n_54358), .D(n_31829
		), .Z(n_296095432));
	notech_ao4 i_145973078(.A(n_54386), .B(n_31893), .C(n_54378), .D(n_31434
		), .Z(n_296295434));
	notech_ao4 i_145873079(.A(n_54405), .B(n_31990), .C(n_31925), .D(n_54398
		), .Z(n_296395435));
	notech_ao4 i_145673081(.A(n_54346), .B(n_31959), .C(n_54336), .D(n_31670
		), .Z(n_296595437));
	notech_ao4 i_145573082(.A(n_54366), .B(n_32023), .C(n_54356), .D(n_31830
		), .Z(n_296695438));
	notech_ao4 i_145373084(.A(n_54386), .B(n_31894), .C(n_54376), .D(n_31435
		), .Z(n_296895440));
	notech_ao4 i_145273085(.A(n_54407), .B(n_31991), .C(n_31926), .D(n_54396
		), .Z(n_296995441));
	notech_ao4 i_145073087(.A(n_54345), .B(n_31960), .C(n_54335), .D(n_31671
		), .Z(n_297195443));
	notech_ao4 i_144973088(.A(n_54365), .B(n_32024), .C(n_54355), .D(n_31831
		), .Z(n_297295444));
	notech_ao4 i_144773090(.A(n_54385), .B(n_31895), .C(n_54375), .D(n_31436
		), .Z(n_297495446));
	notech_ao4 i_144673091(.A(n_54405), .B(n_31992), .C(n_31927), .D(n_54395
		), .Z(n_297595447));
	notech_ao4 i_144473093(.A(n_54345), .B(n_31961), .C(n_54335), .D(n_31672
		), .Z(n_297795449));
	notech_ao4 i_144373094(.A(n_54365), .B(n_32025), .C(n_54355), .D(n_31832
		), .Z(n_297895450));
	notech_ao4 i_144173096(.A(n_54385), .B(n_31896), .C(n_54375), .D(n_31437
		), .Z(n_298095452));
	notech_ao4 i_144073097(.A(n_54404), .B(n_31993), .C(n_31928), .D(n_54395
		), .Z(n_298195453));
	notech_ao4 i_143873099(.A(n_54345), .B(n_31962), .C(n_54336), .D(n_31673
		), .Z(n_298395455));
	notech_ao4 i_143773100(.A(n_54365), .B(n_32026), .C(n_54356), .D(n_31833
		), .Z(n_298495456));
	notech_ao4 i_143573102(.A(n_54385), .B(n_31897), .C(n_54376), .D(n_31438
		), .Z(n_298695458));
	notech_ao4 i_143473103(.A(n_54404), .B(n_31994), .C(n_31929), .D(n_54396
		), .Z(n_298795459));
	notech_ao4 i_143273105(.A(n_54345), .B(n_31963), .C(n_54336), .D(n_31674
		), .Z(n_298995461));
	notech_ao4 i_143173106(.A(n_54365), .B(n_32027), .C(n_54356), .D(n_31834
		), .Z(n_299095462));
	notech_ao4 i_142973108(.A(n_54385), .B(n_31898), .C(n_54376), .D(n_31439
		), .Z(n_299295464));
	notech_ao4 i_142873109(.A(n_54405), .B(n_31995), .C(n_31930), .D(n_54396
		), .Z(n_299395465));
	notech_ao4 i_142473113(.A(n_29047370), .B(n_33169), .C(n_29347373), .D(n_31294
		), .Z(n_299795467));
	notech_ao4 i_142373114(.A(n_30744), .B(n_30967), .C(n_28747367), .D(n_31261
		), .Z(n_299995468));
	notech_ao4 i_142273115(.A(n_29047370), .B(n_33103), .C(n_29347373), .D(n_31295
		), .Z(n_300095469));
	notech_ao4 i_142173116(.A(n_30744), .B(n_30969), .C(n_28747367), .D(n_31262
		), .Z(n_300195470));
	notech_ao4 i_142073117(.A(n_29047370), .B(n_33167), .C(n_29347373), .D(n_31296
		), .Z(n_300295471));
	notech_ao4 i_141973118(.A(n_30744), .B(n_30971), .C(n_28747367), .D(n_31263
		), .Z(n_300395472));
	notech_ao4 i_141873119(.A(n_29047370), .B(n_33118), .C(n_29347373), .D(n_31297
		), .Z(n_300595473));
	notech_ao4 i_141773120(.A(n_30744), .B(n_30973), .C(n_28747367), .D(n_31264
		), .Z(n_300695474));
	notech_ao4 i_141673121(.A(n_29047370), .B(n_33104), .C(n_29347373), .D(n_31298
		), .Z(n_300795475));
	notech_ao4 i_141573122(.A(n_30744), .B(n_30975), .C(n_28747367), .D(n_31265
		), .Z(n_300895476));
	notech_ao4 i_141473123(.A(n_29047370), .B(n_33135), .C(n_29347373), .D(n_31299
		), .Z(n_301095477));
	notech_ao4 i_141373124(.A(n_30744), .B(n_30977), .C(n_28747367), .D(n_31266
		), .Z(n_301395478));
	notech_ao4 i_141273125(.A(n_29047370), .B(n_33166), .C(n_29347373), .D(n_31300
		), .Z(n_301595479));
	notech_ao4 i_141173126(.A(n_30744), .B(n_30979), .C(n_28747367), .D(n_31267
		), .Z(n_301695480));
	notech_ao4 i_141073127(.A(n_29047370), .B(n_33165), .C(n_29347373), .D(n_31301
		), .Z(n_301795481));
	notech_ao4 i_140973128(.A(n_30744), .B(n_30981), .C(n_28747367), .D(n_31268
		), .Z(n_301895482));
	notech_ao4 i_140873129(.A(n_29047370), .B(n_33253), .C(n_29347373), .D(n_31302
		), .Z(n_301995483));
	notech_ao4 i_140773130(.A(n_30744), .B(n_30983), .C(n_28747367), .D(n_31269
		), .Z(n_302095484));
	notech_ao4 i_140673131(.A(n_29047370), .B(n_33168), .C(n_29347373), .D(n_31303
		), .Z(n_302195485));
	notech_ao4 i_140573132(.A(n_30744), .B(n_30985), .C(n_28747367), .D(n_31270
		), .Z(n_302295486));
	notech_ao4 i_140473133(.A(n_29047370), .B(n_33204), .C(n_29347373), .D(n_31304
		), .Z(n_302395487));
	notech_ao4 i_140373134(.A(n_30744), .B(n_30987), .C(n_28747367), .D(n_31271
		), .Z(n_302495488));
	notech_ao4 i_140273135(.A(n_29047370), .B(n_33258), .C(n_29347373), .D(n_31305
		), .Z(n_302595489));
	notech_ao4 i_140173136(.A(n_30744), .B(n_30989), .C(n_28747367), .D(n_31272
		), .Z(n_302795490));
	notech_ao4 i_140073137(.A(n_29047370), .B(n_33250), .C(n_29347373), .D(n_31306
		), .Z(n_302895491));
	notech_ao4 i_139973138(.A(n_30744), .B(n_30991), .C(n_28747367), .D(n_31273
		), .Z(n_302995492));
	notech_ao4 i_139873139(.A(n_29047370), .B(n_33213), .C(n_29347373), .D(n_31307
		), .Z(n_303095493));
	notech_ao4 i_139773140(.A(n_30744), .B(n_30993), .C(n_28747367), .D(n_31274
		), .Z(n_303295494));
	notech_ao4 i_139673141(.A(n_29047370), .B(n_33215), .C(n_29347373), .D(n_31308
		), .Z(n_303595495));
	notech_ao4 i_139573142(.A(n_30744), .B(n_30995), .C(n_28747367), .D(n_31275
		), .Z(n_303795496));
	notech_ao4 i_139473143(.A(n_55247), .B(n_33248), .C(n_55238), .D(n_31309
		), .Z(n_303895497));
	notech_ao4 i_139373144(.A(n_55619), .B(n_30997), .C(n_55258), .D(n_31276
		), .Z(n_303995498));
	notech_ao4 i_139273145(.A(n_55247), .B(n_33199), .C(n_55238), .D(n_31310
		), .Z(n_304095499));
	notech_ao4 i_139173146(.A(n_55619), .B(n_30999), .C(n_55258), .D(n_31277
		), .Z(n_304195500));
	notech_ao4 i_139073147(.A(n_55247), .B(n_33200), .C(n_55238), .D(n_31311
		), .Z(n_304395501));
	notech_ao4 i_138973148(.A(n_55619), .B(n_31002), .C(n_55258), .D(n_31278
		), .Z(n_304495502));
	notech_ao4 i_138873149(.A(n_55247), .B(n_33201), .C(n_55238), .D(n_31312
		), .Z(n_304595503));
	notech_ao4 i_138773150(.A(n_55619), .B(n_31004), .C(n_55258), .D(n_31279
		), .Z(n_304695504));
	notech_ao4 i_138673151(.A(n_55247), .B(n_33202), .C(n_55238), .D(n_31313
		), .Z(n_304895505));
	notech_ao4 i_138573152(.A(n_55619), .B(n_31006), .C(n_55258), .D(n_31280
		), .Z(n_305195506));
	notech_ao4 i_138473153(.A(n_55247), .B(n_33292), .C(n_55238), .D(n_31314
		), .Z(n_305395507));
	notech_ao4 i_138373154(.A(n_55619), .B(n_31008), .C(n_55258), .D(n_31281
		), .Z(n_305495508));
	notech_ao4 i_138273155(.A(n_55247), .B(n_33288), .C(n_55238), .D(n_31315
		), .Z(n_305595509));
	notech_ao4 i_138173156(.A(n_55619), .B(n_31010), .C(n_55258), .D(n_31282
		), .Z(n_305695510));
	notech_ao4 i_138073157(.A(n_55247), .B(n_33284), .C(n_55238), .D(n_31316
		), .Z(n_305795511));
	notech_ao4 i_137973158(.A(n_55619), .B(n_31012), .C(n_55258), .D(n_31283
		), .Z(n_305995512));
	notech_ao4 i_137873159(.A(n_55247), .B(n_33170), .C(n_55238), .D(n_31317
		), .Z(n_306095513));
	notech_ao4 i_137773160(.A(n_55619), .B(n_31014), .C(n_55258), .D(n_31284
		), .Z(n_306195514));
	notech_ao4 i_137673161(.A(n_55247), .B(n_33171), .C(n_55238), .D(n_31318
		), .Z(n_306295515));
	notech_ao4 i_137573162(.A(n_55619), .B(n_31016), .C(n_55258), .D(n_31285
		), .Z(n_306495516));
	notech_ao4 i_137273165(.A(n_55247), .B(n_33198), .C(n_29347373), .D(n_31320
		), .Z(n_306795517));
	notech_ao4 i_137173166(.A(n_30744), .B(n_31020), .C(n_28747367), .D(n_31287
		), .Z(n_306995518));
	notech_ao4 i_137073167(.A(n_55247), .B(n_33195), .C(n_55238), .D(n_31321
		), .Z(n_307095519));
	notech_ao4 i_136973168(.A(n_55619), .B(n_31022), .C(n_55258), .D(n_31288
		), .Z(n_307195520));
	notech_ao4 i_136873169(.A(n_55247), .B(n_33196), .C(n_55238), .D(n_31322
		), .Z(n_307395521));
	notech_ao4 i_136773170(.A(n_55619), .B(n_31024), .C(n_55258), .D(n_31289
		), .Z(n_307595522));
	notech_ao4 i_136673171(.A(n_55247), .B(n_33197), .C(n_55238), .D(n_31323
		), .Z(n_307695523));
	notech_ao4 i_136573172(.A(n_55619), .B(n_31026), .C(n_55258), .D(n_31290
		), .Z(n_307795524));
	notech_ao4 i_136473173(.A(n_55247), .B(n_33194), .C(n_55238), .D(n_31324
		), .Z(n_307895525));
	notech_ao4 i_136373174(.A(n_55619), .B(n_31028), .C(n_55258), .D(n_31291
		), .Z(n_307995526));
	notech_ao4 i_136273175(.A(n_55247), .B(n_33206), .C(n_55238), .D(n_31325
		), .Z(n_308195527));
	notech_ao4 i_136173176(.A(n_55619), .B(n_31030), .C(n_55258), .D(n_31292
		), .Z(n_308495528));
	notech_nand3 i_16317(.A(n_447368057), .B(instrc[103]), .C(n_436467948), 
		.Z(n_308695529));
	notech_ao4 i_129773240(.A(n_436467948), .B(n_33143), .C(n_33176), .D(n_33161
		), .Z(n_308895531));
	notech_nand2 i_66074519(.A(n_447368057), .B(n_176894251), .Z(n_309095532
		));
	notech_ao4 i_129473243(.A(n_309095532), .B(n_33989), .C(n_31294), .D(n_308695529
		), .Z(n_309295533));
	notech_or4 i_64174522(.A(instrc[100]), .B(n_30855), .C(n_30849), .D(instrc
		[102]), .Z(n_309595536));
	notech_ao4 i_129373244(.A(n_447368057), .B(n_30967), .C(n_309595536), .D
		(n_31261), .Z(n_309795537));
	notech_ao4 i_129273245(.A(n_309095532), .B(n_33988), .C(n_308695529), .D
		(n_31295), .Z(n_310095538));
	notech_ao4 i_129173246(.A(n_447368057), .B(n_30969), .C(n_309595536), .D
		(n_31262), .Z(n_310295539));
	notech_ao4 i_129073247(.A(n_309095532), .B(n_33987), .C(n_308695529), .D
		(n_31296), .Z(n_310395540));
	notech_ao4 i_128973248(.A(n_447368057), .B(n_30971), .C(n_309595536), .D
		(n_31263), .Z(n_310495541));
	notech_ao4 i_128873249(.A(n_309095532), .B(n_33986), .C(n_308695529), .D
		(n_31297), .Z(n_310595542));
	notech_ao4 i_128773250(.A(n_447368057), .B(n_30973), .C(n_309595536), .D
		(n_31264), .Z(n_310695543));
	notech_ao4 i_128673251(.A(n_309095532), .B(n_33985), .C(n_308695529), .D
		(n_31298), .Z(n_310895544));
	notech_ao4 i_128573252(.A(n_447368057), .B(n_30975), .C(n_309595536), .D
		(n_31265), .Z(n_310995545));
	notech_ao4 i_128473253(.A(n_309095532), .B(n_33984), .C(n_308695529), .D
		(n_31299), .Z(n_311095546));
	notech_ao4 i_128373254(.A(n_447368057), .B(n_30977), .C(n_309595536), .D
		(n_31266), .Z(n_311195547));
	notech_ao4 i_128273255(.A(n_309095532), .B(n_33983), .C(n_308695529), .D
		(n_31300), .Z(n_311395548));
	notech_ao4 i_128173256(.A(n_447368057), .B(n_30979), .C(n_309595536), .D
		(n_31267), .Z(n_311695549));
	notech_ao4 i_128073257(.A(n_309095532), .B(n_33982), .C(n_308695529), .D
		(n_31301), .Z(n_311895550));
	notech_ao4 i_127973258(.A(n_447368057), .B(n_30981), .C(n_309595536), .D
		(n_31268), .Z(n_311995551));
	notech_ao4 i_127873259(.A(n_309095532), .B(n_33981), .C(n_308695529), .D
		(n_31302), .Z(n_312095552));
	notech_ao4 i_127773260(.A(n_447368057), .B(n_30983), .C(n_309595536), .D
		(n_31269), .Z(n_312195553));
	notech_ao4 i_127673261(.A(n_309095532), .B(n_33980), .C(n_308695529), .D
		(n_31303), .Z(n_312295554));
	notech_ao4 i_127573262(.A(n_447368057), .B(n_30985), .C(n_309595536), .D
		(n_31270), .Z(n_312395555));
	notech_ao4 i_127473263(.A(n_309095532), .B(n_33979), .C(n_308695529), .D
		(n_31304), .Z(n_312495556));
	notech_ao4 i_127373264(.A(n_447368057), .B(n_30987), .C(n_309595536), .D
		(n_31271), .Z(n_312595557));
	notech_ao4 i_127273265(.A(n_309095532), .B(n_33978), .C(n_308695529), .D
		(n_31305), .Z(n_312695558));
	notech_ao4 i_127173266(.A(n_447368057), .B(n_30989), .C(n_309595536), .D
		(n_31272), .Z(n_312795559));
	notech_ao4 i_127073267(.A(n_309095532), .B(n_33977), .C(n_308695529), .D
		(n_31306), .Z(n_312895560));
	notech_ao4 i_126973268(.A(n_447368057), .B(n_30991), .C(n_309595536), .D
		(n_31273), .Z(n_312995561));
	notech_ao4 i_126873269(.A(n_309095532), .B(n_33976), .C(n_308695529), .D
		(n_31307), .Z(n_313095562));
	notech_ao4 i_126773270(.A(n_447368057), .B(n_30993), .C(n_309595536), .D
		(n_31274), .Z(n_313195563));
	notech_ao4 i_126673271(.A(n_309095532), .B(n_33975), .C(n_308695529), .D
		(n_31308), .Z(n_313295564));
	notech_ao4 i_126573272(.A(n_447368057), .B(n_30995), .C(n_309595536), .D
		(n_31275), .Z(n_313395565));
	notech_ao4 i_126473273(.A(n_309095532), .B(n_33974), .C(n_308695529), .D
		(n_31309), .Z(n_313495566));
	notech_ao4 i_126373274(.A(n_55610), .B(n_30997), .C(n_309595536), .D(n_31276
		), .Z(n_313595567));
	notech_ao4 i_126273275(.A(n_54968), .B(n_33973), .C(n_54849), .D(n_31310
		), .Z(n_313695568));
	notech_ao4 i_126173276(.A(n_55610), .B(n_30999), .C(n_54979), .D(n_31277
		), .Z(n_313895569));
	notech_ao4 i_126073277(.A(n_54968), .B(n_33972), .C(n_54849), .D(n_31311
		), .Z(n_314295570));
	notech_ao4 i_125973278(.A(n_55610), .B(n_31002), .C(n_54979), .D(n_31278
		), .Z(n_314395571));
	notech_ao4 i_125873279(.A(n_54968), .B(n_33971), .C(n_54849), .D(n_31312
		), .Z(n_314495572));
	notech_ao4 i_125773280(.A(n_55610), .B(n_31004), .C(n_54979), .D(n_31279
		), .Z(n_314595573));
	notech_ao4 i_125673281(.A(n_54968), .B(n_33970), .C(n_54849), .D(n_31313
		), .Z(n_314795574));
	notech_ao4 i_125573282(.A(n_55610), .B(n_31006), .C(n_54979), .D(n_31280
		), .Z(n_314895575));
	notech_ao4 i_125473283(.A(n_54968), .B(n_33969), .C(n_54849), .D(n_31314
		), .Z(n_314995576));
	notech_ao4 i_125373284(.A(n_55610), .B(n_31008), .C(n_54979), .D(n_31281
		), .Z(n_315095577));
	notech_ao4 i_125273285(.A(n_54968), .B(n_33968), .C(n_54849), .D(n_31315
		), .Z(n_315195578));
	notech_ao4 i_125173286(.A(n_55610), .B(n_31010), .C(n_54979), .D(n_31282
		), .Z(n_315295579));
	notech_ao4 i_125073287(.A(n_54968), .B(n_33967), .C(n_54849), .D(n_31316
		), .Z(n_315395580));
	notech_ao4 i_124973288(.A(n_55610), .B(n_31012), .C(n_54979), .D(n_31283
		), .Z(n_315495581));
	notech_ao4 i_124873289(.A(n_54968), .B(n_33966), .C(n_54849), .D(n_31317
		), .Z(n_315595582));
	notech_ao4 i_124773290(.A(n_55610), .B(n_31014), .C(n_54979), .D(n_31284
		), .Z(n_315695583));
	notech_ao4 i_124673291(.A(n_54968), .B(n_33965), .C(n_54849), .D(n_31318
		), .Z(n_315795584));
	notech_ao4 i_124573292(.A(n_55610), .B(n_31016), .C(n_54979), .D(n_31285
		), .Z(n_315895585));
	notech_ao4 i_124473293(.A(n_54968), .B(n_33964), .C(n_54849), .D(n_31319
		), .Z(n_315995586));
	notech_ao4 i_124373294(.A(n_55610), .B(n_31018), .C(n_54979), .D(n_31286
		), .Z(n_316195587));
	notech_ao4 i_124273295(.A(n_54968), .B(n_33963), .C(n_308695529), .D(n_31320
		), .Z(n_316495588));
	notech_ao4 i_124173296(.A(n_55610), .B(n_31020), .C(n_309595536), .D(n_31287
		), .Z(n_316695589));
	notech_ao4 i_124073297(.A(n_54968), .B(n_33962), .C(n_54849), .D(n_31321
		), .Z(n_316895590));
	notech_ao4 i_123973298(.A(n_55610), .B(n_31022), .C(n_54979), .D(n_31288
		), .Z(n_316995591));
	notech_ao4 i_123873299(.A(n_54968), .B(n_33961), .C(n_54849), .D(n_31322
		), .Z(n_317195592));
	notech_ao4 i_123773300(.A(n_55610), .B(n_31024), .C(n_54979), .D(n_31289
		), .Z(n_317295593));
	notech_ao4 i_123673301(.A(n_54968), .B(n_33960), .C(n_54849), .D(n_31323
		), .Z(n_317395594));
	notech_ao4 i_123573302(.A(n_55610), .B(n_31026), .C(n_54979), .D(n_31290
		), .Z(n_317495595));
	notech_ao4 i_123473303(.A(n_54968), .B(n_33959), .C(n_54849), .D(n_31324
		), .Z(n_317595596));
	notech_ao4 i_123373304(.A(n_55610), .B(n_31028), .C(n_54979), .D(n_31291
		), .Z(n_317695597));
	notech_ao4 i_123273305(.A(n_54968), .B(n_33958), .C(n_54849), .D(n_31325
		), .Z(n_317795598));
	notech_ao4 i_123173306(.A(n_55610), .B(n_31030), .C(n_54979), .D(n_31292
		), .Z(n_317895599));
	notech_ao4 i_122973308(.A(n_33140), .B(n_30865), .C(instrc[97]), .D(instrc
		[98]), .Z(n_318095601));
	notech_nand2 i_66174518(.A(n_447268056), .B(n_176794250), .Z(n_318295602
		));
	notech_or4 i_65874520(.A(n_33159), .B(n_29236), .C(instrc[96]), .D(n_30864
		), .Z(n_318895605));
	notech_ao4 i_122573312(.A(n_31261), .B(n_318895605), .C(n_318295602), .D
		(n_33957), .Z(n_318995606));
	notech_nao3 i_65374521(.A(n_447268056), .B(instrc[99]), .C(n_30751), .Z(n_319295608
		));
	notech_ao4 i_122473313(.A(n_447268056), .B(n_30967), .C(n_319295608), .D
		(n_31294), .Z(n_319395609));
	notech_ao4 i_122373314(.A(n_318895605), .B(n_31262), .C(n_318295602), .D
		(n_33956), .Z(n_319495610));
	notech_ao4 i_122273315(.A(n_447268056), .B(n_30969), .C(n_319295608), .D
		(n_31295), .Z(n_319595611));
	notech_ao4 i_122173316(.A(n_318895605), .B(n_31263), .C(n_318295602), .D
		(n_33955), .Z(n_319695612));
	notech_ao4 i_122073317(.A(n_447268056), .B(n_30971), .C(n_319295608), .D
		(n_31296), .Z(n_319795613));
	notech_ao4 i_121973318(.A(n_318895605), .B(n_31264), .C(n_318295602), .D
		(n_33954), .Z(n_319895614));
	notech_ao4 i_121873319(.A(n_447268056), .B(n_30973), .C(n_319295608), .D
		(n_31297), .Z(n_319995615));
	notech_ao4 i_121773320(.A(n_318895605), .B(n_31265), .C(n_318295602), .D
		(n_33953), .Z(n_320095616));
	notech_ao4 i_121673321(.A(n_447268056), .B(n_30975), .C(n_319295608), .D
		(n_31298), .Z(n_320195617));
	notech_ao4 i_121573322(.A(n_318895605), .B(n_31266), .C(n_318295602), .D
		(n_33952), .Z(n_320295618));
	notech_ao4 i_121473323(.A(n_447268056), .B(n_30977), .C(n_319295608), .D
		(n_31299), .Z(n_320395619));
	notech_ao4 i_121373324(.A(n_318895605), .B(n_31267), .C(n_318295602), .D
		(n_33951), .Z(n_320495620));
	notech_ao4 i_121273325(.A(n_447268056), .B(n_30979), .C(n_319295608), .D
		(n_31300), .Z(n_320595621));
	notech_ao4 i_121173326(.A(n_318895605), .B(n_31268), .C(n_318295602), .D
		(n_33950), .Z(n_320695622));
	notech_ao4 i_121073327(.A(n_447268056), .B(n_30981), .C(n_319295608), .D
		(n_31301), .Z(n_320795623));
	notech_ao4 i_120973328(.A(n_318895605), .B(n_31269), .C(n_318295602), .D
		(n_33949), .Z(n_320895624));
	notech_ao4 i_120873329(.A(n_447268056), .B(n_30983), .C(n_319295608), .D
		(n_31302), .Z(n_320995625));
	notech_ao4 i_120773330(.A(n_318895605), .B(n_31270), .C(n_318295602), .D
		(n_33948), .Z(n_321095626));
	notech_ao4 i_120673331(.A(n_447268056), .B(n_30985), .C(n_319295608), .D
		(n_31303), .Z(n_321195627));
	notech_ao4 i_120573332(.A(n_318895605), .B(n_31271), .C(n_318295602), .D
		(n_33947), .Z(n_321295628));
	notech_ao4 i_120473333(.A(n_447268056), .B(n_30987), .C(n_319295608), .D
		(n_31304), .Z(n_321395629));
	notech_ao4 i_120373334(.A(n_318895605), .B(n_31272), .C(n_318295602), .D
		(n_33946), .Z(n_321495630));
	notech_ao4 i_120273335(.A(n_447268056), .B(n_30989), .C(n_319295608), .D
		(n_31305), .Z(n_321595631));
	notech_ao4 i_120173336(.A(n_318895605), .B(n_31273), .C(n_318295602), .D
		(n_33945), .Z(n_321695632));
	notech_ao4 i_120073337(.A(n_447268056), .B(n_30991), .C(n_319295608), .D
		(n_31306), .Z(n_321795633));
	notech_ao4 i_119973338(.A(n_318895605), .B(n_31274), .C(n_318295602), .D
		(n_33944), .Z(n_321895634));
	notech_ao4 i_119873339(.A(n_447268056), .B(n_30993), .C(n_319295608), .D
		(n_31307), .Z(n_321995635));
	notech_ao4 i_119773340(.A(n_318895605), .B(n_31275), .C(n_318295602), .D
		(n_33943), .Z(n_322095636));
	notech_ao4 i_119673341(.A(n_447268056), .B(n_30995), .C(n_319295608), .D
		(n_31308), .Z(n_322195637));
	notech_ao4 i_119573342(.A(n_318895605), .B(n_31276), .C(n_318295602), .D
		(n_33942), .Z(n_322295638));
	notech_ao4 i_119473343(.A(n_55628), .B(n_30997), .C(n_319295608), .D(n_31309
		), .Z(n_322395639));
	notech_ao4 i_119373344(.A(n_54829), .B(n_31277), .C(n_54820), .D(n_33941
		), .Z(n_322495640));
	notech_ao4 i_119273345(.A(n_55628), .B(n_30999), .C(n_54840), .D(n_31310
		), .Z(n_322595641));
	notech_ao4 i_119173346(.A(n_54829), .B(n_31278), .C(n_54820), .D(n_33940
		), .Z(n_322695642));
	notech_ao4 i_119073347(.A(n_55628), .B(n_31002), .C(n_54840), .D(n_31311
		), .Z(n_322795643));
	notech_ao4 i_118973348(.A(n_54829), .B(n_31279), .C(n_54820), .D(n_33939
		), .Z(n_322895644));
	notech_ao4 i_118873349(.A(n_55628), .B(n_31004), .C(n_54840), .D(n_31312
		), .Z(n_322995645));
	notech_ao4 i_118773350(.A(n_54829), .B(n_31280), .C(n_54820), .D(n_33938
		), .Z(n_323095646));
	notech_ao4 i_118673351(.A(n_55628), .B(n_31006), .C(n_54840), .D(n_31313
		), .Z(n_323195647));
	notech_ao4 i_118573352(.A(n_54829), .B(n_31281), .C(n_54820), .D(n_33937
		), .Z(n_323295648));
	notech_ao4 i_118473353(.A(n_55628), .B(n_31008), .C(n_54840), .D(n_31314
		), .Z(n_323395649));
	notech_ao4 i_118373354(.A(n_54829), .B(n_31282), .C(n_54820), .D(n_33936
		), .Z(n_323495650));
	notech_ao4 i_118273355(.A(n_55628), .B(n_31010), .C(n_54840), .D(n_31315
		), .Z(n_323595651));
	notech_ao4 i_118173356(.A(n_54829), .B(n_31283), .C(n_54820), .D(n_33935
		), .Z(n_323695652));
	notech_ao4 i_118073357(.A(n_55628), .B(n_31012), .C(n_54840), .D(n_31316
		), .Z(n_323795653));
	notech_ao4 i_117973358(.A(n_54829), .B(n_31284), .C(n_54820), .D(n_33934
		), .Z(n_323895654));
	notech_ao4 i_117873359(.A(n_55628), .B(n_31014), .C(n_54840), .D(n_31317
		), .Z(n_323995655));
	notech_ao4 i_117773360(.A(n_54829), .B(n_31285), .C(n_54820), .D(n_33933
		), .Z(n_324095656));
	notech_ao4 i_117673361(.A(n_55628), .B(n_31016), .C(n_31318), .D(n_54840
		), .Z(n_324195657));
	notech_ao4 i_117573362(.A(n_54829), .B(n_31286), .C(n_54820), .D(n_33932
		), .Z(n_324295658));
	notech_ao4 i_117473363(.A(n_55628), .B(n_31018), .C(n_54840), .D(n_31319
		), .Z(n_324395659));
	notech_ao4 i_117373364(.A(n_54829), .B(n_31287), .C(n_318295602), .D(n_33931
		), .Z(n_324495660));
	notech_ao4 i_117273365(.A(n_55628), .B(n_31020), .C(n_319295608), .D(n_31320
		), .Z(n_324595661));
	notech_ao4 i_117173366(.A(n_54829), .B(n_31288), .C(n_54820), .D(n_33930
		), .Z(n_324695662));
	notech_ao4 i_117073367(.A(n_55628), .B(n_31022), .C(n_54840), .D(n_31321
		), .Z(n_324795663));
	notech_ao4 i_116973368(.A(n_54829), .B(n_31289), .C(n_54820), .D(n_33929
		), .Z(n_324895664));
	notech_ao4 i_116873369(.A(n_55628), .B(n_31024), .C(n_54840), .D(n_31322
		), .Z(n_324995665));
	notech_ao4 i_116773370(.A(n_54829), .B(n_31290), .C(n_54820), .D(n_33928
		), .Z(n_325095666));
	notech_ao4 i_116673371(.A(n_55628), .B(n_31026), .C(n_54840), .D(n_31323
		), .Z(n_325195667));
	notech_ao4 i_116573372(.A(n_54829), .B(n_31291), .C(n_54820), .D(n_33927
		), .Z(n_325295668));
	notech_ao4 i_116473373(.A(n_55628), .B(n_31028), .C(n_54840), .D(n_31324
		), .Z(n_325395669));
	notech_ao4 i_116373374(.A(n_54829), .B(n_31292), .C(n_54820), .D(n_33926
		), .Z(n_325495670));
	notech_ao4 i_116273375(.A(n_55628), .B(n_31030), .C(n_54840), .D(n_31325
		), .Z(n_325595671));
	notech_and2 i_88274515(.A(all_cnt[0]), .B(all_cnt[1]), .Z(n_325695672)
		);
	notech_nand3 i_974493(.A(all_cnt[0]), .B(all_cnt[1]), .C(all_cnt[2]), .Z
		(n_325795673));
	notech_ao4 i_160859152(.A(n_55187), .B(n_31628), .C(n_55198), .D(n_31311
		), .Z(n_326295678));
	notech_ao4 i_160759153(.A(n_56002), .B(n_31002), .C(n_55178), .D(n_31278
		), .Z(n_326395679));
	notech_nand2 i_26411(.A(n_61616), .B(n_31369), .Z(n_326695682));
	notech_nand2 i_99136645(.A(n_61616), .B(n_31370), .Z(n_326795683));
	notech_nand2 i_118111(.A(n_142793910), .B(n_142693909), .Z(write_data_27
		[0]));
	notech_nand2 i_218112(.A(n_142993912), .B(n_142893911), .Z(write_data_27
		[1]));
	notech_nand2 i_318113(.A(n_143193914), .B(n_143093913), .Z(write_data_27
		[2]));
	notech_nand2 i_418114(.A(n_143393916), .B(n_143293915), .Z(write_data_27
		[3]));
	notech_nand2 i_618116(.A(n_143593918), .B(n_143493917), .Z(write_data_27
		[5]));
	notech_nand2 i_718117(.A(n_143793920), .B(n_143693919), .Z(write_data_27
		[6]));
	notech_nand2 i_818118(.A(n_143993922), .B(n_143893921), .Z(write_data_27
		[7]));
	notech_nand2 i_918119(.A(n_144193924), .B(n_144093923), .Z(write_data_27
		[8]));
	notech_nand2 i_1018120(.A(n_144393926), .B(n_144293925), .Z(write_data_27
		[9]));
	notech_nand2 i_1118121(.A(n_144593928), .B(n_144493927), .Z(write_data_27
		[10]));
	notech_nand2 i_1218122(.A(n_144793930), .B(n_144693929), .Z(write_data_27
		[11]));
	notech_nand2 i_1318123(.A(n_144993932), .B(n_144893931), .Z(write_data_27
		[12]));
	notech_nand2 i_1418124(.A(n_145193934), .B(n_145093933), .Z(write_data_27
		[13]));
	notech_nand2 i_1518125(.A(n_145393936), .B(n_145293935), .Z(write_data_27
		[14]));
	notech_nand2 i_1618126(.A(n_145593938), .B(n_145493937), .Z(write_data_27
		[15]));
	notech_nand2 i_1718127(.A(n_145793940), .B(n_145693939), .Z(write_data_27
		[16]));
	notech_nand2 i_1918129(.A(n_145993942), .B(n_145893941), .Z(write_data_27
		[18]));
	notech_nand2 i_2018130(.A(n_146193944), .B(n_146093943), .Z(write_data_27
		[19]));
	notech_nand2 i_2118131(.A(n_146393946), .B(n_146293945), .Z(write_data_27
		[20]));
	notech_nand2 i_2218132(.A(n_146593948), .B(n_146493947), .Z(write_data_27
		[21]));
	notech_nand2 i_2318133(.A(n_146793950), .B(n_146693949), .Z(write_data_27
		[22]));
	notech_nand2 i_2418134(.A(n_146993952), .B(n_146893951), .Z(write_data_27
		[23]));
	notech_nand2 i_2518135(.A(n_147193954), .B(n_147093953), .Z(write_data_27
		[24]));
	notech_nand2 i_2618136(.A(n_147393956), .B(n_147293955), .Z(write_data_27
		[25]));
	notech_nand2 i_2718137(.A(n_147593958), .B(n_147493957), .Z(write_data_27
		[26]));
	notech_nand2 i_2818138(.A(n_147793960), .B(n_147693959), .Z(write_data_27
		[27]));
	notech_nand2 i_2918139(.A(n_147993962), .B(n_147893961), .Z(write_data_27
		[28]));
	notech_nand2 i_3018140(.A(n_148193964), .B(n_148093963), .Z(write_data_27
		[29]));
	notech_nand2 i_3118141(.A(n_148393966), .B(n_148293965), .Z(write_data_27
		[30]));
	notech_nand2 i_3218142(.A(n_148593968), .B(n_148493967), .Z(write_data_27
		[31]));
	notech_nand2 i_118239(.A(n_149593978), .B(n_149193974), .Z(write_data_28
		[0]));
	notech_nand2 i_218240(.A(n_149793980), .B(n_149693979), .Z(write_data_28
		[1]));
	notech_nand2 i_318241(.A(n_149993982), .B(n_149893981), .Z(write_data_28
		[2]));
	notech_nand2 i_418242(.A(n_150193984), .B(n_150093983), .Z(write_data_28
		[3]));
	notech_nand2 i_518243(.A(n_150393986), .B(n_150293985), .Z(write_data_28
		[4]));
	notech_nand2 i_618244(.A(n_150593988), .B(n_150493987), .Z(write_data_28
		[5]));
	notech_nand2 i_718245(.A(n_150793990), .B(n_150693989), .Z(write_data_28
		[6]));
	notech_nand2 i_818246(.A(n_150993992), .B(n_150893991), .Z(write_data_28
		[7]));
	notech_nand2 i_918247(.A(n_151193994), .B(n_151093993), .Z(write_data_28
		[8]));
	notech_nand2 i_1018248(.A(n_151393996), .B(n_151293995), .Z(write_data_28
		[9]));
	notech_nand2 i_1118249(.A(n_151593998), .B(n_151493997), .Z(write_data_28
		[10]));
	notech_nand2 i_1218250(.A(n_151794000), .B(n_151693999), .Z(write_data_28
		[11]));
	notech_nand2 i_1318251(.A(n_151994002), .B(n_151894001), .Z(write_data_28
		[12]));
	notech_nand2 i_1418252(.A(n_152194004), .B(n_152094003), .Z(write_data_28
		[13]));
	notech_nand2 i_1518253(.A(n_152394006), .B(n_152294005), .Z(write_data_28
		[14]));
	notech_nand2 i_1618254(.A(n_152594008), .B(n_152494007), .Z(write_data_28
		[15]));
	notech_nand2 i_1718255(.A(n_152794010), .B(n_152694009), .Z(write_data_28
		[16]));
	notech_nand2 i_1818256(.A(n_152994012), .B(n_152894011), .Z(write_data_28
		[17]));
	notech_nand2 i_1918257(.A(n_153194014), .B(n_153094013), .Z(write_data_28
		[18]));
	notech_nand2 i_2018258(.A(n_153394016), .B(n_153294015), .Z(write_data_28
		[19]));
	notech_nand2 i_2118259(.A(n_153594018), .B(n_153494017), .Z(write_data_28
		[20]));
	notech_nand2 i_2218260(.A(n_153794020), .B(n_153694019), .Z(write_data_28
		[21]));
	notech_nand2 i_2318261(.A(n_153994022), .B(n_153894021), .Z(write_data_28
		[22]));
	notech_nand2 i_2418262(.A(n_154194024), .B(n_154094023), .Z(write_data_28
		[23]));
	notech_nand2 i_2518263(.A(n_154394026), .B(n_154294025), .Z(write_data_28
		[24]));
	notech_nand2 i_2618264(.A(n_154594028), .B(n_154494027), .Z(write_data_28
		[25]));
	notech_nand2 i_2718265(.A(n_154794030), .B(n_154694029), .Z(write_data_28
		[26]));
	notech_nand2 i_2818266(.A(n_154994032), .B(n_154894031), .Z(write_data_28
		[27]));
	notech_nand2 i_2918267(.A(n_155194034), .B(n_155094033), .Z(write_data_28
		[28]));
	notech_nand2 i_3018268(.A(n_155394036), .B(n_155294035), .Z(write_data_28
		[29]));
	notech_nand2 i_3118269(.A(n_155594038), .B(n_155494037), .Z(write_data_28
		[30]));
	notech_nand2 i_3218270(.A(n_155794040), .B(n_155694039), .Z(write_data_28
		[31]));
	notech_nand2 i_118623(.A(n_156794050), .B(n_156494047), .Z(write_data_31
		[0]));
	notech_nand2 i_218624(.A(n_156994052), .B(n_156894051), .Z(write_data_31
		[1]));
	notech_nand2 i_318625(.A(n_157194054), .B(n_157094053), .Z(write_data_31
		[2]));
	notech_nand2 i_418626(.A(n_157394056), .B(n_157294055), .Z(write_data_31
		[3]));
	notech_nand2 i_518627(.A(n_157594058), .B(n_157494057), .Z(write_data_31
		[4]));
	notech_nand2 i_618628(.A(n_157794060), .B(n_157694059), .Z(write_data_31
		[5]));
	notech_nand2 i_718629(.A(n_157994062), .B(n_157894061), .Z(write_data_31
		[6]));
	notech_nand2 i_818630(.A(n_158194064), .B(n_158094063), .Z(write_data_31
		[7]));
	notech_nand2 i_918631(.A(n_158394066), .B(n_158294065), .Z(write_data_31
		[8]));
	notech_nand2 i_1018632(.A(n_158594068), .B(n_158494067), .Z(write_data_31
		[9]));
	notech_nand2 i_1118633(.A(n_158794070), .B(n_158694069), .Z(write_data_31
		[10]));
	notech_nand2 i_1218634(.A(n_158994072), .B(n_158894071), .Z(write_data_31
		[11]));
	notech_nand2 i_1318635(.A(n_159194074), .B(n_159094073), .Z(write_data_31
		[12]));
	notech_nand2 i_1418636(.A(n_159394076), .B(n_159294075), .Z(write_data_31
		[13]));
	notech_nand2 i_1518637(.A(n_159594078), .B(n_159494077), .Z(write_data_31
		[14]));
	notech_nand2 i_1618638(.A(n_159794080), .B(n_159694079), .Z(write_data_31
		[15]));
	notech_nand2 i_1718639(.A(n_159994082), .B(n_159894081), .Z(write_data_31
		[16]));
	notech_nand2 i_1818640(.A(n_160194084), .B(n_160094083), .Z(write_data_31
		[17]));
	notech_nand2 i_1918641(.A(n_160394086), .B(n_160294085), .Z(write_data_31
		[18]));
	notech_nand2 i_2018642(.A(n_160594088), .B(n_160494087), .Z(write_data_31
		[19]));
	notech_nand2 i_2118643(.A(n_160794090), .B(n_160694089), .Z(write_data_31
		[20]));
	notech_nand2 i_2218644(.A(n_160994092), .B(n_160894091), .Z(write_data_31
		[21]));
	notech_nand2 i_2318645(.A(n_161194094), .B(n_161094093), .Z(write_data_31
		[22]));
	notech_nand2 i_2418646(.A(n_161394096), .B(n_161294095), .Z(write_data_31
		[23]));
	notech_nand2 i_2518647(.A(n_161594098), .B(n_161494097), .Z(write_data_31
		[24]));
	notech_nand2 i_2618648(.A(n_161794100), .B(n_161694099), .Z(write_data_31
		[25]));
	notech_nand2 i_2718649(.A(n_161994102), .B(n_161894101), .Z(write_data_31
		[26]));
	notech_nand2 i_2818650(.A(n_162194104), .B(n_162094103), .Z(write_data_31
		[27]));
	notech_nand2 i_2918651(.A(n_162394106), .B(n_162294105), .Z(write_data_31
		[28]));
	notech_nand2 i_3018652(.A(n_162594108), .B(n_162494107), .Z(write_data_31
		[29]));
	notech_nand2 i_3118653(.A(n_162794110), .B(n_162694109), .Z(write_data_31
		[30]));
	notech_nand2 i_3218654(.A(n_162994112), .B(n_162894111), .Z(write_data_31
		[31]));
	notech_nand2 i_118751(.A(n_163894121), .B(n_163494117), .Z(write_data_32
		[0]));
	notech_nand2 i_218752(.A(n_164094123), .B(n_163994122), .Z(write_data_32
		[1]));
	notech_nand2 i_318753(.A(n_164294125), .B(n_164194124), .Z(write_data_32
		[2]));
	notech_nand2 i_418754(.A(n_164494127), .B(n_164394126), .Z(write_data_32
		[3]));
	notech_nand2 i_518755(.A(n_164694129), .B(n_164594128), .Z(write_data_32
		[4]));
	notech_nand2 i_618756(.A(n_164894131), .B(n_164794130), .Z(write_data_32
		[5]));
	notech_nand2 i_718757(.A(n_165094133), .B(n_164994132), .Z(write_data_32
		[6]));
	notech_nand2 i_818758(.A(n_165294135), .B(n_165194134), .Z(write_data_32
		[7]));
	notech_nand2 i_918759(.A(n_165494137), .B(n_165394136), .Z(write_data_32
		[8]));
	notech_nand2 i_1018760(.A(n_165694139), .B(n_165594138), .Z(write_data_32
		[9]));
	notech_nand2 i_1118761(.A(n_165894141), .B(n_165794140), .Z(write_data_32
		[10]));
	notech_nand2 i_1218762(.A(n_166094143), .B(n_165994142), .Z(write_data_32
		[11]));
	notech_nand2 i_1318763(.A(n_166294145), .B(n_166194144), .Z(write_data_32
		[12]));
	notech_nand2 i_1418764(.A(n_166494147), .B(n_166394146), .Z(write_data_32
		[13]));
	notech_nand2 i_1518765(.A(n_166694149), .B(n_166594148), .Z(write_data_32
		[14]));
	notech_nand2 i_1618766(.A(n_166894151), .B(n_166794150), .Z(write_data_32
		[15]));
	notech_nand2 i_1718767(.A(n_167094153), .B(n_166994152), .Z(write_data_32
		[16]));
	notech_nand2 i_1818768(.A(n_167294155), .B(n_167194154), .Z(write_data_32
		[17]));
	notech_nand2 i_1918769(.A(n_167494157), .B(n_167394156), .Z(write_data_32
		[18]));
	notech_nand2 i_2018770(.A(n_167694159), .B(n_167594158), .Z(write_data_32
		[19]));
	notech_nand2 i_2118771(.A(n_167894161), .B(n_167794160), .Z(write_data_32
		[20]));
	notech_nand2 i_2218772(.A(n_168094163), .B(n_167994162), .Z(write_data_32
		[21]));
	notech_nand2 i_2318773(.A(n_168294165), .B(n_168194164), .Z(write_data_32
		[22]));
	notech_nand2 i_2418774(.A(n_168494167), .B(n_168394166), .Z(write_data_32
		[23]));
	notech_nand2 i_2518775(.A(n_168694169), .B(n_168594168), .Z(write_data_32
		[24]));
	notech_nand2 i_2618776(.A(n_168894171), .B(n_168794170), .Z(write_data_32
		[25]));
	notech_nand2 i_2718777(.A(n_169094173), .B(n_168994172), .Z(write_data_32
		[26]));
	notech_nand2 i_2818778(.A(n_169294175), .B(n_169194174), .Z(write_data_32
		[27]));
	notech_nand2 i_2918779(.A(n_169494177), .B(n_169394176), .Z(write_data_32
		[28]));
	notech_nand2 i_3018780(.A(n_169694179), .B(n_169594178), .Z(write_data_32
		[29]));
	notech_nand2 i_3118781(.A(n_169894181), .B(n_169794180), .Z(write_data_32
		[30]));
	notech_nand2 i_3218782(.A(n_170094183), .B(n_169994182), .Z(write_data_32
		[31]));
	notech_xor2 i_10975830(.A(\eflags[7] ), .B(\eflags[11] ), .Z(\cond[12] )
		);
	notech_or2 i_117075828(.A(\eflags[6] ), .B(\cond[12] ), .Z(\cond[14] )
		);
	notech_or2 i_95675827(.A(\eflags[0] ), .B(\eflags[6] ), .Z(\cond[6] ));
	notech_mux2 i_3211710(.S(n_61455), .A(cr2[31]), .B(icr2[31]), .Z(n_8293)
		);
	notech_mux2 i_3111709(.S(n_61455), .A(cr2[30]), .B(icr2[30]), .Z(n_8287)
		);
	notech_mux2 i_2211700(.S(n_61455), .A(cr2[21]), .B(icr2[21]), .Z(n_8233)
		);
	notech_mux2 i_1711695(.S(n_61455), .A(cr2[16]), .B(icr2[16]), .Z(n_8203)
		);
	notech_mux2 i_1111689(.S(n_61455), .A(cr2[10]), .B(icr2[10]), .Z(n_8167)
		);
	notech_mux2 i_1011688(.S(n_61455), .A(cr2[9]), .B(icr2[9]), .Z(n_8161)
		);
	notech_mux2 i_911687(.S(n_61455), .A(cr2[8]), .B(icr2[8]), .Z(n_8155));
	notech_mux2 i_811686(.S(n_61455), .A(cr2[7]), .B(icr2[7]), .Z(n_8149));
	notech_mux2 i_711685(.S(n_61451), .A(cr2[6]), .B(icr2[6]), .Z(n_8143));
	notech_mux2 i_611684(.S(n_61451), .A(cr2[5]), .B(icr2[5]), .Z(n_8137));
	notech_mux2 i_511683(.S(n_61451), .A(cr2[4]), .B(icr2[4]), .Z(n_8131));
	notech_mux2 i_411682(.S(n_61455), .A(cr2[3]), .B(icr2[3]), .Z(n_8125));
	notech_mux2 i_311681(.S(n_61455), .A(cr2[2]), .B(icr2[2]), .Z(n_8119));
	notech_mux2 i_211680(.S(n_61455), .A(cr2[1]), .B(icr2[1]), .Z(n_8113));
	notech_mux2 i_111679(.S(n_61455), .A(cr2[0]), .B(icr2[0]), .Z(n_8107));
	notech_and4 i_111967(.A(n_262795108), .B(n_262695107), .C(n_262495105), 
		.D(n_262395104), .Z(to_acu101153[0]));
	notech_and4 i_211968(.A(n_263395114), .B(n_263295113), .C(n_263095111), 
		.D(n_262995110), .Z(to_acu101153[1]));
	notech_and4 i_311969(.A(n_263995120), .B(n_263895119), .C(n_263695117), 
		.D(n_263595116), .Z(to_acu101153[2]));
	notech_and4 i_411970(.A(n_264595126), .B(n_264495125), .C(n_264295123), 
		.D(n_264195122), .Z(to_acu101153[3]));
	notech_and4 i_511971(.A(n_265195132), .B(n_265095131), .C(n_264895129), 
		.D(n_264795128), .Z(to_acu101153[4]));
	notech_and4 i_611972(.A(n_265795138), .B(n_265695137), .C(n_265495135), 
		.D(n_265395134), .Z(to_acu101153[5]));
	notech_and4 i_711973(.A(n_266395144), .B(n_266295143), .C(n_266095141), 
		.D(n_265995140), .Z(to_acu101153[6]));
	notech_and4 i_811974(.A(n_266995150), .B(n_266895149), .C(n_266695147), 
		.D(n_266595146), .Z(to_acu101153[7]));
	notech_and4 i_911975(.A(n_267595156), .B(n_267495155), .C(n_267295153), 
		.D(n_267195152), .Z(to_acu101153[8]));
	notech_and4 i_1011976(.A(n_268195162), .B(n_268095161), .C(n_267895159),
		 .D(n_267795158), .Z(to_acu101153[9]));
	notech_and4 i_1111977(.A(n_268795168), .B(n_268695167), .C(n_268495165),
		 .D(n_268395164), .Z(to_acu101153[10]));
	notech_and4 i_1211978(.A(n_269395174), .B(n_269295173), .C(n_269095171),
		 .D(n_268995170), .Z(to_acu101153[11]));
	notech_and4 i_1311979(.A(n_269995180), .B(n_269895179), .C(n_269695177),
		 .D(n_269595176), .Z(to_acu101153[12]));
	notech_and4 i_1411980(.A(n_270595186), .B(n_270495185), .C(n_270295183),
		 .D(n_270195182), .Z(to_acu101153[13]));
	notech_and4 i_1511981(.A(n_271295192), .B(n_271195191), .C(n_270995189),
		 .D(n_270895188), .Z(to_acu101153[14]));
	notech_and4 i_1811984(.A(n_271895198), .B(n_271795197), .C(n_271595195),
		 .D(n_271495194), .Z(to_acu101153[17]));
	notech_and4 i_2311989(.A(n_272495204), .B(n_272395203), .C(n_272195201),
		 .D(n_272095200), .Z(to_acu101153[22]));
	notech_and4 i_2411990(.A(n_273095210), .B(n_272995209), .C(n_272795207),
		 .D(n_272695206), .Z(to_acu101153[23]));
	notech_and4 i_2511991(.A(n_273695216), .B(n_273595215), .C(n_273395213),
		 .D(n_273295212), .Z(to_acu101153[24]));
	notech_and4 i_2611992(.A(n_274295222), .B(n_274195221), .C(n_273995219),
		 .D(n_273895218), .Z(to_acu101153[25]));
	notech_and4 i_2711993(.A(n_274895228), .B(n_274795227), .C(n_274595225),
		 .D(n_274495224), .Z(to_acu101153[26]));
	notech_and4 i_2811994(.A(n_275695234), .B(n_275595233), .C(n_275395231),
		 .D(n_275195230), .Z(to_acu101153[27]));
	notech_and4 i_2911995(.A(n_276695240), .B(n_276595239), .C(n_276395237),
		 .D(n_276195236), .Z(to_acu101153[28]));
	notech_and4 i_3011996(.A(n_277295246), .B(n_277195245), .C(n_276995243),
		 .D(n_276895242), .Z(to_acu101153[29]));
	notech_and4 i_3111997(.A(n_277895252), .B(n_277795251), .C(n_277595249),
		 .D(n_277495248), .Z(to_acu101153[30]));
	notech_and4 i_3211998(.A(n_278495258), .B(n_278395257), .C(n_278195255),
		 .D(n_278095254), .Z(to_acu101153[31]));
	notech_and4 i_112223(.A(n_280695279), .B(n_280495277), .C(n_279995272), 
		.D(n_279595268), .Z(to_acu101153[32]));
	notech_and4 i_212224(.A(n_281295285), .B(n_281195284), .C(n_280995282), 
		.D(n_280895281), .Z(to_acu101153[33]));
	notech_and4 i_312225(.A(n_281895291), .B(n_281795290), .C(n_281595288), 
		.D(n_281495287), .Z(to_acu101153[34]));
	notech_and4 i_412226(.A(n_282495297), .B(n_282395296), .C(n_282195294), 
		.D(n_282095293), .Z(to_acu101153[35]));
	notech_and4 i_512227(.A(n_283095303), .B(n_282995302), .C(n_282795300), 
		.D(n_282695299), .Z(to_acu101153[36]));
	notech_and4 i_612228(.A(n_283695309), .B(n_283595308), .C(n_283395306), 
		.D(n_283295305), .Z(to_acu101153[37]));
	notech_and4 i_712229(.A(n_284295315), .B(n_284195314), .C(n_283995312), 
		.D(n_283895311), .Z(to_acu101153[38]));
	notech_and4 i_812230(.A(n_284895321), .B(n_284795320), .C(n_284595318), 
		.D(n_284495317), .Z(to_acu101153[39]));
	notech_and4 i_912231(.A(n_285495327), .B(n_285395326), .C(n_285195324), 
		.D(n_285095323), .Z(to_acu101153[40]));
	notech_and4 i_1012232(.A(n_286095333), .B(n_285995332), .C(n_285795330),
		 .D(n_285695329), .Z(to_acu101153[41]));
	notech_and4 i_1112233(.A(n_286695339), .B(n_286595338), .C(n_286395336),
		 .D(n_286295335), .Z(to_acu101153[42]));
	notech_and4 i_1212234(.A(n_287295345), .B(n_287195344), .C(n_286995342),
		 .D(n_286895341), .Z(to_acu101153[43]));
	notech_and4 i_1312235(.A(n_287895351), .B(n_287795350), .C(n_287595348),
		 .D(n_287495347), .Z(to_acu101153[44]));
	notech_and4 i_1412236(.A(n_288495357), .B(n_288395356), .C(n_288195354),
		 .D(n_288095353), .Z(to_acu101153[45]));
	notech_and4 i_1512237(.A(n_289095363), .B(n_288995362), .C(n_288795360),
		 .D(n_288695359), .Z(to_acu101153[46]));
	notech_and4 i_1612238(.A(n_289695369), .B(n_289595368), .C(n_289395366),
		 .D(n_289295365), .Z(to_acu101153[47]));
	notech_and4 i_1712239(.A(n_290295375), .B(n_290195374), .C(n_289995372),
		 .D(n_289895371), .Z(to_acu101153[48]));
	notech_and4 i_1812240(.A(n_290895381), .B(n_290795380), .C(n_290595378),
		 .D(n_290495377), .Z(to_acu101153[49]));
	notech_and4 i_1912241(.A(n_291595387), .B(n_291495386), .C(n_291295384),
		 .D(n_291195383), .Z(to_acu101153[50]));
	notech_and4 i_2012242(.A(n_292195393), .B(n_292095392), .C(n_291895390),
		 .D(n_291795389), .Z(to_acu101153[51]));
	notech_and4 i_2112243(.A(n_292795399), .B(n_292695398), .C(n_292495396),
		 .D(n_292395395), .Z(to_acu101153[52]));
	notech_and4 i_2212244(.A(n_293395405), .B(n_293295404), .C(n_293095402),
		 .D(n_292995401), .Z(to_acu101153[53]));
	notech_and4 i_2312245(.A(n_293995411), .B(n_293895410), .C(n_293695408),
		 .D(n_293595407), .Z(to_acu101153[54]));
	notech_and4 i_2412246(.A(n_294595417), .B(n_294495416), .C(n_294295414),
		 .D(n_294195413), .Z(to_acu101153[55]));
	notech_and4 i_2512247(.A(n_295195423), .B(n_295095422), .C(n_294895420),
		 .D(n_294795419), .Z(to_acu101153[56]));
	notech_and4 i_2612248(.A(n_295795429), .B(n_295695428), .C(n_295495426),
		 .D(n_295395425), .Z(to_acu101153[57]));
	notech_and4 i_2712249(.A(n_296395435), .B(n_296295434), .C(n_296095432),
		 .D(n_295995431), .Z(to_acu101153[58]));
	notech_and4 i_2812250(.A(n_296995441), .B(n_296895440), .C(n_296695438),
		 .D(n_296595437), .Z(to_acu101153[59]));
	notech_and4 i_2912251(.A(n_297595447), .B(n_297495446), .C(n_297295444),
		 .D(n_297195443), .Z(to_acu101153[60]));
	notech_and4 i_3012252(.A(n_298195453), .B(n_298095452), .C(n_297895450),
		 .D(n_297795449), .Z(to_acu101153[61]));
	notech_and4 i_3112253(.A(n_298795459), .B(n_298695458), .C(n_298495456),
		 .D(n_298395455), .Z(to_acu101153[62]));
	notech_and4 i_3212254(.A(n_299395465), .B(n_299295464), .C(n_299095462),
		 .D(n_298995461), .Z(to_acu101153[63]));
	notech_nand2 i_117855(.A(n_299995468), .B(n_299795467), .Z(write_data_25
		[0]));
	notech_nand2 i_217856(.A(n_300195470), .B(n_300095469), .Z(write_data_25
		[1]));
	notech_nand2 i_317857(.A(n_300395472), .B(n_300295471), .Z(write_data_25
		[2]));
	notech_nand2 i_417858(.A(n_300695474), .B(n_300595473), .Z(write_data_25
		[3]));
	notech_nand2 i_517859(.A(n_300895476), .B(n_300795475), .Z(write_data_25
		[4]));
	notech_nand2 i_617860(.A(n_301395478), .B(n_301095477), .Z(write_data_25
		[5]));
	notech_nand2 i_717861(.A(n_301695480), .B(n_301595479), .Z(write_data_25
		[6]));
	notech_nand2 i_817862(.A(n_301895482), .B(n_301795481), .Z(write_data_25
		[7]));
	notech_nand2 i_917863(.A(n_302095484), .B(n_301995483), .Z(write_data_25
		[8]));
	notech_nand2 i_1017864(.A(n_302295486), .B(n_302195485), .Z(write_data_25
		[9]));
	notech_nand2 i_1117865(.A(n_302495488), .B(n_302395487), .Z(write_data_25
		[10]));
	notech_nand2 i_1217866(.A(n_302795490), .B(n_302595489), .Z(write_data_25
		[11]));
	notech_nand2 i_1317867(.A(n_302995492), .B(n_302895491), .Z(write_data_25
		[12]));
	notech_nand2 i_1417868(.A(n_303295494), .B(n_303095493), .Z(write_data_25
		[13]));
	notech_nand2 i_1517869(.A(n_303795496), .B(n_303595495), .Z(write_data_25
		[14]));
	notech_nand2 i_1617870(.A(n_303995498), .B(n_303895497), .Z(write_data_25
		[15]));
	notech_nand2 i_1717871(.A(n_304195500), .B(n_304095499), .Z(write_data_25
		[16]));
	notech_nand2 i_1817872(.A(n_304495502), .B(n_304395501), .Z(write_data_25
		[17]));
	notech_nand2 i_1917873(.A(n_304695504), .B(n_304595503), .Z(write_data_25
		[18]));
	notech_nand2 i_2017874(.A(n_305195506), .B(n_304895505), .Z(write_data_25
		[19]));
	notech_nand2 i_2117875(.A(n_305495508), .B(n_305395507), .Z(write_data_25
		[20]));
	notech_nand2 i_2217876(.A(n_305695510), .B(n_305595509), .Z(write_data_25
		[21]));
	notech_nand2 i_2317877(.A(n_305995512), .B(n_305795511), .Z(write_data_25
		[22]));
	notech_nand2 i_2417878(.A(n_306195514), .B(n_306095513), .Z(write_data_25
		[23]));
	notech_nand2 i_2517879(.A(n_306495516), .B(n_306295515), .Z(write_data_25
		[24]));
	notech_nand2 i_2717881(.A(n_306995518), .B(n_306795517), .Z(write_data_25
		[26]));
	notech_nand2 i_2817882(.A(n_307195520), .B(n_307095519), .Z(write_data_25
		[27]));
	notech_nand2 i_2917883(.A(n_307595522), .B(n_307395521), .Z(write_data_25
		[28]));
	notech_nand2 i_3017884(.A(n_307795524), .B(n_307695523), .Z(write_data_25
		[29]));
	notech_nand2 i_3117885(.A(n_307995526), .B(n_307895525), .Z(write_data_25
		[30]));
	notech_nand2 i_3217886(.A(n_308495528), .B(n_308195527), .Z(write_data_25
		[31]));
	notech_nand2 i_118367(.A(n_309795537), .B(n_309295533), .Z(write_data_29
		[0]));
	notech_nand2 i_218368(.A(n_310295539), .B(n_310095538), .Z(write_data_29
		[1]));
	notech_nand2 i_318369(.A(n_310495541), .B(n_310395540), .Z(write_data_29
		[2]));
	notech_nand2 i_418370(.A(n_310695543), .B(n_310595542), .Z(write_data_29
		[3]));
	notech_nand2 i_518371(.A(n_310995545), .B(n_310895544), .Z(write_data_29
		[4]));
	notech_nand2 i_618372(.A(n_311195547), .B(n_311095546), .Z(write_data_29
		[5]));
	notech_nand2 i_718373(.A(n_311695549), .B(n_311395548), .Z(write_data_29
		[6]));
	notech_nand2 i_818374(.A(n_311995551), .B(n_311895550), .Z(write_data_29
		[7]));
	notech_nand2 i_918375(.A(n_312195553), .B(n_312095552), .Z(write_data_29
		[8]));
	notech_nand2 i_1018376(.A(n_312395555), .B(n_312295554), .Z(write_data_29
		[9]));
	notech_nand2 i_1118377(.A(n_312595557), .B(n_312495556), .Z(write_data_29
		[10]));
	notech_nand2 i_1218378(.A(n_312795559), .B(n_312695558), .Z(write_data_29
		[11]));
	notech_nand2 i_1318379(.A(n_312995561), .B(n_312895560), .Z(write_data_29
		[12]));
	notech_nand2 i_1418380(.A(n_313195563), .B(n_313095562), .Z(write_data_29
		[13]));
	notech_nand2 i_1518381(.A(n_313395565), .B(n_313295564), .Z(write_data_29
		[14]));
	notech_nand2 i_1618382(.A(n_313595567), .B(n_313495566), .Z(write_data_29
		[15]));
	notech_nand2 i_1718383(.A(n_313895569), .B(n_313695568), .Z(write_data_29
		[16]));
	notech_nand2 i_1818384(.A(n_314395571), .B(n_314295570), .Z(write_data_29
		[17]));
	notech_nand2 i_1918385(.A(n_314595573), .B(n_314495572), .Z(write_data_29
		[18]));
	notech_nand2 i_2018386(.A(n_314895575), .B(n_314795574), .Z(write_data_29
		[19]));
	notech_nand2 i_2118387(.A(n_315095577), .B(n_314995576), .Z(write_data_29
		[20]));
	notech_nand2 i_2218388(.A(n_315295579), .B(n_315195578), .Z(write_data_29
		[21]));
	notech_nand2 i_2318389(.A(n_315495581), .B(n_315395580), .Z(write_data_29
		[22]));
	notech_nand2 i_2418390(.A(n_315695583), .B(n_315595582), .Z(write_data_29
		[23]));
	notech_nand2 i_2518391(.A(n_315895585), .B(n_315795584), .Z(write_data_29
		[24]));
	notech_nand2 i_2618392(.A(n_316195587), .B(n_315995586), .Z(write_data_29
		[25]));
	notech_nand2 i_2718393(.A(n_316695589), .B(n_316495588), .Z(write_data_29
		[26]));
	notech_nand2 i_2818394(.A(n_316995591), .B(n_316895590), .Z(write_data_29
		[27]));
	notech_nand2 i_2918395(.A(n_317295593), .B(n_317195592), .Z(write_data_29
		[28]));
	notech_nand2 i_3018396(.A(n_317495595), .B(n_317395594), .Z(write_data_29
		[29]));
	notech_nand2 i_3118397(.A(n_317695597), .B(n_317595596), .Z(write_data_29
		[30]));
	notech_nand2 i_3218398(.A(n_317895599), .B(n_317795598), .Z(write_data_29
		[31]));
	notech_nand2 i_118495(.A(n_319395609), .B(n_318995606), .Z(write_data_30
		[0]));
	notech_nand2 i_218496(.A(n_319595611), .B(n_319495610), .Z(write_data_30
		[1]));
	notech_nand2 i_318497(.A(n_319795613), .B(n_319695612), .Z(write_data_30
		[2]));
	notech_nand2 i_418498(.A(n_319995615), .B(n_319895614), .Z(write_data_30
		[3]));
	notech_nand2 i_518499(.A(n_320195617), .B(n_320095616), .Z(write_data_30
		[4]));
	notech_nand2 i_618500(.A(n_320395619), .B(n_320295618), .Z(write_data_30
		[5]));
	notech_nand2 i_718501(.A(n_320595621), .B(n_320495620), .Z(write_data_30
		[6]));
	notech_nand2 i_818502(.A(n_320795623), .B(n_320695622), .Z(write_data_30
		[7]));
	notech_nand2 i_918503(.A(n_320995625), .B(n_320895624), .Z(write_data_30
		[8]));
	notech_nand2 i_1018504(.A(n_321195627), .B(n_321095626), .Z(write_data_30
		[9]));
	notech_nand2 i_1118505(.A(n_321395629), .B(n_321295628), .Z(write_data_30
		[10]));
	notech_nand2 i_1218506(.A(n_321595631), .B(n_321495630), .Z(write_data_30
		[11]));
	notech_nand2 i_1318507(.A(n_321795633), .B(n_321695632), .Z(write_data_30
		[12]));
	notech_nand2 i_1418508(.A(n_321995635), .B(n_321895634), .Z(write_data_30
		[13]));
	notech_nand2 i_1518509(.A(n_322195637), .B(n_322095636), .Z(write_data_30
		[14]));
	notech_nand2 i_1618510(.A(n_322395639), .B(n_322295638), .Z(write_data_30
		[15]));
	notech_nand2 i_1718511(.A(n_322595641), .B(n_322495640), .Z(write_data_30
		[16]));
	notech_nand2 i_1818512(.A(n_322795643), .B(n_322695642), .Z(write_data_30
		[17]));
	notech_nand2 i_1918513(.A(n_322995645), .B(n_322895644), .Z(write_data_30
		[18]));
	notech_nand2 i_2018514(.A(n_323195647), .B(n_323095646), .Z(write_data_30
		[19]));
	notech_nand2 i_2118515(.A(n_323395649), .B(n_323295648), .Z(write_data_30
		[20]));
	notech_nand2 i_2218516(.A(n_323595651), .B(n_323495650), .Z(write_data_30
		[21]));
	notech_nand2 i_2318517(.A(n_323795653), .B(n_323695652), .Z(write_data_30
		[22]));
	notech_nand2 i_2418518(.A(n_323995655), .B(n_323895654), .Z(write_data_30
		[23]));
	notech_nand2 i_2518519(.A(n_324195657), .B(n_324095656), .Z(write_data_30
		[24]));
	notech_nand2 i_2618520(.A(n_324395659), .B(n_324295658), .Z(write_data_30
		[25]));
	notech_nand2 i_2718521(.A(n_324595661), .B(n_324495660), .Z(write_data_30
		[26]));
	notech_nand2 i_2818522(.A(n_324795663), .B(n_324695662), .Z(write_data_30
		[27]));
	notech_nand2 i_2918523(.A(n_324995665), .B(n_324895664), .Z(write_data_30
		[28]));
	notech_nand2 i_3018524(.A(n_325195667), .B(n_325095666), .Z(write_data_30
		[29]));
	notech_nand2 i_3118525(.A(n_325395669), .B(n_325295668), .Z(write_data_30
		[30]));
	notech_nand2 i_3218526(.A(n_325595671), .B(n_325495670), .Z(write_data_30
		[31]));
	notech_ao4 i_6327530(.A(n_56380), .B(n_33003), .C(n_59109), .D(n_33001),
		 .Z(n_8094));
	notech_ao4 i_6227529(.A(n_56380), .B(n_33002), .C(n_59109), .D(n_33000),
		 .Z(n_8089));
	notech_ao4 i_6127528(.A(n_59104), .B(n_32999), .C(n_56380), .D(n_33001),
		 .Z(n_8084));
	notech_ao4 i_6027527(.A(n_56380), .B(n_33000), .C(n_59104), .D(n_32998),
		 .Z(n_8079));
	notech_ao4 i_5927526(.A(n_56380), .B(n_32999), .C(n_59104), .D(n_32997),
		 .Z(n_8074));
	notech_ao4 i_5827525(.A(n_56380), .B(n_32998), .C(n_59104), .D(n_32996),
		 .Z(n_8069));
	notech_ao4 i_5727524(.A(n_56380), .B(n_32997), .C(n_59104), .D(n_32995),
		 .Z(n_8064));
	notech_ao4 i_5627523(.A(n_56379), .B(n_32996), .C(n_59104), .D(n_32994),
		 .Z(n_8059));
	notech_ao4 i_5527522(.A(n_56379), .B(n_32995), .C(n_59104), .D(n_32993),
		 .Z(n_8054));
	notech_ao4 i_5427521(.A(n_56379), .B(n_32994), .C(n_59104), .D(n_32992),
		 .Z(n_8049));
	notech_ao4 i_5327520(.A(n_56379), .B(n_32993), .C(n_59104), .D(n_32991),
		 .Z(n_8044));
	notech_ao4 i_5227519(.A(n_56379), .B(n_32992), .C(n_59104), .D(n_32990),
		 .Z(n_8039));
	notech_ao4 i_5127518(.A(n_56379), .B(n_32991), .C(n_59104), .D(n_32989),
		 .Z(n_8034));
	notech_ao4 i_5027517(.A(n_56379), .B(n_32990), .C(n_59109), .D(n_32988),
		 .Z(n_8029));
	notech_ao4 i_4927516(.A(n_56380), .B(n_32989), .C(n_59109), .D(n_32987),
		 .Z(n_8024));
	notech_ao4 i_4827515(.A(n_56383), .B(n_32988), .C(n_59109), .D(n_32986),
		 .Z(n_8019));
	notech_ao4 i_4727514(.A(n_56383), .B(n_32987), .C(n_59109), .D(n_32985),
		 .Z(n_8014));
	notech_ao4 i_4627513(.A(n_56383), .B(n_32986), .C(n_59109), .D(n_32984),
		 .Z(n_8009));
	notech_ao4 i_4527512(.A(n_56383), .B(n_32985), .C(n_59114), .D(n_32983),
		 .Z(n_8004));
	notech_ao4 i_4427511(.A(n_56383), .B(n_32984), .C(n_59109), .D(n_32982),
		 .Z(n_7999));
	notech_ao4 i_4327510(.A(n_56383), .B(n_32983), .C(n_59109), .D(n_32981),
		 .Z(n_7994));
	notech_ao4 i_4227509(.A(n_56383), .B(n_32982), .C(n_59109), .D(n_32980),
		 .Z(n_7989));
	notech_ao4 i_4127508(.A(n_56383), .B(n_32981), .C(n_59109), .D(n_32979),
		 .Z(n_7984));
	notech_ao4 i_4027507(.A(n_56380), .B(n_32980), .C(n_59109), .D(n_32978),
		 .Z(n_7979));
	notech_ao4 i_3927506(.A(n_56380), .B(n_32979), .C(n_59109), .D(n_32977),
		 .Z(n_7974));
	notech_ao4 i_3827505(.A(n_56380), .B(n_32978), .C(n_59109), .D(n_32976),
		 .Z(n_7969));
	notech_ao4 i_3727504(.A(n_56380), .B(n_32977), .C(n_59109), .D(n_32975),
		 .Z(n_7964));
	notech_ao4 i_3627503(.A(n_56383), .B(n_32976), .C(n_59109), .D(n_32974),
		 .Z(n_7959));
	notech_ao4 i_3527502(.A(n_56383), .B(n_32975), .C(n_59109), .D(n_32973),
		 .Z(n_7954));
	notech_ao4 i_3427501(.A(n_56380), .B(n_32974), .C(n_59109), .D(n_32972),
		 .Z(n_7949));
	notech_and2 i_17488(.A(opb[0]), .B(n_61656), .Z(n_326895684));
	notech_and2 i_17489(.A(n_61656), .B(opb[1]), .Z(n_326995685));
	notech_and2 i_17490(.A(opb[2]), .B(n_61656), .Z(n_327095686));
	notech_and2 i_17491(.A(opb[3]), .B(n_61656), .Z(n_327195687));
	notech_and2 i_17492(.A(opb[4]), .B(n_61656), .Z(n_327295688));
	notech_and2 i_17493(.A(opb[5]), .B(n_61656), .Z(n_327395689));
	notech_and2 i_17494(.A(n_61656), .B(opb[6]), .Z(n_327495690));
	notech_and2 i_17495(.A(n_61656), .B(opb[8]), .Z(n_327595691));
	notech_and2 i_17496(.A(n_61656), .B(opb[9]), .Z(n_327695692));
	notech_and2 i_17497(.A(n_61656), .B(opb[10]), .Z(n_327795693));
	notech_and2 i_17498(.A(opb[11]), .B(n_61660), .Z(n_327895694));
	notech_and2 i_17499(.A(opb[12]), .B(n_61661), .Z(n_327995695));
	notech_and2 i_17500(.A(opb[13]), .B(n_61661), .Z(n_328095696));
	notech_and2 i_17501(.A(n_61661), .B(opb[14]), .Z(n_328195697));
	notech_ao3 i_17502(.A(n_61730), .B(opb[15]), .C(n_61880), .Z(n_328295698
		));
	notech_nand2 i_1818128(.A(n_326395679), .B(n_326295678), .Z(write_data_27
		[17]));
	notech_ao4 i_222466(.A(n_31370), .B(n_326695682), .C(n_326795683), .D(n_31369
		), .Z(n_8327));
	notech_and2 i_17455(.A(pt_fault), .B(n_33829), .Z(n_16495863));
	notech_and2 i_26593(.A(had_lgjmp), .B(\nbus_14542[31] ), .Z(pg_en));
	notech_nao3 i_261(.A(n_303060659), .B(instrc[125]), .C(n_303260661), .Z(n_2924
		));
	notech_nand3 i_235(.A(n_302460653), .B(n_304860677), .C(instrc[63]), .Z(n_2923
		));
	notech_or2 i_246(.A(n_302260651), .B(n_33146), .Z(n_2922));
	notech_nand3 i_247(.A(n_304060669), .B(n_1816), .C(instrc[55]), .Z(n_2921
		));
	notech_nao3 i_234(.A(n_303060659), .B(instrc[127]), .C(n_303260661), .Z(n_291060622
		));
	notech_nand3 i_206(.A(n_302460653), .B(n_304860677), .C(instrc[59]), .Z(n_2909
		));
	notech_or2 i_219(.A(n_302260651), .B(n_33145), .Z(n_290860621));
	notech_nand3 i_220(.A(n_304060669), .B(n_1816), .C(instrc[51]), .Z(n_2907
		));
	notech_nao3 i_205(.A(n_303060659), .B(n_61828), .C(n_303260661), .Z(n_2896
		));
	notech_nand3 i_179(.A(n_302460653), .B(n_304860677), .C(instrc[56]), .Z(n_2895
		));
	notech_or2 i_190(.A(n_302260651), .B(n_33144), .Z(n_2894));
	notech_nand3 i_191(.A(n_304060669), .B(n_1816), .C(instrc[48]), .Z(n_2893
		));
	notech_mux2 i_112255(.S(n_61275), .A(n_1411), .B(regs_14[0]), .Z(pc_out[
		0]));
	notech_mux2 i_212256(.S(n_61275), .A(n_1412), .B(regs_14[1]), .Z(pc_out[
		1]));
	notech_mux2 i_312257(.S(n_61275), .A(n_1413), .B(regs_14[2]), .Z(pc_out[
		2]));
	notech_mux2 i_412258(.S(n_61275), .A(n_1414), .B(regs_14[3]), .Z(pc_out[
		3]));
	notech_mux2 i_512259(.S(n_61275), .A(n_1415), .B(regs_14[4]), .Z(pc_out[
		4]));
	notech_mux2 i_612260(.S(n_61275), .A(n_1416), .B(regs_14[5]), .Z(pc_out[
		5]));
	notech_mux2 i_712261(.S(n_61275), .A(n_1417), .B(regs_14[6]), .Z(pc_out[
		6]));
	notech_mux2 i_812262(.S(n_61275), .A(n_1418), .B(regs_14[7]), .Z(pc_out[
		7]));
	notech_mux2 i_912263(.S(n_61275), .A(n_1419), .B(regs_14[8]), .Z(pc_out[
		8]));
	notech_mux2 i_1012264(.S(n_61275), .A(n_1420), .B(regs_14[9]), .Z(pc_out
		[9]));
	notech_mux2 i_1112265(.S(n_61275), .A(n_1421), .B(regs_14[10]), .Z(pc_out
		[10]));
	notech_mux2 i_1212266(.S(n_61275), .A(n_1422), .B(regs_14[11]), .Z(pc_out
		[11]));
	notech_mux2 i_1312267(.S(n_61275), .A(n_1423), .B(regs_14[12]), .Z(pc_out
		[12]));
	notech_mux2 i_1412268(.S(n_61275), .A(n_1424), .B(regs_14[13]), .Z(pc_out
		[13]));
	notech_mux2 i_1512269(.S(n_61275), .A(n_1425), .B(regs_14[14]), .Z(pc_out
		[14]));
	notech_mux2 i_1612270(.S(n_61275), .A(n_1426), .B(regs_14[15]), .Z(pc_out
		[15]));
	notech_mux2 i_1712271(.S(n_61275), .A(n_1427), .B(regs_14[16]), .Z(pc_out
		[16]));
	notech_mux2 i_1812272(.S(n_61279), .A(n_1428), .B(regs_14[17]), .Z(pc_out
		[17]));
	notech_mux2 i_1912273(.S(n_61279), .A(n_1429), .B(regs_14[18]), .Z(pc_out
		[18]));
	notech_mux2 i_2012274(.S(n_61279), .A(n_1430), .B(regs_14[19]), .Z(pc_out
		[19]));
	notech_mux2 i_2112275(.S(n_61279), .A(n_1431), .B(regs_14[20]), .Z(pc_out
		[20]));
	notech_mux2 i_2212276(.S(n_61279), .A(n_1432), .B(regs_14[21]), .Z(pc_out
		[21]));
	notech_mux2 i_2312277(.S(n_61281), .A(n_1433), .B(regs_14[22]), .Z(pc_out
		[22]));
	notech_mux2 i_2412278(.S(n_61281), .A(n_1434), .B(regs_14[23]), .Z(pc_out
		[23]));
	notech_mux2 i_2512279(.S(n_61279), .A(n_1435), .B(regs_14[24]), .Z(pc_out
		[24]));
	notech_mux2 i_2612280(.S(n_61281), .A(n_1436), .B(regs_14[25]), .Z(pc_out
		[25]));
	notech_mux2 i_2712281(.S(n_61279), .A(n_1437), .B(regs_14[26]), .Z(pc_out
		[26]));
	notech_mux2 i_2812282(.S(n_61279), .A(n_1438), .B(regs_14[27]), .Z(pc_out
		[27]));
	notech_mux2 i_2912283(.S(n_61275), .A(n_1439), .B(regs_14[28]), .Z(pc_out
		[28]));
	notech_mux2 i_3012284(.S(n_61279), .A(n_1440), .B(regs_14[29]), .Z(pc_out
		[29]));
	notech_mux2 i_3112285(.S(n_61279), .A(n_1441), .B(regs_14[30]), .Z(pc_out
		[30]));
	notech_mux2 i_3212286(.S(n_61279), .A(n_1442), .B(regs_14[31]), .Z(pc_out
		[31]));
	notech_nand2 i_12375829(.A(n_33829), .B(n_61094), .Z(\nbus_11278[0] ));
	notech_mux2 i_3011708(.S(n_61455), .A(cr2[29]), .B(icr2[29]), .Z(n_8281)
		);
	notech_mux2 i_2911707(.S(n_61456), .A(cr2[28]), .B(icr2[28]), .Z(n_8275)
		);
	notech_mux2 i_2811706(.S(n_61456), .A(cr2[27]), .B(icr2[27]), .Z(n_8269)
		);
	notech_mux2 i_2711705(.S(n_61456), .A(cr2[26]), .B(icr2[26]), .Z(n_8263)
		);
	notech_mux2 i_2611704(.S(n_61456), .A(cr2[25]), .B(icr2[25]), .Z(n_8257)
		);
	notech_mux2 i_2511703(.S(n_61456), .A(cr2[24]), .B(icr2[24]), .Z(n_8251)
		);
	notech_mux2 i_2411702(.S(n_61456), .A(cr2[23]), .B(icr2[23]), .Z(n_8245)
		);
	notech_mux2 i_2311701(.S(n_61456), .A(cr2[22]), .B(icr2[22]), .Z(n_8239)
		);
	notech_mux2 i_2111699(.S(n_61456), .A(cr2[20]), .B(icr2[20]), .Z(n_8227)
		);
	notech_mux2 i_2011698(.S(n_61456), .A(cr2[19]), .B(icr2[19]), .Z(n_8221)
		);
	notech_mux2 i_1911697(.S(n_61456), .A(cr2[18]), .B(icr2[18]), .Z(n_8215)
		);
	notech_mux2 i_1811696(.S(n_61455), .A(cr2[17]), .B(icr2[17]), .Z(n_8209)
		);
	notech_mux2 i_1611694(.S(n_61456), .A(cr2[15]), .B(icr2[15]), .Z(n_8197)
		);
	notech_mux2 i_1511693(.S(n_61456), .A(cr2[14]), .B(icr2[14]), .Z(n_8191)
		);
	notech_mux2 i_1411692(.S(n_61456), .A(cr2[13]), .B(icr2[13]), .Z(n_8185)
		);
	notech_mux2 i_1311691(.S(n_61456), .A(cr2[12]), .B(icr2[12]), .Z(n_8179)
		);
	notech_mux2 i_1211690(.S(n_61447), .A(cr2[11]), .B(icr2[11]), .Z(n_8173)
		);
	notech_mux2 i_3211742(.S(n_56952), .A(n_848), .B(n_847), .Z(n_17885));
	notech_mux2 i_3111741(.S(n_56951), .A(n_846), .B(n_845), .Z(n_17878));
	notech_mux2 i_3011740(.S(n_56952), .A(n_844), .B(n_843), .Z(n_17871));
	notech_mux2 i_2911739(.S(n_56952), .A(n_842), .B(n_841), .Z(n_17864));
	notech_mux2 i_2811738(.S(n_56952), .A(n_840), .B(n_839), .Z(n_17857));
	notech_mux2 i_2711737(.S(n_56951), .A(n_838), .B(n_837), .Z(n_17850));
	notech_mux2 i_2611736(.S(n_56951), .A(n_836), .B(n_835), .Z(n_17843));
	notech_mux2 i_2511735(.S(n_56951), .A(n_834), .B(n_833), .Z(n_17836));
	notech_mux2 i_2411734(.S(n_56951), .A(n_832), .B(n_831), .Z(n_17829));
	notech_mux2 i_2311733(.S(n_56951), .A(n_830), .B(n_829), .Z(n_17822));
	notech_mux2 i_2211732(.S(n_56952), .A(n_828), .B(n_827), .Z(n_17815));
	notech_mux2 i_2111731(.S(n_56952), .A(n_826), .B(n_825), .Z(n_17808));
	notech_mux2 i_2011730(.S(n_56952), .A(n_824), .B(n_823), .Z(n_17801));
	notech_mux2 i_1911729(.S(n_56952), .A(n_822), .B(n_821), .Z(n_17794));
	notech_mux2 i_1811728(.S(n_56952), .A(n_820), .B(n_819), .Z(n_17787));
	notech_mux2 i_1711727(.S(n_56952), .A(n_818), .B(n_817), .Z(n_17780));
	notech_mux2 i_1611726(.S(n_56952), .A(n_816), .B(n_815), .Z(n_17773));
	notech_mux2 i_1511725(.S(n_56952), .A(n_814), .B(n_813), .Z(n_17766));
	notech_mux2 i_1411724(.S(n_56952), .A(n_812), .B(n_811), .Z(n_17759));
	notech_mux2 i_1311723(.S(n_56952), .A(n_810), .B(n_809), .Z(n_17752));
	notech_mux2 i_1211722(.S(n_56951), .A(n_808), .B(n_807), .Z(n_17745));
	notech_mux2 i_1111721(.S(n_56952), .A(n_806), .B(n_805), .Z(n_17738));
	notech_mux2 i_1011720(.S(n_56952), .A(n_804), .B(n_803), .Z(n_17731));
	notech_mux2 i_911719(.S(n_56952), .A(n_802), .B(n_801), .Z(n_17724));
	notech_mux2 i_811718(.S(n_56952), .A(n_800), .B(n_799), .Z(n_17717));
	notech_mux2 i_711717(.S(n_56952), .A(n_798), .B(n_797), .Z(n_17710));
	notech_mux2 i_611716(.S(n_56952), .A(n_796), .B(n_795), .Z(n_17703));
	notech_mux2 i_511715(.S(n_56951), .A(n_794), .B(n_793), .Z(n_17696));
	notech_mux2 i_411714(.S(n_56951), .A(n_792), .B(n_791), .Z(n_17689));
	notech_mux2 i_311713(.S(n_56951), .A(n_790), .B(n_789), .Z(n_17682));
	notech_mux2 i_211712(.S(n_56951), .A(n_788), .B(n_787), .Z(n_17675));
	notech_mux2 i_111711(.S(n_56951), .A(n_786), .B(n_785), .Z(n_17668));
	notech_reg_set fsmf_reg_0(.CP(n_63362), .D(n_61898), .SD(n_62441), .Q(fsmf
		[0]));
	notech_reg_set fsmf_reg_1(.CP(n_63362), .D(n_61912), .SD(n_62441), .Q(fsmf
		[1]));
	notech_reg_set fsmf_reg_2(.CP(n_63362), .D(fsm[2]), .SD(n_62441), .Q(fsmf
		[2]));
	notech_reg_set fsmf_reg_3(.CP(n_63362), .D(fsm[3]), .SD(n_62441), .Q(fsmf
		[3]));
	notech_reg fsmf_reg_4(.CP(n_63362), .D(fsm[4]), .CD(n_62437), .Q(fsmf[4]
		));
	notech_reg calc_sz_reg_0(.CP(n_63362), .D(n_20813), .CD(n_62441), .Q(calc_sz
		[0]));
	notech_mux2 i_460(.S(n_330181778), .A(instrc[108]), .B(calc_sz[0]), .Z(n_20813
		));
	notech_reg calc_sz_reg_1(.CP(n_63362), .D(n_20820), .CD(n_62441), .Q(calc_sz
		[1]));
	notech_mux2 i_60598763(.S(n_330181778), .A(instrc[109]), .B(calc_sz[1]),
		 .Z(n_20820));
	notech_reg calc_sz_reg_2(.CP(n_63362), .D(n_20826), .CD(n_62441), .Q(calc_sz
		[2]));
	notech_mux2 i_65198762(.S(n_330181778), .A(instrc[110]), .B(calc_sz[2]),
		 .Z(n_20826));
	notech_reg calc_sz_reg_3(.CP(n_63362), .D(n_20832), .CD(n_62441), .Q(calc_sz
		[3]));
	notech_mux2 i_71898761(.S(n_330181778), .A(instrc[111]), .B(calc_sz[3]),
		 .Z(n_20832));
	notech_reg tsc_reg_0(.CP(n_63362), .D(n_328), .CD(n_62441), .Q(tsc[0])
		);
	notech_reg tsc_reg_1(.CP(n_63362), .D(n_330), .CD(n_62441), .Q(tsc[1])
		);
	notech_reg tsc_reg_2(.CP(n_63362), .D(n_332), .CD(n_62443), .Q(tsc[2])
		);
	notech_reg tsc_reg_3(.CP(n_63466), .D(n_334), .CD(n_62443), .Q(tsc[3])
		);
	notech_reg tsc_reg_4(.CP(n_63466), .D(n_336), .CD(n_62443), .Q(tsc[4])
		);
	notech_reg tsc_reg_5(.CP(n_63466), .D(n_338), .CD(n_62443), .Q(tsc[5])
		);
	notech_reg tsc_reg_6(.CP(n_63466), .D(n_340), .CD(n_62443), .Q(tsc[6])
		);
	notech_reg tsc_reg_7(.CP(n_63466), .D(n_342), .CD(n_62444), .Q(tsc[7])
		);
	notech_reg tsc_reg_8(.CP(n_63466), .D(n_344), .CD(n_62444), .Q(tsc[8])
		);
	notech_reg tsc_reg_9(.CP(n_63466), .D(n_346), .CD(n_62444), .Q(tsc[9])
		);
	notech_reg tsc_reg_10(.CP(n_63466), .D(n_348), .CD(n_62444), .Q(tsc[10])
		);
	notech_reg tsc_reg_11(.CP(n_63466), .D(n_350), .CD(n_62443), .Q(tsc[11])
		);
	notech_reg tsc_reg_12(.CP(n_63466), .D(n_352), .CD(n_62443), .Q(tsc[12])
		);
	notech_reg tsc_reg_13(.CP(n_63466), .D(n_354), .CD(n_62443), .Q(tsc[13])
		);
	notech_reg tsc_reg_14(.CP(n_63466), .D(n_356), .CD(n_62441), .Q(tsc[14])
		);
	notech_reg tsc_reg_15(.CP(n_63466), .D(n_358), .CD(n_62441), .Q(tsc[15])
		);
	notech_reg tsc_reg_16(.CP(n_63466), .D(n_360), .CD(n_62443), .Q(tsc[16])
		);
	notech_reg tsc_reg_17(.CP(n_63466), .D(n_362), .CD(n_62443), .Q(tsc[17])
		);
	notech_reg tsc_reg_18(.CP(n_63466), .D(n_364), .CD(n_62443), .Q(tsc[18])
		);
	notech_reg tsc_reg_19(.CP(n_63466), .D(n_366), .CD(n_62443), .Q(tsc[19])
		);
	notech_reg tsc_reg_20(.CP(n_63466), .D(n_368), .CD(n_62443), .Q(tsc[20])
		);
	notech_reg tsc_reg_21(.CP(n_63466), .D(n_370), .CD(n_62435), .Q(tsc[21])
		);
	notech_reg tsc_reg_22(.CP(n_63464), .D(n_372), .CD(n_62436), .Q(tsc[22])
		);
	notech_reg tsc_reg_23(.CP(n_63464), .D(n_374), .CD(n_62435), .Q(tsc[23])
		);
	notech_reg tsc_reg_24(.CP(n_63526), .D(n_376), .CD(n_62435), .Q(tsc[24])
		);
	notech_reg tsc_reg_25(.CP(n_63526), .D(n_378), .CD(n_62436), .Q(tsc[25])
		);
	notech_reg tsc_reg_26(.CP(n_63526), .D(n_380), .CD(n_62436), .Q(tsc[26])
		);
	notech_reg tsc_reg_27(.CP(n_63526), .D(n_382), .CD(n_62436), .Q(tsc[27])
		);
	notech_reg tsc_reg_28(.CP(n_63526), .D(n_384), .CD(n_62436), .Q(tsc[28])
		);
	notech_reg tsc_reg_29(.CP(n_63526), .D(n_386), .CD(n_62436), .Q(tsc[29])
		);
	notech_reg tsc_reg_30(.CP(n_63526), .D(n_388), .CD(n_62435), .Q(tsc[30])
		);
	notech_reg tsc_reg_31(.CP(n_63526), .D(n_390), .CD(n_62435), .Q(tsc[31])
		);
	notech_reg tsc_reg_32(.CP(n_63526), .D(n_392), .CD(n_62435), .Q(tsc[32])
		);
	notech_reg tsc_reg_33(.CP(n_63526), .D(n_394), .CD(n_62435), .Q(tsc[33])
		);
	notech_reg tsc_reg_34(.CP(n_63526), .D(n_396), .CD(n_62435), .Q(tsc[34])
		);
	notech_reg tsc_reg_35(.CP(n_63526), .D(n_398), .CD(n_62435), .Q(tsc[35])
		);
	notech_reg tsc_reg_36(.CP(n_63526), .D(n_400), .CD(n_62435), .Q(tsc[36])
		);
	notech_reg tsc_reg_37(.CP(n_63526), .D(n_402), .CD(n_62435), .Q(tsc[37])
		);
	notech_reg tsc_reg_38(.CP(n_63526), .D(n_404), .CD(n_62435), .Q(tsc[38])
		);
	notech_reg tsc_reg_39(.CP(n_63526), .D(n_406), .CD(n_62435), .Q(tsc[39])
		);
	notech_reg tsc_reg_40(.CP(n_63526), .D(n_408), .CD(n_62437), .Q(tsc[40])
		);
	notech_reg tsc_reg_41(.CP(n_63526), .D(n_410), .CD(n_62437), .Q(tsc[41])
		);
	notech_reg tsc_reg_42(.CP(n_63464), .D(n_412), .CD(n_62437), .Q(tsc[42])
		);
	notech_reg tsc_reg_43(.CP(n_63464), .D(n_414), .CD(n_62437), .Q(tsc[43])
		);
	notech_reg tsc_reg_44(.CP(n_63464), .D(n_416), .CD(n_62437), .Q(tsc[44])
		);
	notech_reg tsc_reg_45(.CP(n_63464), .D(n_418), .CD(n_62437), .Q(tsc[45])
		);
	notech_reg tsc_reg_46(.CP(n_63464), .D(n_420), .CD(n_62437), .Q(tsc[46])
		);
	notech_reg tsc_reg_47(.CP(n_63464), .D(n_422), .CD(n_62437), .Q(tsc[47])
		);
	notech_reg tsc_reg_48(.CP(n_63464), .D(n_424), .CD(n_62437), .Q(tsc[48])
		);
	notech_reg tsc_reg_49(.CP(n_63464), .D(n_426), .CD(n_62437), .Q(tsc[49])
		);
	notech_reg tsc_reg_50(.CP(n_63464), .D(n_428), .CD(n_62436), .Q(tsc[50])
		);
	notech_reg tsc_reg_51(.CP(n_63464), .D(n_430), .CD(n_62436), .Q(tsc[51])
		);
	notech_reg tsc_reg_52(.CP(n_63526), .D(n_432), .CD(n_62436), .Q(tsc[52])
		);
	notech_reg tsc_reg_53(.CP(n_63462), .D(n_434), .CD(n_62436), .Q(tsc[53])
		);
	notech_reg tsc_reg_54(.CP(n_63462), .D(n_436), .CD(n_62436), .Q(tsc[54])
		);
	notech_reg tsc_reg_55(.CP(n_63522), .D(n_438), .CD(n_62437), .Q(tsc[55])
		);
	notech_reg tsc_reg_56(.CP(n_63522), .D(n_440), .CD(n_62437), .Q(tsc[56])
		);
	notech_reg tsc_reg_57(.CP(n_63522), .D(n_442), .CD(n_62436), .Q(tsc[57])
		);
	notech_reg tsc_reg_58(.CP(n_63522), .D(n_444), .CD(n_62436), .Q(tsc[58])
		);
	notech_reg tsc_reg_59(.CP(n_63522), .D(n_446), .CD(n_62449), .Q(tsc[59])
		);
	notech_reg tsc_reg_60(.CP(n_63522), .D(n_448), .CD(n_62449), .Q(tsc[60])
		);
	notech_reg tsc_reg_61(.CP(n_63522), .D(n_450), .CD(n_62449), .Q(tsc[61])
		);
	notech_reg tsc_reg_62(.CP(n_63522), .D(n_452), .CD(n_62449), .Q(tsc[62])
		);
	notech_reg tsc_reg_63(.CP(n_63522), .D(n_454), .CD(n_62449), .Q(tsc[63])
		);
	notech_reg_set first_rep_reg(.CP(n_63522), .D(n_21004), .SD(n_62449), .Q
		(first_rep));
	notech_mux2 i_2426(.S(n_14216), .A(first_rep), .B(n_30524), .Z(n_21004)
		);
	notech_reg_set fecx_reg(.CP(n_63606), .D(n_21010), .SD(1'b1), .Q(fecx)
		);
	notech_mux2 i_2434(.S(n_8484), .A(fecx), .B(n_30730), .Z(n_21010));
	notech_reg sav_ecx_reg_0(.CP(n_63606), .D(n_21016), .CD(n_62449), .Q(sav_ecx
		[0]));
	notech_mux2 i_2442(.S(n_58832), .A(ecx[0]), .B(sav_ecx[0]), .Z(n_21016)
		);
	notech_reg sav_ecx_reg_1(.CP(n_63606), .D(n_21022), .CD(n_62449), .Q(sav_ecx
		[1]));
	notech_mux2 i_2450(.S(n_58832), .A(ecx[1]), .B(sav_ecx[1]), .Z(n_21022)
		);
	notech_reg sav_ecx_reg_2(.CP(n_63606), .D(n_21028), .CD(n_62449), .Q(sav_ecx
		[2]));
	notech_mux2 i_2458(.S(n_58832), .A(ecx[2]), .B(sav_ecx[2]), .Z(n_21028)
		);
	notech_nao3 i_178(.A(n_303060659), .B(n_61786), .C(n_303260661), .Z(n_2882
		));
	notech_reg sav_ecx_reg_3(.CP(n_63606), .D(n_21035), .CD(n_62448), .Q(sav_ecx
		[3]));
	notech_mux2 i_2466(.S(n_58832), .A(ecx[3]), .B(sav_ecx[3]), .Z(n_21035)
		);
	notech_nand3 i_148(.A(n_302460653), .B(n_304860677), .C(instrc[58]), .Z(n_2881
		));
	notech_reg sav_ecx_reg_4(.CP(n_63606), .D(n_21042), .CD(n_62448), .Q(sav_ecx
		[4]));
	notech_mux2 i_2474(.S(n_58832), .A(ecx[4]), .B(sav_ecx[4]), .Z(n_21042)
		);
	notech_or2 i_159(.A(n_302260651), .B(n_33151), .Z(n_2880));
	notech_reg sav_ecx_reg_5(.CP(n_63606), .D(n_21049), .CD(n_62448), .Q(sav_ecx
		[5]));
	notech_mux2 i_2482(.S(n_58833), .A(ecx[5]), .B(sav_ecx[5]), .Z(n_21049)
		);
	notech_nand3 i_163(.A(n_304060669), .B(n_1816), .C(instrc[50]), .Z(n_2879
		));
	notech_reg sav_ecx_reg_6(.CP(n_63606), .D(n_21057), .CD(n_62448), .Q(sav_ecx
		[6]));
	notech_mux2 i_2490(.S(n_58833), .A(ecx[6]), .B(sav_ecx[6]), .Z(n_21057)
		);
	notech_reg sav_ecx_reg_7(.CP(n_63606), .D(n_21064), .CD(n_62448), .Q(sav_ecx
		[7]));
	notech_mux2 i_2498(.S(n_58833), .A(ecx[7]), .B(sav_ecx[7]), .Z(n_21064)
		);
	notech_reg sav_ecx_reg_8(.CP(n_63606), .D(n_21071), .CD(n_62448), .Q(sav_ecx
		[8]));
	notech_mux2 i_2506(.S(n_58832), .A(ecx[8]), .B(sav_ecx[8]), .Z(n_21071)
		);
	notech_reg sav_ecx_reg_9(.CP(n_63606), .D(n_21078), .CD(n_62448), .Q(sav_ecx
		[9]));
	notech_mux2 i_2514(.S(n_58832), .A(ecx[9]), .B(sav_ecx[9]), .Z(n_21078)
		);
	notech_reg sav_ecx_reg_10(.CP(n_63606), .D(n_21085), .CD(n_62448), .Q(sav_ecx
		[10]));
	notech_mux2 i_2522(.S(n_58833), .A(ecx[10]), .B(sav_ecx[10]), .Z(n_21085
		));
	notech_reg sav_ecx_reg_11(.CP(n_63606), .D(n_21093), .CD(n_62448), .Q(sav_ecx
		[11]));
	notech_mux2 i_2530(.S(n_58827), .A(ecx[11]), .B(sav_ecx[11]), .Z(n_21093
		));
	notech_reg sav_ecx_reg_12(.CP(n_63606), .D(n_21100), .CD(n_62448), .Q(sav_ecx
		[12]));
	notech_mux2 i_2538(.S(n_58827), .A(ecx[12]), .B(sav_ecx[12]), .Z(n_21100
		));
	notech_reg sav_ecx_reg_13(.CP(n_63606), .D(n_21107), .CD(n_62452), .Q(sav_ecx
		[13]));
	notech_mux2 i_2546(.S(n_58827), .A(ecx[13]), .B(sav_ecx[13]), .Z(n_21107
		));
	notech_reg sav_ecx_reg_14(.CP(n_63606), .D(n_21114), .CD(n_62452), .Q(sav_ecx
		[14]));
	notech_mux2 i_2554(.S(n_58827), .A(ecx[14]), .B(sav_ecx[14]), .Z(n_21114
		));
	notech_reg sav_ecx_reg_15(.CP(n_63606), .D(n_21121), .CD(n_62452), .Q(sav_ecx
		[15]));
	notech_mux2 i_2562(.S(n_58827), .A(ecx[15]), .B(sav_ecx[15]), .Z(n_21121
		));
	notech_reg sav_ecx_reg_16(.CP(n_63606), .D(n_21128), .CD(n_62452), .Q(sav_ecx
		[16]));
	notech_mux2 i_2570(.S(n_58827), .A(ecx[16]), .B(sav_ecx[16]), .Z(n_21128
		));
	notech_nao3 i_147(.A(n_303060659), .B(n_61944), .C(n_303260661), .Z(n_2868
		));
	notech_reg sav_ecx_reg_17(.CP(n_63522), .D(n_21134), .CD(n_62452), .Q(sav_ecx
		[17]));
	notech_mux2 i_2578(.S(n_58832), .A(ecx[17]), .B(sav_ecx[17]), .Z(n_21134
		));
	notech_and4 i_227949(.A(n_2865), .B(n_313460762), .C(n_2853), .D(n_2866)
		, .Z(n_2867));
	notech_reg sav_ecx_reg_18(.CP(n_63606), .D(n_21140), .CD(n_62453), .Q(sav_ecx
		[18]));
	notech_mux2 i_2586(.S(n_58832), .A(ecx[18]), .B(sav_ecx[18]), .Z(n_21140
		));
	notech_nand3 i_115(.A(n_302460653), .B(n_304860677), .C(instrc[57]), .Z(n_2866
		));
	notech_reg sav_ecx_reg_19(.CP(n_63524), .D(n_21146), .CD(n_62453), .Q(sav_ecx
		[19]));
	notech_mux2 i_2594(.S(n_58832), .A(ecx[19]), .B(sav_ecx[19]), .Z(n_21146
		));
	notech_or2 i_132(.A(n_302260651), .B(n_33150), .Z(n_2865));
	notech_reg sav_ecx_reg_20(.CP(n_63524), .D(n_21152), .CD(n_62452), .Q(sav_ecx
		[20]));
	notech_mux2 i_2602(.S(n_58832), .A(ecx[20]), .B(sav_ecx[20]), .Z(n_21152
		));
	notech_nand3 i_133(.A(n_304060669), .B(n_1816), .C(instrc[49]), .Z(n_2864
		));
	notech_reg sav_ecx_reg_21(.CP(n_63524), .D(n_21158), .CD(n_62452), .Q(sav_ecx
		[21]));
	notech_mux2 i_2610(.S(n_58832), .A(ecx[21]), .B(sav_ecx[21]), .Z(n_21158
		));
	notech_reg sav_ecx_reg_22(.CP(n_63524), .D(n_21164), .CD(n_62452), .Q(sav_ecx
		[22]));
	notech_mux2 i_2618(.S(n_58832), .A(ecx[22]), .B(sav_ecx[22]), .Z(n_21164
		));
	notech_reg sav_ecx_reg_23(.CP(n_63524), .D(n_21170), .CD(n_62449), .Q(sav_ecx
		[23]));
	notech_mux2 i_2626(.S(n_58835), .A(ecx[23]), .B(sav_ecx[23]), .Z(n_21170
		));
	notech_reg sav_ecx_reg_24(.CP(n_63524), .D(n_21176), .CD(n_62449), .Q(sav_ecx
		[24]));
	notech_mux2 i_2634(.S(n_58835), .A(ecx[24]), .B(sav_ecx[24]), .Z(n_21176
		));
	notech_reg sav_ecx_reg_25(.CP(n_63524), .D(n_21182), .CD(n_62449), .Q(sav_ecx
		[25]));
	notech_mux2 i_2642(.S(n_58835), .A(ecx[25]), .B(sav_ecx[25]), .Z(n_21182
		));
	notech_reg sav_ecx_reg_26(.CP(n_63524), .D(n_21188), .CD(n_62449), .Q(sav_ecx
		[26]));
	notech_mux2 i_2650(.S(n_58835), .A(ecx[26]), .B(sav_ecx[26]), .Z(n_21188
		));
	notech_reg sav_ecx_reg_27(.CP(n_63524), .D(n_21194), .CD(n_62452), .Q(sav_ecx
		[27]));
	notech_mux2 i_2658(.S(n_58835), .A(ecx[27]), .B(sav_ecx[27]), .Z(n_21194
		));
	notech_reg sav_ecx_reg_28(.CP(n_63524), .D(n_21200), .CD(n_62452), .Q(sav_ecx
		[28]));
	notech_mux2 i_2666(.S(n_58835), .A(ecx[28]), .B(sav_ecx[28]), .Z(n_21200
		));
	notech_reg sav_ecx_reg_29(.CP(n_63524), .D(n_21206), .CD(n_62452), .Q(sav_ecx
		[29]));
	notech_mux2 i_2674(.S(n_58835), .A(ecx[29]), .B(sav_ecx[29]), .Z(n_21206
		));
	notech_reg sav_ecx_reg_30(.CP(n_63524), .D(n_21212), .CD(n_62452), .Q(sav_ecx
		[30]));
	notech_mux2 i_2682(.S(n_58835), .A(ecx[30]), .B(sav_ecx[30]), .Z(n_21212
		));
	notech_reg sav_ecx_reg_31(.CP(n_63524), .D(n_21218), .CD(n_62452), .Q(sav_ecx
		[31]));
	notech_mux2 i_2690(.S(n_58835), .A(ecx[31]), .B(sav_ecx[31]), .Z(n_21218
		));
	notech_nao3 i_114(.A(n_303060659), .B(n_61964), .C(n_303260661), .Z(n_2853
		));
	notech_reg fesp_reg(.CP(n_63524), .D(n_21224), .CD(n_62446), .Q(fesp));
	notech_mux2 i_2698(.S(n_8555), .A(fesp), .B(n_315692475), .Z(n_21224));
	notech_ao3 i_87(.A(n_1817), .B(n_23350), .C(n_1806), .Z(n_2852));
	notech_reg_set sav_esp_reg_0(.CP(n_63524), .D(n_21230), .SD(1'b1), .Q(sav_esp
		[0]));
	notech_mux2 i_2706(.S(n_348389365), .A(regs_4[0]), .B(sav_esp[0]), .Z(n_21230
		));
	notech_reg_set sav_esp_reg_1(.CP(n_63524), .D(n_21236), .SD(1'b1), .Q(sav_esp
		[1]));
	notech_mux2 i_2714(.S(n_348389365), .A(regs_4[1]), .B(sav_esp[1]), .Z(n_21236
		));
	notech_nand3 i_203137445(.A(n_61094), .B(n_61616), .C(n_30714), .Z(n_35412112
		));
	notech_reg_set sav_esp_reg_2(.CP(n_63524), .D(n_21242), .SD(1'b1), .Q(sav_esp
		[2]));
	notech_mux2 i_2722(.S(n_348389365), .A(regs_4[2]), .B(sav_esp[2]), .Z(n_21242
		));
	notech_ao4 i_30837611(.A(n_2848), .B(n_57633), .C(n_32308), .D(n_32215),
		 .Z(n_2850));
	notech_reg_set sav_esp_reg_3(.CP(n_63524), .D(n_21248), .SD(1'b1), .Q(sav_esp
		[3]));
	notech_mux2 i_2730(.S(n_348389365), .A(regs_4[3]), .B(sav_esp[3]), .Z(n_21248
		));
	notech_reg_set sav_esp_reg_4(.CP(n_63524), .D(n_21254), .SD(1'b1), .Q(sav_esp
		[4]));
	notech_mux2 i_2738(.S(n_348389365), .A(regs_4[4]), .B(sav_esp[4]), .Z(n_21254
		));
	notech_nand3 i_185937467(.A(n_61819), .B(n_32315), .C(n_61092), .Z(n_2848
		));
	notech_reg_set sav_esp_reg_5(.CP(n_63462), .D(n_21260), .SD(1'b1), .Q(sav_esp
		[5]));
	notech_mux2 i_2746(.S(n_348389365), .A(regs_4[5]), .B(sav_esp[5]), .Z(n_21260
		));
	notech_reg_set sav_esp_reg_6(.CP(n_63462), .D(n_21266), .SD(1'b1), .Q(sav_esp
		[6]));
	notech_mux2 i_2754(.S(n_348389365), .A(regs_4[6]), .B(sav_esp[6]), .Z(n_21266
		));
	notech_reg_set sav_esp_reg_7(.CP(n_63462), .D(n_21272), .SD(1'b1), .Q(sav_esp
		[7]));
	notech_mux2 i_2762(.S(n_348389365), .A(regs_4[7]), .B(sav_esp[7]), .Z(n_21272
		));
	notech_nand2 i_96737507(.A(instrc[112]), .B(n_32158), .Z(n_2845));
	notech_reg_set sav_esp_reg_8(.CP(n_63462), .D(n_21278), .SD(1'b1), .Q(sav_esp
		[8]));
	notech_mux2 i_2770(.S(n_348389365), .A(regs_4[8]), .B(sav_esp[8]), .Z(n_21278
		));
	notech_ao4 i_132236354(.A(n_32273), .B(n_275660605), .C(n_60188), .D(n_30788
		), .Z(n_2844));
	notech_reg_set sav_esp_reg_9(.CP(n_63462), .D(n_21284), .SD(1'b1), .Q(sav_esp
		[9]));
	notech_mux2 i_2778(.S(n_348389365), .A(regs_4[9]), .B(sav_esp[9]), .Z(n_21284
		));
	notech_reg_set sav_esp_reg_10(.CP(n_63462), .D(n_21290), .SD(1'b1), .Q(sav_esp
		[10]));
	notech_mux2 i_2786(.S(n_348389365), .A(regs_4[10]), .B(sav_esp[10]), .Z(n_21290
		));
	notech_and4 i_12037556(.A(n_312460752), .B(n_309860726), .C(n_61819), .D
		(n_32583), .Z(n_63212389));
	notech_reg_set sav_esp_reg_11(.CP(n_63462), .D(n_21296), .SD(1'b1), .Q(sav_esp
		[11]));
	notech_mux2 i_2794(.S(n_348389365), .A(regs_4[11]), .B(sav_esp[11]), .Z(n_21296
		));
	notech_reg_set sav_esp_reg_12(.CP(n_63462), .D(n_21302), .SD(1'b1), .Q(sav_esp
		[12]));
	notech_mux2 i_2802(.S(n_348389365), .A(regs_4[12]), .B(sav_esp[12]), .Z(n_21302
		));
	notech_reg_set sav_esp_reg_13(.CP(n_63462), .D(n_21309), .SD(1'b1), .Q(sav_esp
		[13]));
	notech_mux2 i_2810(.S(n_348389365), .A(regs_4[13]), .B(sav_esp[13]), .Z(n_21309
		));
	notech_reg_set sav_esp_reg_14(.CP(n_63462), .D(n_21316), .SD(1'b1), .Q(sav_esp
		[14]));
	notech_mux2 i_2818(.S(n_348389365), .A(regs_4[14]), .B(sav_esp[14]), .Z(n_21316
		));
	notech_mux2 i_76337562(.S(n_2819), .A(n_2770), .B(n_72112478), .Z(n_72012477
		));
	notech_reg_set sav_esp_reg_15(.CP(n_63522), .D(n_21324), .SD(1'b1), .Q(sav_esp
		[15]));
	notech_mux2 i_2826(.S(n_348389365), .A(regs_4[15]), .B(sav_esp[15]), .Z(n_21324
		));
	notech_nand3 i_2130556(.A(n_58696), .B(n_2835), .C(n_2793), .Z(n_72112478
		));
	notech_reg_set sav_esp_reg_16(.CP(n_63516), .D(n_21331), .SD(1'b1), .Q(sav_esp
		[16]));
	notech_mux2 i_2834(.S(n_55568), .A(regs_4[16]), .B(sav_esp[16]), .Z(n_21331
		));
	notech_reg_set sav_esp_reg_17(.CP(n_63460), .D(n_21339), .SD(1'b1), .Q(sav_esp
		[17]));
	notech_mux2 i_2842(.S(n_55568), .A(regs_4[17]), .B(sav_esp[17]), .Z(n_21339
		));
	notech_reg_set sav_esp_reg_18(.CP(n_63516), .D(n_21346), .SD(1'b1), .Q(sav_esp
		[18]));
	notech_mux2 i_2851(.S(n_55568), .A(regs_4[18]), .B(sav_esp[18]), .Z(n_21346
		));
	notech_reg_set sav_esp_reg_19(.CP(n_63516), .D(n_21354), .SD(1'b1), .Q(sav_esp
		[19]));
	notech_mux2 i_2859(.S(n_55568), .A(regs_4[19]), .B(sav_esp[19]), .Z(n_21354
		));
	notech_ao4 i_137236305(.A(n_60440), .B(n_2815), .C(n_31369), .D(n_2789),
		 .Z(n_2836));
	notech_reg_set sav_esp_reg_20(.CP(n_63516), .D(n_21361), .SD(1'b1), .Q(sav_esp
		[20]));
	notech_mux2 i_2868(.S(n_55568), .A(regs_4[20]), .B(sav_esp[20]), .Z(n_21361
		));
	notech_ao4 i_136936308(.A(n_2787), .B(n_31372), .C(n_58707), .D(n_2786),
		 .Z(n_2835));
	notech_reg_set sav_esp_reg_21(.CP(n_63516), .D(n_21369), .SD(1'b1), .Q(sav_esp
		[21]));
	notech_mux2 i_2876(.S(n_55568), .A(regs_4[21]), .B(sav_esp[21]), .Z(n_21369
		));
	notech_reg_set sav_esp_reg_22(.CP(n_63516), .D(n_21376), .SD(1'b1), .Q(sav_esp
		[22]));
	notech_mux2 i_2884(.S(n_55568), .A(regs_4[22]), .B(sav_esp[22]), .Z(n_21376
		));
	notech_ao4 i_137536302(.A(n_2823), .B(n_2789), .C(n_60440), .D(n_2815), 
		.Z(n_2833));
	notech_reg_set sav_esp_reg_23(.CP(n_63516), .D(n_21384), .SD(1'b1), .Q(sav_esp
		[23]));
	notech_mux2 i_2892(.S(n_55568), .A(regs_4[23]), .B(sav_esp[23]), .Z(n_21384
		));
	notech_reg_set sav_esp_reg_24(.CP(n_63516), .D(n_21391), .SD(1'b1), .Q(sav_esp
		[24]));
	notech_mux2 i_2900(.S(n_55568), .A(regs_4[24]), .B(sav_esp[24]), .Z(n_21391
		));
	notech_ao4 i_137736300(.A(n_60431), .B(n_31370), .C(n_60440), .D(n_31371
		), .Z(n_2831));
	notech_reg_set sav_esp_reg_25(.CP(n_63516), .D(n_21399), .SD(1'b1), .Q(sav_esp
		[25]));
	notech_mux2 i_2908(.S(n_55568), .A(regs_4[25]), .B(sav_esp[25]), .Z(n_21399
		));
	notech_or2 i_207837442(.A(n_60422), .B(instrc[115]), .Z(n_2830));
	notech_reg_set sav_esp_reg_26(.CP(n_63516), .D(n_21406), .SD(1'b1), .Q(sav_esp
		[26]));
	notech_mux2 i_2916(.S(n_55568), .A(regs_4[26]), .B(sav_esp[26]), .Z(n_21406
		));
	notech_or2 i_90537508(.A(instrc[113]), .B(n_32157), .Z(n_2829));
	notech_reg_set sav_esp_reg_27(.CP(n_63516), .D(n_21414), .SD(1'b1), .Q(sav_esp
		[27]));
	notech_mux2 i_2924(.S(n_55568), .A(regs_4[27]), .B(sav_esp[27]), .Z(n_21414
		));
	notech_reg_set sav_esp_reg_28(.CP(n_63602), .D(n_21421), .SD(1'b1), .Q(sav_esp
		[28]));
	notech_mux2 i_2932(.S(n_55568), .A(regs_4[28]), .B(sav_esp[28]), .Z(n_21421
		));
	notech_ao4 i_138036298(.A(all_cnt[3]), .B(n_2822), .C(n_2778), .D(n_2826
		), .Z(n_2827));
	notech_reg_set sav_esp_reg_29(.CP(n_63602), .D(n_21429), .SD(1'b1), .Q(sav_esp
		[29]));
	notech_mux2 i_2940(.S(n_55568), .A(regs_4[29]), .B(sav_esp[29]), .Z(n_21429
		));
	notech_or2 i_138136297(.A(all_cnt[2]), .B(n_2825), .Z(n_2826));
	notech_reg_set sav_esp_reg_30(.CP(n_63602), .D(n_21436), .SD(1'b1), .Q(sav_esp
		[30]));
	notech_mux2 i_2948(.S(n_55568), .A(regs_4[30]), .B(sav_esp[30]), .Z(n_21436
		));
	notech_ao4 i_101337505(.A(all_cnt[1]), .B(n_31000), .C(n_60440), .D(n_2824
		), .Z(n_2825));
	notech_reg_set sav_esp_reg_31(.CP(n_63602), .D(n_21444), .SD(1'b1), .Q(sav_esp
		[31]));
	notech_mux2 i_2956(.S(n_55568), .A(regs_4[31]), .B(sav_esp[31]), .Z(n_21444
		));
	notech_and2 i_3737430(.A(all_cnt[1]), .B(n_31000), .Z(n_2824));
	notech_reg sav_esi_reg_0(.CP(n_63602), .D(n_21451), .CD(n_62446), .Q(sav_esi
		[0]));
	notech_mux2 i_2964(.S(n_58835), .A(regs_6[0]), .B(sav_esi[0]), .Z(n_21451
		));
	notech_and2 i_96837510(.A(n_60422), .B(n_31369), .Z(n_2823));
	notech_reg sav_esi_reg_1(.CP(n_63602), .D(n_21459), .CD(n_62446), .Q(sav_esi
		[1]));
	notech_mux2 i_2972(.S(n_58835), .A(regs_6[1]), .B(sav_esi[1]), .Z(n_21459
		));
	notech_xor2 i_52044(.A(instrc[115]), .B(n_2820), .Z(n_2822));
	notech_reg sav_esi_reg_2(.CP(n_63602), .D(n_21466), .CD(n_62446), .Q(sav_esi
		[2]));
	notech_mux2 i_2980(.S(n_58835), .A(regs_6[2]), .B(sav_esi[2]), .Z(n_21466
		));
	notech_nand3 i_102537504(.A(n_60440), .B(n_60431), .C(instrc[115]), .Z(n_2821
		));
	notech_reg sav_esi_reg_3(.CP(n_63602), .D(n_21472), .CD(n_62446), .Q(sav_esi
		[3]));
	notech_mux2 i_2988(.S(n_58833), .A(regs_6[3]), .B(sav_esi[3]), .Z(n_21472
		));
	notech_nand2 i_88137509(.A(n_60440), .B(n_60431), .Z(n_2820));
	notech_reg sav_esi_reg_4(.CP(n_63602), .D(n_21478), .CD(n_62446), .Q(sav_esi
		[4]));
	notech_mux2 i_2996(.S(n_58833), .A(regs_6[4]), .B(sav_esi[4]), .Z(n_21478
		));
	notech_and2 i_530744(.A(n_275860607), .B(n_275760606), .Z(n_2819));
	notech_reg sav_esi_reg_5(.CP(n_63602), .D(n_21484), .CD(n_62446), .Q(sav_esi
		[5]));
	notech_mux2 i_3004(.S(n_58833), .A(regs_6[5]), .B(sav_esi[5]), .Z(n_21484
		));
	notech_or4 i_3943(.A(all_cnt[3]), .B(n_31369), .C(all_cnt[1]), .D(all_cnt
		[2]), .Z(n_75912515));
	notech_reg sav_esi_reg_6(.CP(n_63602), .D(n_21490), .CD(n_62446), .Q(sav_esi
		[6]));
	notech_mux2 i_3012(.S(n_58833), .A(regs_6[6]), .B(sav_esi[6]), .Z(n_21490
		));
	notech_or4 i_8637412(.A(all_cnt[0]), .B(all_cnt[3]), .C(all_cnt[1]), .D(all_cnt
		[2]), .Z(n_76412520));
	notech_reg sav_esi_reg_7(.CP(n_63602), .D(n_21496), .CD(n_62446), .Q(sav_esi
		[7]));
	notech_mux2 i_3020(.S(n_58833), .A(regs_6[7]), .B(sav_esi[7]), .Z(n_21496
		));
	notech_reg sav_esi_reg_8(.CP(n_63602), .D(n_21502), .CD(n_62446), .Q(sav_esi
		[8]));
	notech_mux2 i_3028(.S(n_58833), .A(regs_6[8]), .B(sav_esi[8]), .Z(n_21502
		));
	notech_or4 i_189237462(.A(n_61717), .B(n_61880), .C(n_61864), .D(tcmp), 
		.Z(n_76712523));
	notech_reg sav_esi_reg_9(.CP(n_63602), .D(n_21508), .CD(n_62444), .Q(sav_esi
		[9]));
	notech_mux2 i_3036(.S(n_58833), .A(regs_6[9]), .B(sav_esi[9]), .Z(n_21508
		));
	notech_ao4 i_141036274(.A(n_331960947), .B(n_30287), .C(n_335660984), .D
		(n_57656), .Z(n_2817));
	notech_reg sav_esi_reg_10(.CP(n_63602), .D(n_21514), .CD(n_62444), .Q(sav_esi
		[10]));
	notech_mux2 i_3044(.S(n_58835), .A(regs_6[10]), .B(sav_esi[10]), .Z(n_21514
		));
	notech_or4 i_3950(.A(all_cnt[2]), .B(n_31370), .C(all_cnt[3]), .D(n_31369
		), .Z(n_77012526));
	notech_reg sav_esi_reg_11(.CP(n_63602), .D(n_21520), .CD(n_62444), .Q(sav_esi
		[11]));
	notech_mux2 i_3052(.S(n_58835), .A(regs_6[11]), .B(sav_esi[11]), .Z(n_21520
		));
	notech_reg sav_esi_reg_12(.CP(n_63602), .D(n_21526), .CD(n_62444), .Q(sav_esi
		[12]));
	notech_mux2 i_3060(.S(n_58833), .A(regs_6[12]), .B(sav_esi[12]), .Z(n_21526
		));
	notech_or4 i_3960(.A(n_31370), .B(n_31371), .C(all_cnt[0]), .D(all_cnt[3
		]), .Z(n_77712533));
	notech_reg sav_esi_reg_13(.CP(n_63602), .D(n_21532), .CD(n_62444), .Q(sav_esi
		[13]));
	notech_mux2 i_3068(.S(n_58833), .A(regs_6[13]), .B(sav_esi[13]), .Z(n_21532
		));
	notech_nand2 i_191237460(.A(n_33155), .B(n_33141), .Z(n_77812534));
	notech_reg sav_esi_reg_14(.CP(n_63602), .D(n_21538), .CD(n_62444), .Q(sav_esi
		[14]));
	notech_mux2 i_3076(.S(n_58833), .A(regs_6[14]), .B(sav_esi[14]), .Z(n_21538
		));
	notech_reg sav_esi_reg_15(.CP(n_63666), .D(n_21544), .CD(n_62444), .Q(sav_esi
		[15]));
	notech_mux2 i_3084(.S(n_58827), .A(regs_6[15]), .B(sav_esi[15]), .Z(n_21544
		));
	notech_nand2 i_170237473(.A(all_cnt[1]), .B(all_cnt[2]), .Z(n_2815));
	notech_reg sav_esi_reg_16(.CP(n_63600), .D(n_21550), .CD(n_62444), .Q(sav_esi
		[16]));
	notech_mux2 i_3092(.S(n_58820), .A(regs_6[16]), .B(sav_esi[16]), .Z(n_21550
		));
	notech_nand2 i_191337459(.A(n_33154), .B(n_33138), .Z(n_78212538));
	notech_reg sav_esi_reg_17(.CP(n_63666), .D(n_21556), .CD(n_62444), .Q(sav_esi
		[17]));
	notech_mux2 i_3100(.S(n_58820), .A(regs_6[17]), .B(sav_esi[17]), .Z(n_21556
		));
	notech_and4 i_3957(.A(n_31372), .B(all_cnt[0]), .C(n_31370), .D(all_cnt[
		2]), .Z(n_78412540));
	notech_reg sav_esi_reg_18(.CP(n_63666), .D(n_21562), .CD(n_62447), .Q(sav_esi
		[18]));
	notech_mux2 i_3108(.S(n_58820), .A(regs_6[18]), .B(sav_esi[18]), .Z(n_21562
		));
	notech_and2 i_154737482(.A(n_31372), .B(all_cnt[0]), .Z(n_2814));
	notech_reg sav_esi_reg_19(.CP(n_63666), .D(n_21568), .CD(n_62447), .Q(sav_esi
		[19]));
	notech_mux2 i_3116(.S(n_58820), .A(regs_6[19]), .B(sav_esi[19]), .Z(n_21568
		));
	notech_reg sav_esi_reg_20(.CP(n_63666), .D(n_21574), .CD(n_62447), .Q(sav_esi
		[20]));
	notech_mux2 i_3124(.S(n_58820), .A(regs_6[20]), .B(sav_esi[20]), .Z(n_21574
		));
	notech_nand2 i_207737443(.A(n_31370), .B(all_cnt[2]), .Z(n_79512551));
	notech_reg sav_esi_reg_21(.CP(n_63666), .D(n_21580), .CD(n_62447), .Q(sav_esi
		[21]));
	notech_mux2 i_3132(.S(n_58820), .A(regs_6[21]), .B(sav_esi[21]), .Z(n_21580
		));
	notech_reg sav_esi_reg_22(.CP(n_63666), .D(n_21586), .CD(n_62447), .Q(sav_esi
		[22]));
	notech_mux2 i_3140(.S(n_58833), .A(regs_6[22]), .B(sav_esi[22]), .Z(n_21586
		));
	notech_reg sav_esi_reg_23(.CP(n_63666), .D(n_21592), .CD(n_62448), .Q(sav_esi
		[23]));
	notech_mux2 i_3148(.S(n_58833), .A(regs_6[23]), .B(sav_esi[23]), .Z(n_21592
		));
	notech_reg sav_esi_reg_24(.CP(n_63666), .D(n_21598), .CD(n_62448), .Q(sav_esi
		[24]));
	notech_mux2 i_3156(.S(n_58833), .A(regs_6[24]), .B(sav_esi[24]), .Z(n_21598
		));
	notech_nand2 i_7637422(.A(n_31371), .B(all_cnt[1]), .Z(n_80312559));
	notech_reg sav_esi_reg_25(.CP(n_63666), .D(n_21604), .CD(n_62447), .Q(sav_esi
		[25]));
	notech_mux2 i_3164(.S(n_58833), .A(regs_6[25]), .B(sav_esi[25]), .Z(n_21604
		));
	notech_nand2 i_154937481(.A(n_31369), .B(n_31372), .Z(n_80512561));
	notech_reg sav_esi_reg_26(.CP(n_63666), .D(n_21610), .CD(n_62448), .Q(sav_esi
		[26]));
	notech_mux2 i_3172(.S(n_58833), .A(regs_6[26]), .B(sav_esi[26]), .Z(n_21610
		));
	notech_nao3 i_58537534(.A(n_61819), .B(n_31249), .C(n_30804), .Z(n_2810)
		);
	notech_reg sav_esi_reg_27(.CP(n_63666), .D(n_21616), .CD(n_62447), .Q(sav_esi
		[27]));
	notech_mux2 i_3180(.S(n_58833), .A(regs_6[27]), .B(sav_esi[27]), .Z(n_21616
		));
	notech_reg sav_esi_reg_28(.CP(n_63666), .D(n_21622), .CD(n_62446), .Q(sav_esi
		[28]));
	notech_mux2 i_3188(.S(n_58820), .A(regs_6[28]), .B(sav_esi[28]), .Z(n_21622
		));
	notech_reg sav_esi_reg_29(.CP(n_63666), .D(n_21628), .CD(n_62447), .Q(sav_esi
		[29]));
	notech_mux2 i_3196(.S(n_58820), .A(regs_6[29]), .B(sav_esi[29]), .Z(n_21628
		));
	notech_reg sav_esi_reg_30(.CP(n_63666), .D(n_21634), .CD(n_62446), .Q(sav_esi
		[30]));
	notech_mux2 i_3204(.S(n_58820), .A(regs_6[30]), .B(sav_esi[30]), .Z(n_21634
		));
	notech_reg sav_esi_reg_31(.CP(n_63666), .D(n_21640), .CD(n_62446), .Q(sav_esi
		[31]));
	notech_mux2 i_3212(.S(n_58820), .A(regs_6[31]), .B(sav_esi[31]), .Z(n_21640
		));
	notech_or2 i_184660736(.A(n_335660984), .B(n_57656), .Z(n_2805));
	notech_reg sav_edi_reg_0(.CP(n_63666), .D(n_21646), .CD(n_62447), .Q(sav_edi
		[0]));
	notech_mux2 i_3220(.S(n_58820), .A(regs_7[0]), .B(sav_edi[0]), .Z(n_21646
		));
	notech_reg sav_edi_reg_1(.CP(n_63666), .D(n_21652), .CD(n_62447), .Q(sav_edi
		[1]));
	notech_mux2 i_3228(.S(n_58820), .A(regs_7[1]), .B(sav_edi[1]), .Z(n_21652
		));
	notech_reg sav_edi_reg_2(.CP(n_63666), .D(n_21658), .CD(n_62447), .Q(sav_edi
		[2]));
	notech_mux2 i_3236(.S(n_58820), .A(regs_7[2]), .B(sav_edi[2]), .Z(n_21658
		));
	notech_reg sav_edi_reg_3(.CP(n_63600), .D(n_21664), .CD(n_62447), .Q(sav_edi
		[3]));
	notech_mux2 i_3244(.S(n_58820), .A(regs_7[3]), .B(sav_edi[3]), .Z(n_21664
		));
	notech_reg sav_edi_reg_4(.CP(n_63600), .D(n_21670), .CD(n_62447), .Q(sav_edi
		[4]));
	notech_mux2 i_3252(.S(n_58820), .A(regs_7[4]), .B(sav_edi[4]), .Z(n_21670
		));
	notech_reg sav_edi_reg_5(.CP(n_63600), .D(n_21676), .CD(n_62424), .Q(sav_edi
		[5]));
	notech_mux2 i_3260(.S(n_58820), .A(regs_7[5]), .B(sav_edi[5]), .Z(n_21676
		));
	notech_or2 i_67536914(.A(n_340361031), .B(n_31370), .Z(n_2799));
	notech_reg sav_edi_reg_6(.CP(n_63600), .D(n_21682), .CD(n_62424), .Q(sav_edi
		[6]));
	notech_mux2 i_3268(.S(n_58820), .A(regs_7[6]), .B(sav_edi[6]), .Z(n_21682
		));
	notech_reg sav_edi_reg_7(.CP(n_63600), .D(n_21688), .CD(n_62424), .Q(sav_edi
		[7]));
	notech_mux2 i_3276(.S(n_58820), .A(regs_7[7]), .B(sav_edi[7]), .Z(n_21688
		));
	notech_reg sav_edi_reg_8(.CP(n_63600), .D(n_21694), .CD(n_62424), .Q(sav_edi
		[8]));
	notech_mux2 i_3284(.S(n_58827), .A(regs_7[8]), .B(sav_edi[8]), .Z(n_21694
		));
	notech_or2 i_67636913(.A(n_60431), .B(n_31371), .Z(n_2796));
	notech_reg sav_edi_reg_9(.CP(n_63600), .D(n_21700), .CD(n_62424), .Q(sav_edi
		[9]));
	notech_mux2 i_3292(.S(n_58827), .A(regs_7[9]), .B(sav_edi[9]), .Z(n_21700
		));
	notech_reg sav_edi_reg_10(.CP(n_63600), .D(n_21706), .CD(n_62424), .Q(sav_edi
		[10]));
	notech_mux2 i_3300(.S(n_58827), .A(regs_7[10]), .B(sav_edi[10]), .Z(n_21706
		));
	notech_reg sav_edi_reg_11(.CP(n_63600), .D(n_21712), .CD(n_62424), .Q(sav_edi
		[11]));
	notech_mux2 i_3308(.S(n_58827), .A(regs_7[11]), .B(sav_edi[11]), .Z(n_21712
		));
	notech_or2 i_66636923(.A(instrc[115]), .B(n_2788), .Z(n_2793));
	notech_reg sav_edi_reg_12(.CP(n_63600), .D(n_21718), .CD(n_62424), .Q(sav_edi
		[12]));
	notech_mux2 i_3316(.S(n_58827), .A(regs_7[12]), .B(sav_edi[12]), .Z(n_21718
		));
	notech_or4 i_27084(.A(n_61880), .B(n_339461022), .C(n_61717), .D(\opcode[3] 
		), .Z(n_32314));
	notech_reg sav_edi_reg_13(.CP(n_63600), .D(n_21724), .CD(n_62424), .Q(sav_edi
		[13]));
	notech_mux2 i_3324(.S(n_58827), .A(regs_7[13]), .B(sav_edi[13]), .Z(n_21724
		));
	notech_reg sav_edi_reg_14(.CP(n_63516), .D(n_21730), .CD(n_62423), .Q(sav_edi
		[14]));
	notech_mux2 i_3332(.S(n_58827), .A(regs_7[14]), .B(sav_edi[14]), .Z(n_21730
		));
	notech_ao3 i_27088(.A(n_61661), .B(\opcode[3] ), .C(n_339461022), .Z(n_32310
		));
	notech_reg sav_edi_reg_15(.CP(n_63460), .D(n_21736), .CD(n_62423), .Q(sav_edi
		[15]));
	notech_mux2 i_3340(.S(n_58827), .A(regs_7[15]), .B(sav_edi[15]), .Z(n_21736
		));
	notech_reg sav_edi_reg_16(.CP(n_63604), .D(n_21742), .CD(n_62423), .Q(sav_edi
		[16]));
	notech_mux2 i_3348(.S(n_58827), .A(regs_7[16]), .B(sav_edi[16]), .Z(n_21742
		));
	notech_or2 i_35887(.A(n_390464435), .B(n_23763), .Z(n_23511));
	notech_reg sav_edi_reg_17(.CP(n_63518), .D(n_21748), .CD(n_62423), .Q(sav_edi
		[17]));
	notech_mux2 i_3356(.S(n_58827), .A(regs_7[17]), .B(sav_edi[17]), .Z(n_21748
		));
	notech_or2 i_35888(.A(n_334560973), .B(n_23763), .Z(n_23510));
	notech_reg sav_edi_reg_18(.CP(n_63518), .D(n_21754), .CD(n_62423), .Q(sav_edi
		[18]));
	notech_mux2 i_3364(.S(n_58827), .A(regs_7[18]), .B(sav_edi[18]), .Z(n_21754
		));
	notech_reg sav_edi_reg_19(.CP(n_63518), .D(n_21760), .CD(n_62423), .Q(sav_edi
		[19]));
	notech_mux2 i_3372(.S(n_58827), .A(regs_7[19]), .B(sav_edi[19]), .Z(n_21760
		));
	notech_reg sav_edi_reg_20(.CP(n_63518), .D(n_21766), .CD(n_62423), .Q(sav_edi
		[20]));
	notech_mux2 i_3380(.S(n_58832), .A(regs_7[20]), .B(sav_edi[20]), .Z(n_21766
		));
	notech_and3 i_19337333(.A(n_340361031), .B(n_2815), .C(n_2831), .Z(n_2789
		));
	notech_reg sav_edi_reg_21(.CP(n_63518), .D(n_21772), .CD(n_62423), .Q(sav_edi
		[21]));
	notech_mux2 i_3388(.S(n_58832), .A(regs_7[21]), .B(sav_edi[21]), .Z(n_21772
		));
	notech_and4 i_19237334(.A(n_2796), .B(n_2799), .C(n_2836), .D(n_31372), 
		.Z(n_2788));
	notech_reg sav_edi_reg_22(.CP(n_63518), .D(n_21778), .CD(n_62423), .Q(sav_edi
		[22]));
	notech_mux2 i_3396(.S(n_58832), .A(regs_7[22]), .B(sav_edi[22]), .Z(n_21778
		));
	notech_and3 i_19137335(.A(n_2833), .B(n_2799), .C(n_2796), .Z(n_2787));
	notech_reg sav_edi_reg_23(.CP(n_63518), .D(n_21784), .CD(n_62423), .Q(sav_edi
		[23]));
	notech_mux2 i_3404(.S(n_58832), .A(regs_7[23]), .B(sav_edi[23]), .Z(n_21784
		));
	notech_and2 i_19037336(.A(n_2815), .B(n_2831), .Z(n_2786));
	notech_reg sav_edi_reg_24(.CP(n_63518), .D(n_21790), .CD(n_62425), .Q(sav_edi
		[24]));
	notech_mux2 i_3412(.S(n_58832), .A(regs_7[24]), .B(sav_edi[24]), .Z(n_21790
		));
	notech_reg sav_edi_reg_25(.CP(n_63518), .D(n_21796), .CD(n_62425), .Q(sav_edi
		[25]));
	notech_mux2 i_3420(.S(n_58832), .A(regs_7[25]), .B(sav_edi[25]), .Z(n_21796
		));
	notech_reg sav_edi_reg_26(.CP(n_63518), .D(n_21802), .CD(n_62425), .Q(sav_edi
		[26]));
	notech_mux2 i_3428(.S(n_58835), .A(regs_7[26]), .B(sav_edi[26]), .Z(n_21802
		));
	notech_reg sav_edi_reg_27(.CP(n_63604), .D(n_21808), .CD(n_62425), .Q(sav_edi
		[27]));
	notech_mux2 i_3436(.S(n_58835), .A(regs_7[27]), .B(sav_edi[27]), .Z(n_21808
		));
	notech_reg sav_edi_reg_28(.CP(n_63604), .D(n_21814), .CD(n_62425), .Q(sav_edi
		[28]));
	notech_mux2 i_3444(.S(n_58835), .A(regs_7[28]), .B(sav_edi[28]), .Z(n_21814
		));
	notech_reg sav_edi_reg_29(.CP(n_63604), .D(n_21820), .CD(n_62426), .Q(sav_edi
		[29]));
	notech_mux2 i_3452(.S(n_58835), .A(regs_7[29]), .B(sav_edi[29]), .Z(n_21820
		));
	notech_reg sav_edi_reg_30(.CP(n_63604), .D(n_21826), .CD(n_62426), .Q(sav_edi
		[30]));
	notech_mux2 i_3460(.S(n_58835), .A(regs_7[30]), .B(sav_edi[30]), .Z(n_21826
		));
	notech_reg sav_edi_reg_31(.CP(n_63604), .D(n_21832), .CD(n_62425), .Q(sav_edi
		[31]));
	notech_mux2 i_3468(.S(n_58835), .A(regs_7[31]), .B(sav_edi[31]), .Z(n_21832
		));
	notech_and2 i_7737421(.A(n_2822), .B(all_cnt[3]), .Z(n_2778));
	notech_reg fepc_reg(.CP(n_63604), .D(n_21838), .CD(n_62425), .Q(fepc));
	notech_mux2 i_3476(.S(n_10020), .A(fepc), .B(n_10023), .Z(n_21838));
	notech_and3 i_14437356(.A(n_31000), .B(all_cnt[1]), .C(all_cnt[2]), .Z(n_2777
		));
	notech_reg_set sav_epc_reg_0(.CP(n_63604), .D(n_21844), .SD(1'b1), .Q(sav_epc
		[0]));
	notech_mux2 i_3484(.S(n_30894), .A(sav_epc[0]), .B(regs_14[0]), .Z(n_21844
		));
	notech_reg_set sav_epc_reg_1(.CP(n_63604), .D(n_21850), .SD(1'b1), .Q(sav_epc
		[1]));
	notech_mux2 i_3492(.S(n_30894), .A(sav_epc[1]), .B(regs_14[1]), .Z(n_21850
		));
	notech_and2 i_14337357(.A(all_cnt[2]), .B(n_2825), .Z(n_2775));
	notech_reg_set sav_epc_reg_2(.CP(n_63604), .D(n_21856), .SD(1'b1), .Q(sav_epc
		[2]));
	notech_mux2 i_3500(.S(n_30894), .A(sav_epc[2]), .B(regs_14[2]), .Z(n_21856
		));
	notech_reg_set sav_epc_reg_3(.CP(n_63604), .D(n_21862), .SD(1'b1), .Q(sav_epc
		[3]));
	notech_mux2 i_3508(.S(n_30894), .A(sav_epc[3]), .B(regs_14[3]), .Z(n_21862
		));
	notech_ao4 i_14237358(.A(n_2829), .B(n_2777), .C(n_58716), .D(n_2775), .Z
		(n_2773));
	notech_reg_set sav_epc_reg_4(.CP(n_63604), .D(n_21868), .SD(1'b1), .Q(sav_epc
		[4]));
	notech_mux2 i_3516(.S(n_30894), .A(sav_epc[4]), .B(regs_14[4]), .Z(n_21868
		));
	notech_or2 i_65236937(.A(n_2773), .B(n_2778), .Z(n_2772));
	notech_reg_set sav_epc_reg_5(.CP(n_63604), .D(n_21874), .SD(1'b1), .Q(sav_epc
		[5]));
	notech_mux2 i_3524(.S(n_30894), .A(sav_epc[5]), .B(regs_14[5]), .Z(n_21874
		));
	notech_reg_set sav_epc_reg_6(.CP(n_63604), .D(n_21880), .SD(1'b1), .Q(sav_epc
		[6]));
	notech_mux2 i_3532(.S(n_30894), .A(sav_epc[6]), .B(regs_14[6]), .Z(n_21880
		));
	notech_and3 i_14137359(.A(n_2821), .B(n_2827), .C(n_2772), .Z(n_2770));
	notech_reg_set sav_epc_reg_7(.CP(n_63604), .D(n_21886), .SD(1'b1), .Q(sav_epc
		[7]));
	notech_mux2 i_3540(.S(n_30894), .A(sav_epc[7]), .B(regs_14[7]), .Z(n_21886
		));
	notech_reg_set sav_epc_reg_8(.CP(n_63604), .D(n_21892), .SD(1'b1), .Q(sav_epc
		[8]));
	notech_mux2 i_3548(.S(n_30894), .A(sav_epc[8]), .B(regs_14[8]), .Z(n_21892
		));
	notech_reg_set sav_epc_reg_9(.CP(n_63604), .D(n_21898), .SD(1'b1), .Q(sav_epc
		[9]));
	notech_mux2 i_3556(.S(n_30894), .A(sav_epc[9]), .B(regs_14[9]), .Z(n_21898
		));
	notech_nand2 i_47537086(.A(n_115942600), .B(n_32342), .Z(n_276760616));
	notech_reg_set sav_epc_reg_10(.CP(n_63604), .D(n_21904), .SD(1'b1), .Q(sav_epc
		[10]));
	notech_mux2 i_3564(.S(n_30894), .A(sav_epc[10]), .B(regs_14[10]), .Z(n_21904
		));
	notech_and4 i_46637095(.A(n_32310), .B(n_61092), .C(n_32323), .D(n_57199
		), .Z(n_276660615));
	notech_reg_set sav_epc_reg_11(.CP(n_63604), .D(n_21910), .SD(1'b1), .Q(sav_epc
		[11]));
	notech_mux2 i_3572(.S(n_30894), .A(sav_epc[11]), .B(regs_14[11]), .Z(n_21910
		));
	notech_reg_set sav_epc_reg_12(.CP(n_63518), .D(n_21916), .SD(1'b1), .Q(sav_epc
		[12]));
	notech_mux2 i_3580(.S(n_30894), .A(sav_epc[12]), .B(regs_14[12]), .Z(n_21916
		));
	notech_and4 i_46437097(.A(n_32310), .B(n_61092), .C(n_32321), .D(n_57199
		), .Z(n_276460613));
	notech_reg_set sav_epc_reg_13(.CP(n_63518), .D(n_21922), .SD(1'b1), .Q(sav_epc
		[13]));
	notech_mux2 i_3588(.S(n_30894), .A(sav_epc[13]), .B(regs_14[13]), .Z(n_21922
		));
	notech_reg_set sav_epc_reg_14(.CP(n_63520), .D(n_21928), .SD(1'b1), .Q(sav_epc
		[14]));
	notech_mux2 i_3596(.S(n_30894), .A(sav_epc[14]), .B(regs_14[14]), .Z(n_21928
		));
	notech_reg_set sav_epc_reg_15(.CP(n_63520), .D(n_21934), .SD(1'b1), .Q(sav_epc
		[15]));
	notech_mux2 i_3604(.S(n_30894), .A(sav_epc[15]), .B(regs_14[15]), .Z(n_21934
		));
	notech_reg_set sav_epc_reg_16(.CP(n_63520), .D(n_21940), .SD(1'b1), .Q(sav_epc
		[16]));
	notech_mux2 i_3612(.S(n_55771), .A(sav_epc[16]), .B(regs_14[16]), .Z(n_21940
		));
	notech_reg_set sav_epc_reg_17(.CP(n_63520), .D(n_21946), .SD(1'b1), .Q(sav_epc
		[17]));
	notech_mux2 i_3620(.S(n_55771), .A(sav_epc[17]), .B(regs_14[17]), .Z(n_21946
		));
	notech_reg_set sav_epc_reg_18(.CP(n_63520), .D(n_21952), .SD(1'b1), .Q(sav_epc
		[18]));
	notech_mux2 i_3628(.S(n_55771), .A(sav_epc[18]), .B(regs_14[18]), .Z(n_21952
		));
	notech_xor2 i_21237314(.A(sav_cs[1]), .B(n_31368), .Z(n_275860607));
	notech_reg_set sav_epc_reg_19(.CP(n_63520), .D(n_21958), .SD(1'b1), .Q(sav_epc
		[19]));
	notech_mux2 i_3636(.S(n_55771), .A(sav_epc[19]), .B(regs_14[19]), .Z(n_21958
		));
	notech_xor2 i_21137315(.A(sav_cs[0]), .B(n_31367), .Z(n_275760606));
	notech_reg_set sav_epc_reg_20(.CP(n_63520), .D(n_21964), .SD(1'b1), .Q(sav_epc
		[20]));
	notech_mux2 i_3644(.S(n_55771), .A(sav_epc[20]), .B(regs_14[20]), .Z(n_21964
		));
	notech_ao4 i_124837499(.A(n_63792), .B(n_61958), .C(n_61056), .D(n_30788
		), .Z(n_275660605));
	notech_reg_set sav_epc_reg_21(.CP(n_63520), .D(n_21970), .SD(1'b1), .Q(sav_epc
		[21]));
	notech_mux2 i_3652(.S(n_55771), .A(sav_epc[21]), .B(regs_14[21]), .Z(n_21970
		));
	notech_or4 i_187437466(.A(n_58583), .B(n_61786), .C(n_61766), .D(n_275660605
		), .Z(n_26618));
	notech_reg_set sav_epc_reg_22(.CP(n_63520), .D(n_21976), .SD(1'b1), .Q(sav_epc
		[22]));
	notech_mux2 i_3660(.S(n_55771), .A(sav_epc[22]), .B(regs_14[22]), .Z(n_21976
		));
	notech_and3 i_166637475(.A(n_57705), .B(n_57686), .C(n_33152), .Z(n_275560604
		));
	notech_reg_set sav_epc_reg_23(.CP(n_63520), .D(n_21982), .SD(1'b1), .Q(sav_epc
		[23]));
	notech_mux2 i_3668(.S(n_55771), .A(sav_epc[23]), .B(regs_14[23]), .Z(n_21982
		));
	notech_nor2 i_131037496(.A(n_339461022), .B(n_61616), .Z(n_32315));
	notech_reg_set sav_epc_reg_24(.CP(n_63520), .D(n_21988), .SD(1'b1), .Q(sav_epc
		[24]));
	notech_mux2 i_3676(.S(n_55771), .A(sav_epc[24]), .B(regs_14[24]), .Z(n_21988
		));
	notech_reg_set sav_epc_reg_25(.CP(n_63520), .D(n_21994), .SD(1'b1), .Q(sav_epc
		[25]));
	notech_mux2 i_3684(.S(n_55771), .A(sav_epc[25]), .B(regs_14[25]), .Z(n_21994
		));
	notech_or4 i_22837551(.A(n_61815), .B(n_57535), .C(n_61864), .D(n_57656)
		, .Z(n_32292));
	notech_reg_set sav_epc_reg_26(.CP(n_63520), .D(n_22000), .SD(1'b1), .Q(sav_epc
		[26]));
	notech_mux2 i_3692(.S(n_55771), .A(sav_epc[26]), .B(regs_14[26]), .Z(n_22000
		));
	notech_or4 i_22737552(.A(n_61815), .B(n_57535), .C(n_61864), .D(n_57633)
		, .Z(n_32308));
	notech_reg_set sav_epc_reg_27(.CP(n_63520), .D(n_22006), .SD(1'b1), .Q(sav_epc
		[27]));
	notech_mux2 i_3700(.S(n_55771), .A(sav_epc[27]), .B(regs_14[27]), .Z(n_22006
		));
	notech_or4 i_22637553(.A(n_61815), .B(n_57672), .C(n_57535), .D(n_61864)
		, .Z(n_32288));
	notech_reg_set sav_epc_reg_28(.CP(n_63520), .D(n_22012), .SD(1'b1), .Q(sav_epc
		[28]));
	notech_mux2 i_3708(.S(n_55771), .A(sav_epc[28]), .B(regs_14[28]), .Z(n_22012
		));
	notech_or4 i_22537554(.A(n_61815), .B(n_57535), .C(n_61864), .D(n_57662)
		, .Z(n_32290));
	notech_reg_set sav_epc_reg_29(.CP(n_63520), .D(n_22018), .SD(1'b1), .Q(sav_epc
		[29]));
	notech_mux2 i_3716(.S(n_55771), .A(sav_epc[29]), .B(regs_14[29]), .Z(n_22018
		));
	notech_nand2 i_104937595(.A(n_391064441), .B(n_23759), .Z(n_23615));
	notech_reg_set sav_epc_reg_30(.CP(n_63520), .D(n_22024), .SD(1'b1), .Q(sav_epc
		[30]));
	notech_mux2 i_3724(.S(n_55771), .A(sav_epc[30]), .B(regs_14[30]), .Z(n_22024
		));
	notech_or4 i_10288(.A(instrc[115]), .B(n_60422), .C(n_2829), .D(n_32290)
		, .Z(n_275360602));
	notech_reg_set sav_epc_reg_31(.CP(n_63520), .D(n_22030), .SD(1'b1), .Q(sav_epc
		[31]));
	notech_mux2 i_3732(.S(n_55771), .A(sav_epc[31]), .B(regs_14[31]), .Z(n_22030
		));
	notech_reg_set all_cnt_reg_0(.CP(n_63520), .D(n_22036), .SD(1'b1), .Q(all_cnt
		[0]));
	notech_mux2 i_3740(.S(\nbus_11280[0] ), .A(all_cnt[0]), .B(n_30758), .Z(n_22036
		));
	notech_reg_set all_cnt_reg_1(.CP(n_63460), .D(n_22042), .SD(1'b1), .Q(all_cnt
		[1]));
	notech_mux2 i_3748(.S(\nbus_11280[0] ), .A(all_cnt[1]), .B(n_30897), .Z(n_22042
		));
	notech_ao4 i_179741563(.A(n_58592), .B(n_32021), .C(n_58561), .D(n_31989
		), .Z(n_275060599));
	notech_reg_set all_cnt_reg_2(.CP(n_63460), .D(n_22048), .SD(1'b1), .Q(all_cnt
		[2]));
	notech_mux2 i_3756(.S(\nbus_11280[0] ), .A(all_cnt[2]), .B(n_177094253),
		 .Z(n_22048));
	notech_ao4 i_179841562(.A(n_58570), .B(n_31433), .C(n_57524), .D(n_33116
		), .Z(n_274960598));
	notech_reg_set all_cnt_reg_3(.CP(n_63460), .D(n_22054), .SD(1'b1), .Q(all_cnt
		[3]));
	notech_mux2 i_3764(.S(\nbus_11280[0] ), .A(all_cnt[3]), .B(n_177194254),
		 .Z(n_22054));
	notech_and2 i_180441558(.A(n_274760596), .B(n_274660595), .Z(n_274860597
		));
	notech_reg regs_reg_14_0(.CP(n_63460), .D(n_22060), .CD(n_62425), .Q(regs_14
		[0]));
	notech_mux2 i_3772(.S(n_30448), .A(n_19894), .B(regs_14[0]), .Z(n_22060)
		);
	notech_ao4 i_180141560(.A(n_57444), .B(n_31597), .C(n_57429), .D(n_31957
		), .Z(n_274760596));
	notech_reg regs_reg_14_1(.CP(n_63460), .D(n_22066), .CD(n_62424), .Q(regs_14
		[1]));
	notech_mux2 i_3780(.S(n_30448), .A(n_19900), .B(regs_14[1]), .Z(n_22066)
		);
	notech_ao4 i_180341559(.A(n_57412), .B(n_31924), .C(n_57401), .D(n_31892
		), .Z(n_274660595));
	notech_reg regs_reg_14_2(.CP(n_63460), .D(n_22072), .CD(n_62424), .Q(regs_14
		[2]));
	notech_mux2 i_3788(.S(n_30448), .A(n_4410), .B(regs_14[2]), .Z(n_22072)
		);
	notech_and4 i_181541550(.A(n_274360592), .B(n_274260591), .C(n_2740), .D
		(n_2739), .Z(n_274560594));
	notech_reg regs_reg_14_3(.CP(n_63460), .D(n_22078), .CD(n_62424), .Q(regs_14
		[3]));
	notech_mux2 i_3796(.S(n_30448), .A(n_4409), .B(regs_14[3]), .Z(n_22078)
		);
	notech_reg regs_reg_14_4(.CP(n_63460), .D(n_22084), .CD(n_62424), .Q(regs_14
		[4]));
	notech_mux2 i_3804(.S(n_30448), .A(n_4408), .B(regs_14[4]), .Z(n_22084)
		);
	notech_ao4 i_180641556(.A(n_57512), .B(n_31860), .C(n_58550), .D(n_31828
		), .Z(n_274360592));
	notech_reg regs_reg_14_5(.CP(n_63460), .D(n_22090), .CD(n_62425), .Q(regs_14
		[5]));
	notech_mux2 i_3812(.S(n_30448), .A(n_19924), .B(regs_14[5]), .Z(n_22090)
		);
	notech_ao4 i_180741555(.A(n_57500), .B(n_31796), .C(n_57489), .D(n_31764
		), .Z(n_274260591));
	notech_reg regs_reg_14_6(.CP(n_63460), .D(n_22096), .CD(n_62425), .Q(regs_14
		[6]));
	notech_mux2 i_3820(.S(n_30448), .A(n_19930), .B(regs_14[6]), .Z(n_22096)
		);
	notech_reg regs_reg_14_7(.CP(n_63600), .D(n_22102), .CD(n_62425), .Q(regs_14
		[7]));
	notech_mux2 i_3828(.S(n_30448), .A(n_19936), .B(regs_14[7]), .Z(n_22102)
		);
	notech_ao4 i_180941553(.A(n_57622), .B(n_33115), .C(n_57476), .D(n_31732
		), .Z(n_2740));
	notech_reg regs_reg_14_8(.CP(n_63458), .D(n_22108), .CD(n_62425), .Q(regs_14
		[8]));
	notech_mux2 i_3836(.S(n_30448), .A(n_19942), .B(regs_14[8]), .Z(n_22108)
		);
	notech_ao4 i_181041552(.A(n_57467), .B(n_31700), .C(n_57456), .D(n_31668
		), .Z(n_2739));
	notech_reg regs_reg_14_9(.CP(n_63458), .D(n_22114), .CD(n_62425), .Q(regs_14
		[9]));
	notech_mux2 i_3844(.S(n_30448), .A(n_4422), .B(regs_14[9]), .Z(n_22114)
		);
	notech_reg_set regs_reg_14_10(.CP(n_63508), .D(n_22120), .SD(n_62420), .Q
		(regs_14[10]));
	notech_mux2 i_3852(.S(n_30448), .A(n_389464425), .B(regs_14[10]), .Z(n_22120
		));
	notech_reg_set regs_reg_14_11(.CP(n_63508), .D(n_22126), .SD(n_62420), .Q
		(regs_14[11]));
	notech_mux2 i_3860(.S(n_30448), .A(n_446368047), .B(regs_14[11]), .Z(n_22126
		));
	notech_ao4 i_181641549(.A(n_58592), .B(n_32020), .C(n_58561), .D(n_31988
		), .Z(n_273660587));
	notech_reg_set regs_reg_14_12(.CP(n_63508), .D(n_22132), .SD(n_62420), .Q
		(regs_14[12]));
	notech_mux2 i_3868(.S(n_30448), .A(n_446268046), .B(regs_14[12]), .Z(n_22132
		));
	notech_ao4 i_181741548(.A(n_58570), .B(n_31432), .C(n_57524), .D(n_33114
		), .Z(n_273560586));
	notech_reg_set regs_reg_14_13(.CP(n_63508), .D(n_22138), .SD(n_62420), .Q
		(regs_14[13]));
	notech_mux2 i_3876(.S(n_30448), .A(n_389364424), .B(regs_14[13]), .Z(n_22138
		));
	notech_and2 i_182141544(.A(n_273360584), .B(n_273160583), .Z(n_273460585
		));
	notech_reg_set regs_reg_14_14(.CP(n_63508), .D(n_22144), .SD(n_62420), .Q
		(regs_14[14]));
	notech_mux2 i_3885(.S(n_30448), .A(n_19978), .B(regs_14[14]), .Z(n_22144
		));
	notech_ao4 i_181941546(.A(n_57444), .B(n_31596), .C(n_57429), .D(n_31956
		), .Z(n_273360584));
	notech_reg_set regs_reg_14_15(.CP(n_63508), .D(n_22150), .SD(n_62420), .Q
		(regs_14[15]));
	notech_mux2 i_3893(.S(n_30448), .A(n_446168045), .B(regs_14[15]), .Z(n_22150
		));
	notech_ao4 i_182041545(.A(n_57412), .B(n_31923), .C(n_57401), .D(n_31891
		), .Z(n_273160583));
	notech_reg_set regs_reg_14_16(.CP(n_63508), .D(n_22156), .SD(n_62420), .Q
		(regs_14[16]));
	notech_mux2 i_3901(.S(n_57045), .A(n_19990), .B(regs_14[16]), .Z(n_22156
		));
	notech_and4 i_182941536(.A(n_272860580), .B(n_272760579), .C(n_272560577
		), .D(n_272460576), .Z(n_273060582));
	notech_reg_set regs_reg_14_17(.CP(n_63508), .D(n_22162), .SD(n_62420), .Q
		(regs_14[17]));
	notech_mux2 i_3909(.S(n_57045), .A(n_19996), .B(regs_14[17]), .Z(n_22162
		));
	notech_reg_set regs_reg_14_18(.CP(n_63508), .D(n_22168), .SD(n_62420), .Q
		(regs_14[18]));
	notech_mux2 i_3917(.S(n_57045), .A(n_20002), .B(regs_14[18]), .Z(n_22168
		));
	notech_ao4 i_182341542(.A(n_57512), .B(n_31859), .C(n_58550), .D(n_31827
		), .Z(n_272860580));
	notech_reg_set regs_reg_14_19(.CP(n_63508), .D(n_22174), .SD(n_62420), .Q
		(regs_14[19]));
	notech_mux2 i_3925(.S(n_57045), .A(n_20008), .B(regs_14[19]), .Z(n_22174
		));
	notech_ao4 i_182441541(.A(n_57500), .B(n_31795), .C(n_57489), .D(n_31763
		), .Z(n_272760579));
	notech_reg regs_reg_14_20(.CP(n_63592), .D(n_22180), .CD(n_62419), .Q(regs_14
		[20]));
	notech_mux2 i_3933(.S(n_57045), .A(n_20014), .B(regs_14[20]), .Z(n_22180
		));
	notech_reg regs_reg_14_21(.CP(n_63592), .D(n_22186), .CD(n_62419), .Q(regs_14
		[21]));
	notech_mux2 i_3941(.S(n_57045), .A(n_20020), .B(regs_14[21]), .Z(n_22186
		));
	notech_ao4 i_182641539(.A(n_57622), .B(n_33113), .C(n_57480), .D(n_31731
		), .Z(n_272560577));
	notech_reg regs_reg_14_22(.CP(n_63592), .D(n_22192), .CD(n_62419), .Q(regs_14
		[22]));
	notech_mux2 i_3952(.S(n_57045), .A(n_20026), .B(regs_14[22]), .Z(n_22192
		));
	notech_ao4 i_182741538(.A(n_57467), .B(n_31699), .C(n_57456), .D(n_31667
		), .Z(n_272460576));
	notech_reg regs_reg_14_23(.CP(n_63592), .D(n_22198), .CD(n_62419), .Q(regs_14
		[23]));
	notech_mux2 i_3963(.S(n_57045), .A(n_20032), .B(regs_14[23]), .Z(n_22198
		));
	notech_reg regs_reg_14_24(.CP(n_63592), .D(n_22204), .CD(n_62419), .Q(regs_14
		[24]));
	notech_mux2 i_3971(.S(n_57045), .A(n_20038), .B(regs_14[24]), .Z(n_22204
		));
	notech_reg regs_reg_14_25(.CP(n_63592), .D(n_22210), .CD(n_62419), .Q(regs_14
		[25]));
	notech_mux2 i_3979(.S(n_57045), .A(n_20044), .B(regs_14[25]), .Z(n_22210
		));
	notech_ao4 i_183041535(.A(n_58596), .B(n_32019), .C(n_58565), .D(n_31987
		), .Z(n_272160573));
	notech_reg regs_reg_14_26(.CP(n_63592), .D(n_22216), .CD(n_62419), .Q(regs_14
		[26]));
	notech_mux2 i_3987(.S(n_57045), .A(n_20050), .B(regs_14[26]), .Z(n_22216
		));
	notech_ao4 i_183141534(.A(n_58570), .B(n_31431), .C(n_57524), .D(n_33112
		), .Z(n_272060572));
	notech_reg regs_reg_14_27(.CP(n_63592), .D(n_22222), .CD(n_62419), .Q(regs_14
		[27]));
	notech_mux2 i_3995(.S(n_57045), .A(n_20056), .B(regs_14[27]), .Z(n_22222
		));
	notech_and2 i_183641530(.A(n_271860570), .B(n_271760569), .Z(n_271960571
		));
	notech_reg regs_reg_14_28(.CP(n_63592), .D(n_22228), .CD(n_62419), .Q(regs_14
		[28]));
	notech_mux2 i_4003(.S(n_57045), .A(n_20062), .B(regs_14[28]), .Z(n_22228
		));
	notech_ao4 i_183341532(.A(n_57444), .B(n_31595), .C(n_57429), .D(n_31955
		), .Z(n_271860570));
	notech_reg regs_reg_14_29(.CP(n_63592), .D(n_22234), .CD(n_62421), .Q(regs_14
		[29]));
	notech_mux2 i_4011(.S(n_57045), .A(n_20068), .B(regs_14[29]), .Z(n_22234
		));
	notech_ao4 i_183441531(.A(n_57412), .B(n_31922), .C(n_57406), .D(n_31890
		), .Z(n_271760569));
	notech_reg regs_reg_14_30(.CP(n_63592), .D(n_22240), .CD(n_62421), .Q(regs_14
		[30]));
	notech_mux2 i_4019(.S(n_57045), .A(n_20074), .B(regs_14[30]), .Z(n_22240
		));
	notech_and4 i_184541522(.A(n_271460566), .B(n_271360565), .C(n_271160563
		), .D(n_270960562), .Z(n_271660568));
	notech_reg regs_reg_14_31(.CP(n_63592), .D(n_22246), .CD(n_62421), .Q(regs_14
		[31]));
	notech_mux2 i_4027(.S(n_57045), .A(n_20080), .B(regs_14[31]), .Z(n_22246
		));
	notech_reg regs_reg_13_0(.CP(n_63592), .D(n_22252), .CD(n_62421), .Q(gs[
		0]));
	notech_mux2 i_4035(.S(n_173966175), .A(n_195666383), .B(gs[0]), .Z(n_22252
		));
	notech_ao4 i_183941528(.A(n_57512), .B(n_31858), .C(n_58550), .D(n_31826
		), .Z(n_271460566));
	notech_reg regs_reg_13_1(.CP(n_63592), .D(n_22258), .CD(n_62421), .Q(gs[
		1]));
	notech_mux2 i_4043(.S(n_173966175), .A(n_30440), .B(gs[1]), .Z(n_22258)
		);
	notech_ao4 i_184041527(.A(n_57500), .B(n_31794), .C(n_57489), .D(n_31762
		), .Z(n_271360565));
	notech_reg regs_reg_13_2(.CP(n_63592), .D(n_22264), .CD(n_62423), .Q(gs[
		2]));
	notech_mux2 i_4051(.S(n_173966175), .A(n_194466371), .B(n_56951), .Z(n_22264
		));
	notech_reg regs_reg_13_3(.CP(n_63592), .D(n_22270), .CD(n_62423), .Q(gs[
		3]));
	notech_mux2 i_4059(.S(n_173966175), .A(n_19586), .B(gs[3]), .Z(n_22270)
		);
	notech_ao4 i_184241525(.A(n_57622), .B(n_33111), .C(n_57480), .D(n_31730
		), .Z(n_271160563));
	notech_reg regs_reg_13_4(.CP(n_63592), .D(n_22276), .CD(n_62421), .Q(gs[
		4]));
	notech_mux2 i_4067(.S(n_173966175), .A(n_19592), .B(gs[4]), .Z(n_22276)
		);
	notech_ao4 i_184341524(.A(n_57471), .B(n_31698), .C(n_57456), .D(n_31666
		), .Z(n_270960562));
	notech_reg regs_reg_13_5(.CP(n_63592), .D(n_22282), .CD(n_62423), .Q(gs[
		5]));
	notech_mux2 i_4075(.S(n_173966175), .A(n_4365), .B(gs[5]), .Z(n_22282)
		);
	notech_reg regs_reg_13_6(.CP(n_63592), .D(n_22288), .CD(n_62421), .Q(gs[
		6]));
	notech_mux2 i_4083(.S(n_173966175), .A(n_193166358), .B(gs[6]), .Z(n_22288
		));
	notech_reg regs_reg_13_7(.CP(n_63590), .D(n_22294), .CD(n_62420), .Q(gs[
		7]));
	notech_mux2 i_4091(.S(n_173966175), .A(n_1505), .B(gs[7]), .Z(n_22294)
		);
	notech_ao4 i_201041367(.A(n_58596), .B(n_32005), .C(n_58565), .D(n_31973
		), .Z(n_270660559));
	notech_reg regs_reg_13_8(.CP(n_63590), .D(n_22300), .CD(n_62421), .Q(gs[
		8]));
	notech_mux2 i_4099(.S(n_173966175), .A(n_446468048), .B(gs[8]), .Z(n_22300
		));
	notech_ao4 i_201141366(.A(n_58574), .B(n_31417), .C(n_57524), .D(n_33131
		), .Z(n_270560558));
	notech_reg regs_reg_13_9(.CP(n_63662), .D(n_22306), .CD(n_62420), .Q(gs[
		9]));
	notech_mux2 i_4107(.S(n_173966175), .A(n_191866345), .B(gs[9]), .Z(n_22306
		));
	notech_and2 i_201541362(.A(n_270360556), .B(n_270260555), .Z(n_270460557
		));
	notech_reg regs_reg_13_10(.CP(n_63662), .D(n_22312), .CD(n_62420), .Q(gs
		[10]));
	notech_mux2 i_4115(.S(n_173966175), .A(n_167462706), .B(gs[10]), .Z(n_22312
		));
	notech_ao4 i_201341364(.A(n_57444), .B(n_31581), .C(n_57429), .D(n_31940
		), .Z(n_270360556));
	notech_reg regs_reg_13_11(.CP(n_63662), .D(n_22318), .CD(n_62421), .Q(gs
		[11]));
	notech_mux2 i_4123(.S(n_173966175), .A(n_190766334), .B(gs[11]), .Z(n_22318
		));
	notech_ao4 i_201441363(.A(n_57412), .B(n_31908), .C(n_57406), .D(n_31876
		), .Z(n_270260555));
	notech_reg regs_reg_13_12(.CP(n_63662), .D(n_22324), .CD(n_62421), .Q(gs
		[12]));
	notech_mux2 i_4131(.S(n_173966175), .A(n_189666323), .B(gs[12]), .Z(n_22324
		));
	notech_and4 i_202441354(.A(n_269960552), .B(n_269860551), .C(n_269660549
		), .D(n_269560548), .Z(n_270160554));
	notech_reg regs_reg_13_13(.CP(n_63662), .D(n_22331), .CD(n_62421), .Q(gs
		[13]));
	notech_mux2 i_4139(.S(n_173966175), .A(n_166362695), .B(gs[13]), .Z(n_22331
		));
	notech_reg regs_reg_13_14(.CP(n_63662), .D(n_22337), .CD(n_62421), .Q(gs
		[14]));
	notech_mux2 i_4147(.S(n_173966175), .A(n_30447), .B(gs[14]), .Z(n_22337)
		);
	notech_ao4 i_201741360(.A(n_57512), .B(n_31844), .C(n_58550), .D(n_31812
		), .Z(n_269960552));
	notech_reg regs_reg_13_15(.CP(n_63662), .D(n_22343), .CD(n_62421), .Q(gs
		[15]));
	notech_mux2 i_4155(.S(n_173966175), .A(n_187466301), .B(gs[15]), .Z(n_22343
		));
	notech_ao4 i_201841359(.A(n_57500), .B(n_31780), .C(n_57489), .D(n_31748
		), .Z(n_269860551));
	notech_reg regs_reg_13_16(.CP(n_63662), .D(n_22349), .CD(n_62432), .Q(gs
		[16]));
	notech_mux2 i_4163(.S(n_55820), .A(n_19664), .B(gs[16]), .Z(n_22349));
	notech_reg regs_reg_13_17(.CP(n_63662), .D(n_22355), .CD(n_62432), .Q(gs
		[17]));
	notech_mux2 i_4171(.S(n_55820), .A(n_19670), .B(gs[17]), .Z(n_22355));
	notech_ao4 i_202041357(.A(n_57622), .B(n_33132), .C(n_57480), .D(n_31716
		), .Z(n_269660549));
	notech_reg regs_reg_13_18(.CP(n_63662), .D(n_22361), .CD(n_62431), .Q(gs
		[18]));
	notech_mux2 i_4179(.S(n_55820), .A(n_19676), .B(gs[18]), .Z(n_22361));
	notech_ao4 i_202141356(.A(n_57471), .B(n_31684), .C(n_57456), .D(n_31652
		), .Z(n_269560548));
	notech_reg regs_reg_13_19(.CP(n_63662), .D(n_22367), .CD(n_62431), .Q(gs
		[19]));
	notech_mux2 i_4187(.S(n_55820), .A(n_19682), .B(gs[19]), .Z(n_22367));
	notech_reg regs_reg_13_20(.CP(n_63662), .D(n_22373), .CD(n_62432), .Q(gs
		[20]));
	notech_mux2 i_4195(.S(n_55820), .A(n_19688), .B(gs[20]), .Z(n_22373));
	notech_reg regs_reg_13_21(.CP(n_63662), .D(n_22379), .CD(n_62432), .Q(gs
		[21]));
	notech_mux2 i_4203(.S(n_55820), .A(n_19694), .B(gs[21]), .Z(n_22379));
	notech_ao4 i_204041339(.A(n_58596), .B(n_32003), .C(n_58565), .D(n_31971
		), .Z(n_269260545));
	notech_reg regs_reg_13_22(.CP(n_63662), .D(n_22385), .CD(n_62432), .Q(gs
		[22]));
	notech_mux2 i_4211(.S(n_55820), .A(n_19700), .B(gs[22]), .Z(n_22385));
	notech_ao4 i_204241338(.A(n_58574), .B(n_31415), .C(n_57524), .D(n_33121
		), .Z(n_269160544));
	notech_reg regs_reg_13_23(.CP(n_63662), .D(n_22391), .CD(n_62432), .Q(gs
		[23]));
	notech_mux2 i_4219(.S(n_55820), .A(n_19706), .B(gs[23]), .Z(n_22391));
	notech_and2 i_204641334(.A(n_268960542), .B(n_268660541), .Z(n_269060543
		));
	notech_reg regs_reg_13_24(.CP(n_63662), .D(n_22397), .CD(n_62432), .Q(gs
		[24]));
	notech_mux2 i_4227(.S(n_55820), .A(n_3442), .B(gs[24]), .Z(n_22397));
	notech_ao4 i_204441336(.A(n_57444), .B(n_31579), .C(n_57429), .D(n_31938
		), .Z(n_268960542));
	notech_reg regs_reg_13_25(.CP(n_63662), .D(n_22403), .CD(n_62431), .Q(gs
		[25]));
	notech_mux2 i_4235(.S(n_55820), .A(n_19718), .B(gs[25]), .Z(n_22403));
	notech_ao4 i_204541335(.A(n_57412), .B(n_31906), .C(n_57406), .D(n_31874
		), .Z(n_268660541));
	notech_reg regs_reg_13_26(.CP(n_63662), .D(n_22409), .CD(n_62431), .Q(gs
		[26]));
	notech_mux2 i_4243(.S(n_55820), .A(n_19724), .B(gs[26]), .Z(n_22409));
	notech_and4 i_205441326(.A(n_268360538), .B(n_268260537), .C(n_268060535
		), .D(n_267960534), .Z(n_268560540));
	notech_reg regs_reg_13_27(.CP(n_63590), .D(n_22415), .CD(n_62431), .Q(gs
		[27]));
	notech_mux2 i_4251(.S(n_55820), .A(n_19730), .B(gs[27]), .Z(n_22415));
	notech_reg regs_reg_13_28(.CP(n_63590), .D(n_22421), .CD(n_62431), .Q(gs
		[28]));
	notech_mux2 i_4259(.S(n_55820), .A(n_19736), .B(gs[28]), .Z(n_22421));
	notech_ao4 i_204841332(.A(n_57512), .B(n_31842), .C(n_58550), .D(n_31810
		), .Z(n_268360538));
	notech_reg regs_reg_13_29(.CP(n_63590), .D(n_22427), .CD(n_62431), .Q(gs
		[29]));
	notech_mux2 i_4267(.S(n_55820), .A(n_30402), .B(gs[29]), .Z(n_22427));
	notech_ao4 i_204941331(.A(n_57500), .B(n_31778), .C(n_57489), .D(n_31746
		), .Z(n_268260537));
	notech_reg regs_reg_13_30(.CP(n_63590), .D(n_22433), .CD(n_62431), .Q(gs
		[30]));
	notech_mux2 i_4275(.S(n_55820), .A(n_19748), .B(gs[30]), .Z(n_22433));
	notech_reg regs_reg_13_31(.CP(n_63590), .D(n_22439), .CD(n_62431), .Q(gs
		[31]));
	notech_mux2 i_4283(.S(n_55820), .A(n_19754), .B(gs[31]), .Z(n_22439));
	notech_ao4 i_205141329(.A(n_57622), .B(n_33122), .C(n_57480), .D(n_31714
		), .Z(n_268060535));
	notech_reg regs_reg_12_0(.CP(n_63590), .D(n_22445), .CD(n_62431), .Q(regs_12
		[0]));
	notech_mux2 i_4291(.S(n_212880631), .A(n_201966439), .B(regs_12[0]), .Z(n_22445
		));
	notech_ao4 i_205241328(.A(n_57471), .B(n_31682), .C(n_57456), .D(n_31650
		), .Z(n_267960534));
	notech_reg regs_reg_12_1(.CP(n_63590), .D(n_22451), .CD(n_62431), .Q(regs_12
		[1]));
	notech_mux2 i_4299(.S(n_212880631), .A(n_439967983), .B(regs_12[1]), .Z(n_22451
		));
	notech_reg regs_reg_12_2(.CP(n_63590), .D(n_22458), .CD(n_62431), .Q(regs_12
		[2]));
	notech_mux2 i_4307(.S(n_212880631), .A(n_1545), .B(regs_12[2]), .Z(n_22458
		));
	notech_reg regs_reg_12_3(.CP(n_63590), .D(n_22464), .CD(n_62434), .Q(regs_12
		[3]));
	notech_mux2 i_4315(.S(n_212880631), .A(n_19238), .B(regs_12[3]), .Z(n_22464
		));
	notech_ao4 i_205541325(.A(n_58596), .B(n_32002), .C(n_58565), .D(n_31970
		), .Z(n_267660531));
	notech_reg regs_reg_12_4(.CP(n_63590), .D(n_22473), .CD(n_62434), .Q(regs_12
		[4]));
	notech_mux2 i_4323(.S(n_212880631), .A(n_19244), .B(regs_12[4]), .Z(n_22473
		));
	notech_ao4 i_205641324(.A(n_58574), .B(n_31414), .C(n_57529), .D(n_33123
		), .Z(n_267560530));
	notech_reg regs_reg_12_5(.CP(n_63662), .D(n_22482), .CD(n_62434), .Q(regs_12
		[5]));
	notech_mux2 i_4331(.S(n_212880631), .A(n_4366), .B(regs_12[5]), .Z(n_22482
		));
	notech_and2 i_206041320(.A(n_267360528), .B(n_267260527), .Z(n_267460529
		));
	notech_reg regs_reg_12_6(.CP(n_63658), .D(n_22488), .CD(n_62434), .Q(regs_12
		[6]));
	notech_mux2 i_4339(.S(n_212880631), .A(n_1531), .B(regs_12[6]), .Z(n_22488
		));
	notech_ao4 i_205841322(.A(n_57449), .B(n_31578), .C(n_57429), .D(n_31937
		), .Z(n_267360528));
	notech_reg regs_reg_12_7(.CP(n_63588), .D(n_22494), .CD(n_62434), .Q(regs_12
		[7]));
	notech_mux2 i_4347(.S(n_212880631), .A(n_1518), .B(regs_12[7]), .Z(n_22494
		));
	notech_ao4 i_205941321(.A(n_57412), .B(n_31905), .C(n_57406), .D(n_31873
		), .Z(n_267260527));
	notech_reg regs_reg_12_8(.CP(n_63658), .D(n_22500), .CD(n_62434), .Q(regs_12
		[8]));
	notech_mux2 i_4355(.S(n_212880631), .A(n_446568049), .B(regs_12[8]), .Z(n_22500
		));
	notech_and4 i_206841312(.A(n_266960524), .B(n_266860523), .C(n_266660521
		), .D(n_266560520), .Z(n_267160526));
	notech_reg regs_reg_12_9(.CP(n_63658), .D(n_22506), .CD(n_62434), .Q(regs_12
		[9]));
	notech_mux2 i_4363(.S(n_212880631), .A(n_200266427), .B(regs_12[9]), .Z(n_22506
		));
	notech_reg regs_reg_12_10(.CP(n_63658), .D(n_22512), .CD(n_62434), .Q(regs_12
		[10]));
	notech_mux2 i_4371(.S(n_212880631), .A(n_383764368), .B(regs_12[10]), .Z
		(n_22512));
	notech_ao4 i_206241318(.A(n_57512), .B(n_31841), .C(n_58550), .D(n_31809
		), .Z(n_266960524));
	notech_reg regs_reg_12_11(.CP(n_63658), .D(n_22518), .CD(n_62434), .Q(regs_12
		[11]));
	notech_mux2 i_4379(.S(n_212880631), .A(n_198966416), .B(regs_12[11]), .Z
		(n_22518));
	notech_ao4 i_206341317(.A(n_57500), .B(n_31777), .C(n_57489), .D(n_31745
		), .Z(n_266860523));
	notech_reg regs_reg_12_12(.CP(n_63658), .D(n_22524), .CD(n_62434), .Q(regs_12
		[12]));
	notech_mux2 i_4387(.S(n_212880631), .A(n_197866405), .B(regs_12[12]), .Z
		(n_22524));
	notech_reg regs_reg_12_13(.CP(n_63658), .D(n_22530), .CD(n_62432), .Q(regs_12
		[13]));
	notech_mux2 i_4395(.S(n_212880631), .A(n_168562717), .B(regs_12[13]), .Z
		(n_22530));
	notech_ao4 i_206541315(.A(n_57622), .B(n_33124), .C(n_57480), .D(n_31713
		), .Z(n_266660521));
	notech_reg regs_reg_12_14(.CP(n_63658), .D(n_22536), .CD(n_62432), .Q(regs_12
		[14]));
	notech_mux2 i_4403(.S(n_212880631), .A(n_30384), .B(regs_12[14]), .Z(n_22536
		));
	notech_ao4 i_206641314(.A(n_57471), .B(n_31681), .C(n_57461), .D(n_31649
		), .Z(n_266560520));
	notech_reg regs_reg_12_15(.CP(n_63658), .D(n_22542), .CD(n_62432), .Q(regs_12
		[15]));
	notech_mux2 i_4411(.S(n_212880631), .A(n_196766394), .B(regs_12[15]), .Z
		(n_22542));
	notech_reg regs_reg_12_16(.CP(n_63658), .D(n_22548), .CD(n_62432), .Q(regs_12
		[16]));
	notech_mux2 i_4419(.S(n_55840), .A(n_19316), .B(regs_12[16]), .Z(n_22548
		));
	notech_reg regs_reg_12_17(.CP(n_63658), .D(n_22554), .CD(n_62432), .Q(regs_12
		[17]));
	notech_mux2 i_4427(.S(n_55840), .A(n_19322), .B(regs_12[17]), .Z(n_22554
		));
	notech_ao4 i_206941311(.A(n_58596), .B(n_32001), .C(n_58565), .D(n_31969
		), .Z(n_266260517));
	notech_reg regs_reg_12_18(.CP(n_63658), .D(n_22560), .CD(n_62434), .Q(regs_12
		[18]));
	notech_mux2 i_4435(.S(n_55840), .A(n_19328), .B(regs_12[18]), .Z(n_22560
		));
	notech_ao4 i_207041310(.A(n_58574), .B(n_31413), .C(n_57524), .D(n_33125
		), .Z(n_266160516));
	notech_reg regs_reg_12_19(.CP(n_63690), .D(n_22566), .CD(n_62434), .Q(regs_12
		[19]));
	notech_mux2 i_4443(.S(n_55840), .A(n_19334), .B(regs_12[19]), .Z(n_22566
		));
	notech_and2 i_207441306(.A(n_265960514), .B(n_265860513), .Z(n_266060515
		));
	notech_reg regs_reg_12_20(.CP(n_63690), .D(n_22572), .CD(n_62432), .Q(regs_12
		[20]));
	notech_mux2 i_4451(.S(n_55840), .A(n_19340), .B(regs_12[20]), .Z(n_22572
		));
	notech_ao4 i_207241308(.A(n_57444), .B(n_31577), .C(n_57429), .D(n_31936
		), .Z(n_265960514));
	notech_reg regs_reg_12_21(.CP(n_63690), .D(n_22578), .CD(n_62434), .Q(regs_12
		[21]));
	notech_mux2 i_4459(.S(n_55840), .A(n_19346), .B(regs_12[21]), .Z(n_22578
		));
	notech_ao4 i_207341307(.A(n_57417), .B(n_31904), .C(n_57406), .D(n_31872
		), .Z(n_265860513));
	notech_reg regs_reg_12_22(.CP(n_63690), .D(n_22584), .CD(n_62429), .Q(regs_12
		[22]));
	notech_mux2 i_4467(.S(n_55840), .A(n_19352), .B(regs_12[22]), .Z(n_22584
		));
	notech_and4 i_208241298(.A(n_265560510), .B(n_265460509), .C(n_265260507
		), .D(n_265160506), .Z(n_265760512));
	notech_reg regs_reg_12_23(.CP(n_63690), .D(n_22590), .CD(n_62429), .Q(regs_12
		[23]));
	notech_mux2 i_4475(.S(n_55840), .A(n_19358), .B(regs_12[23]), .Z(n_22590
		));
	notech_reg regs_reg_12_24(.CP(n_63690), .D(n_22596), .CD(n_62426), .Q(regs_12
		[24]));
	notech_mux2 i_4483(.S(n_55840), .A(n_30913), .B(regs_12[24]), .Z(n_22596
		));
	notech_ao4 i_207641304(.A(n_57512), .B(n_31840), .C(n_58550), .D(n_31808
		), .Z(n_265560510));
	notech_reg regs_reg_12_25(.CP(n_63690), .D(n_22602), .CD(n_62429), .Q(regs_12
		[25]));
	notech_mux2 i_4491(.S(n_55840), .A(n_347367644), .B(regs_12[25]), .Z(n_22602
		));
	notech_ao4 i_207741303(.A(n_57500), .B(n_31776), .C(n_57489), .D(n_31744
		), .Z(n_265460509));
	notech_reg regs_reg_12_26(.CP(n_63690), .D(n_22608), .CD(n_62429), .Q(regs_12
		[26]));
	notech_mux2 i_4499(.S(n_55840), .A(n_19376), .B(regs_12[26]), .Z(n_22608
		));
	notech_reg regs_reg_12_27(.CP(n_63690), .D(n_22614), .CD(n_62429), .Q(regs_12
		[27]));
	notech_mux2 i_4507(.S(n_55840), .A(n_19382), .B(regs_12[27]), .Z(n_22614
		));
	notech_ao4 i_207941301(.A(n_57622), .B(n_33126), .C(n_57480), .D(n_31712
		), .Z(n_265260507));
	notech_reg regs_reg_12_28(.CP(n_63690), .D(n_22620), .CD(n_62429), .Q(regs_12
		[28]));
	notech_mux2 i_4515(.S(n_55840), .A(n_19388), .B(regs_12[28]), .Z(n_22620
		));
	notech_ao4 i_208041300(.A(n_57471), .B(n_31680), .C(n_57456), .D(n_31648
		), .Z(n_265160506));
	notech_reg regs_reg_12_29(.CP(n_63690), .D(n_22626), .CD(n_62429), .Q(regs_12
		[29]));
	notech_mux2 i_4523(.S(n_55840), .A(n_30403), .B(regs_12[29]), .Z(n_22626
		));
	notech_reg regs_reg_12_30(.CP(n_63690), .D(n_22632), .CD(n_62429), .Q(regs_12
		[30]));
	notech_mux2 i_4531(.S(n_55840), .A(n_19400), .B(regs_12[30]), .Z(n_22632
		));
	notech_reg regs_reg_12_31(.CP(n_63690), .D(n_22638), .CD(n_62426), .Q(regs_12
		[31]));
	notech_mux2 i_4539(.S(n_55840), .A(n_19406), .B(regs_12[31]), .Z(n_22638
		));
	notech_ao4 i_208341297(.A(n_58592), .B(n_32000), .C(n_58561), .D(n_31968
		), .Z(n_264860503));
	notech_reg regs_reg_11_0(.CP(n_63690), .D(n_22644), .CD(n_62426), .Q(regs_11
		[0]));
	notech_mux2 i_4547(.S(n_176766199), .A(n_30388), .B(regs_11[0]), .Z(n_22644
		));
	notech_ao4 i_208441296(.A(n_58574), .B(n_31412), .C(n_57524), .D(n_33127
		), .Z(n_264760502));
	notech_reg regs_reg_11_1(.CP(n_63690), .D(n_22650), .CD(n_62426), .Q(regs_11
		[1]));
	notech_mux2 i_4555(.S(n_176766199), .A(n_4368), .B(regs_11[1]), .Z(n_22650
		));
	notech_and2 i_208841292(.A(n_264560500), .B(n_264460499), .Z(n_264660501
		));
	notech_reg regs_reg_11_2(.CP(n_63690), .D(n_22656), .CD(n_62426), .Q(regs_11
		[2]));
	notech_mux2 i_4563(.S(n_176766199), .A(n_172062752), .B(regs_11[2]), .Z(n_22656
		));
	notech_ao4 i_208641294(.A(n_57444), .B(n_31576), .C(n_57429), .D(n_31935
		), .Z(n_264560500));
	notech_reg regs_reg_11_3(.CP(n_63690), .D(n_22662), .CD(n_62426), .Q(regs_11
		[3]));
	notech_mux2 i_4571(.S(n_176766199), .A(n_18890), .B(regs_11[3]), .Z(n_22662
		));
	notech_ao4 i_208741293(.A(n_57412), .B(n_31903), .C(n_57406), .D(n_31871
		), .Z(n_264460499));
	notech_reg regs_reg_11_4(.CP(n_63690), .D(n_22668), .CD(n_62426), .Q(regs_11
		[4]));
	notech_mux2 i_4579(.S(n_176766199), .A(n_18896), .B(regs_11[4]), .Z(n_22668
		));
	notech_and4 i_209641284(.A(n_264160496), .B(n_264060495), .C(n_2638), .D
		(n_2637), .Z(n_264360498));
	notech_reg regs_reg_11_5(.CP(n_63658), .D(n_22674), .CD(n_62426), .Q(regs_11
		[5]));
	notech_mux2 i_4587(.S(n_176766199), .A(n_4367), .B(regs_11[5]), .Z(n_22674
		));
	notech_reg regs_reg_11_6(.CP(n_63690), .D(n_22680), .CD(n_62426), .Q(regs_11
		[6]));
	notech_mux2 i_4595(.S(n_176766199), .A(n_18908), .B(regs_11[6]), .Z(n_22680
		));
	notech_ao4 i_209041290(.A(n_57512), .B(n_31839), .C(n_58550), .D(n_31807
		), .Z(n_264160496));
	notech_reg regs_reg_11_7(.CP(n_63660), .D(n_22686), .CD(n_62426), .Q(regs_11
		[7]));
	notech_mux2 i_4603(.S(n_176766199), .A(n_18914), .B(regs_11[7]), .Z(n_22686
		));
	notech_ao4 i_209141289(.A(n_57500), .B(n_31775), .C(n_57489), .D(n_31743
		), .Z(n_264060495));
	notech_reg regs_reg_11_8(.CP(n_63660), .D(n_22692), .CD(n_62426), .Q(regs_11
		[8]));
	notech_mux2 i_4611(.S(n_176766199), .A(n_18920), .B(regs_11[8]), .Z(n_22692
		));
	notech_reg regs_reg_11_9(.CP(n_63660), .D(n_22698), .CD(n_62430), .Q(regs_11
		[9]));
	notech_mux2 i_4619(.S(n_176766199), .A(n_216480665), .B(regs_11[9]), .Z(n_22698
		));
	notech_ao4 i_209341287(.A(n_57622), .B(n_33128), .C(n_57480), .D(n_31711
		), .Z(n_2638));
	notech_reg regs_reg_11_10(.CP(n_63660), .D(n_22704), .CD(n_62430), .Q(regs_11
		[10]));
	notech_mux2 i_4627(.S(n_176766199), .A(n_170762739), .B(regs_11[10]), .Z
		(n_22704));
	notech_ao4 i_209441286(.A(n_57467), .B(n_31679), .C(n_57456), .D(n_31647
		), .Z(n_2637));
	notech_reg regs_reg_11_11(.CP(n_63660), .D(n_22710), .CD(n_62430), .Q(regs_11
		[11]));
	notech_mux2 i_4635(.S(n_176766199), .A(n_205466472), .B(regs_11[11]), .Z
		(n_22710));
	notech_reg regs_reg_11_12(.CP(n_63660), .D(n_22716), .CD(n_62430), .Q(regs_11
		[12]));
	notech_mux2 i_4643(.S(n_176766199), .A(n_204266461), .B(regs_11[12]), .Z
		(n_22716));
	notech_reg regs_reg_11_13(.CP(n_63660), .D(n_22722), .CD(n_62430), .Q(regs_11
		[13]));
	notech_mux2 i_4651(.S(n_176766199), .A(n_169662728), .B(regs_11[13]), .Z
		(n_22722));
	notech_ao4 i_209741283(.A(n_58592), .B(n_31999), .C(n_58561), .D(n_31967
		), .Z(n_2634));
	notech_reg regs_reg_11_14(.CP(n_63660), .D(n_22728), .CD(n_62430), .Q(regs_11
		[14]));
	notech_mux2 i_4659(.S(n_176766199), .A(n_30385), .B(regs_11[14]), .Z(n_22728
		));
	notech_ao4 i_209841282(.A(n_58574), .B(n_31411), .C(n_57524), .D(n_33119
		), .Z(n_2633));
	notech_reg regs_reg_11_15(.CP(n_63660), .D(n_22734), .CD(n_62431), .Q(regs_11
		[15]));
	notech_mux2 i_4667(.S(n_176766199), .A(n_203066450), .B(regs_11[15]), .Z
		(n_22734));
	notech_and2 i_210241278(.A(n_2631), .B(n_2630), .Z(n_2632));
	notech_reg regs_reg_11_16(.CP(n_63660), .D(n_22740), .CD(n_62430), .Q(regs_11
		[16]));
	notech_mux2 i_4675(.S(n_55851), .A(n_18968), .B(regs_11[16]), .Z(n_22740
		));
	notech_ao4 i_210041280(.A(n_57444), .B(n_31575), .C(n_57429), .D(n_31934
		), .Z(n_2631));
	notech_reg regs_reg_11_17(.CP(n_63660), .D(n_22749), .CD(n_62430), .Q(regs_11
		[17]));
	notech_mux2 i_4683(.S(n_55851), .A(n_18974), .B(regs_11[17]), .Z(n_22749
		));
	notech_ao4 i_210141279(.A(n_57412), .B(n_31902), .C(n_57406), .D(n_31870
		), .Z(n_2630));
	notech_reg regs_reg_11_18(.CP(n_63660), .D(n_22756), .CD(n_62430), .Q(regs_11
		[18]));
	notech_mux2 i_4691(.S(n_55851), .A(n_18980), .B(regs_11[18]), .Z(n_22756
		));
	notech_and4 i_211041270(.A(n_2627), .B(n_2626), .C(n_2624), .D(n_2623), 
		.Z(n_2629));
	notech_reg regs_reg_11_19(.CP(n_63660), .D(n_22762), .CD(n_62429), .Q(regs_11
		[19]));
	notech_mux2 i_4699(.S(n_55851), .A(n_18986), .B(regs_11[19]), .Z(n_22762
		));
	notech_reg regs_reg_11_20(.CP(n_63660), .D(n_22768), .CD(n_62429), .Q(regs_11
		[20]));
	notech_mux2 i_4707(.S(n_55851), .A(n_18992), .B(regs_11[20]), .Z(n_22768
		));
	notech_ao4 i_210441276(.A(n_57512), .B(n_31838), .C(n_58550), .D(n_31806
		), .Z(n_2627));
	notech_reg regs_reg_11_21(.CP(n_63660), .D(n_22774), .CD(n_62429), .Q(regs_11
		[21]));
	notech_mux2 i_4715(.S(n_55851), .A(n_18998), .B(regs_11[21]), .Z(n_22774
		));
	notech_ao4 i_210541275(.A(n_57500), .B(n_31774), .C(n_57489), .D(n_31742
		), .Z(n_2626));
	notech_reg regs_reg_11_22(.CP(n_63660), .D(n_22780), .CD(n_62429), .Q(regs_11
		[22]));
	notech_mux2 i_4723(.S(n_55851), .A(n_348567653), .B(regs_11[22]), .Z(n_22780
		));
	notech_reg regs_reg_11_23(.CP(n_63660), .D(n_22787), .CD(n_62429), .Q(regs_11
		[23]));
	notech_mux2 i_4731(.S(n_55851), .A(n_19010), .B(regs_11[23]), .Z(n_22787
		));
	notech_ao4 i_210741273(.A(n_57622), .B(n_33120), .C(n_57480), .D(n_31710
		), .Z(n_2624));
	notech_reg regs_reg_11_24(.CP(n_63660), .D(n_22793), .CD(n_62430), .Q(regs_11
		[24]));
	notech_mux2 i_4739(.S(n_55851), .A(n_19016), .B(regs_11[24]), .Z(n_22793
		));
	notech_ao4 i_210841272(.A(n_57467), .B(n_31678), .C(n_57456), .D(n_31646
		), .Z(n_2623));
	notech_reg regs_reg_11_25(.CP(n_63660), .D(n_22799), .CD(n_62430), .Q(regs_11
		[25]));
	notech_mux2 i_4747(.S(n_55851), .A(n_19022), .B(regs_11[25]), .Z(n_22799
		));
	notech_reg regs_reg_11_26(.CP(n_63588), .D(n_22805), .CD(n_62430), .Q(regs_11
		[26]));
	notech_mux2 i_4755(.S(n_55851), .A(n_19028), .B(regs_11[26]), .Z(n_22805
		));
	notech_reg regs_reg_11_27(.CP(n_63588), .D(n_22811), .CD(n_62430), .Q(regs_11
		[27]));
	notech_mux2 i_4763(.S(n_55851), .A(n_19034), .B(regs_11[27]), .Z(n_22811
		));
	notech_ao4 i_211141269(.A(n_58592), .B(n_31997), .C(n_58561), .D(n_31965
		), .Z(n_2620));
	notech_reg regs_reg_11_28(.CP(n_63588), .D(n_22817), .CD(n_62474), .Q(regs_11
		[28]));
	notech_mux2 i_4771(.S(n_55851), .A(n_19040), .B(regs_11[28]), .Z(n_22817
		));
	notech_ao4 i_211241268(.A(n_58574), .B(n_31409), .C(n_57524), .D(n_33133
		), .Z(n_2619));
	notech_reg regs_reg_11_29(.CP(n_63588), .D(n_22823), .CD(n_62474), .Q(regs_11
		[29]));
	notech_mux2 i_4779(.S(n_55851), .A(n_30404), .B(regs_11[29]), .Z(n_22823
		));
	notech_and2 i_211641264(.A(n_2617), .B(n_2616), .Z(n_2618));
	notech_reg regs_reg_11_30(.CP(n_63588), .D(n_22829), .CD(n_62474), .Q(regs_11
		[30]));
	notech_mux2 i_4787(.S(n_55851), .A(n_19052), .B(regs_11[30]), .Z(n_22829
		));
	notech_ao4 i_211441266(.A(n_57444), .B(n_31573), .C(n_57429), .D(n_31932
		), .Z(n_2617));
	notech_reg regs_reg_11_31(.CP(n_63588), .D(n_22835), .CD(n_62474), .Q(regs_11
		[31]));
	notech_mux2 i_4795(.S(n_55851), .A(n_19058), .B(regs_11[31]), .Z(n_22835
		));
	notech_ao4 i_211541265(.A(n_57412), .B(n_31900), .C(n_57406), .D(n_31868
		), .Z(n_2616));
	notech_reg regs_reg_10_0(.CP(n_63588), .D(n_22841), .CD(n_62474), .Q(regs_10
		[0]));
	notech_mux2 i_4803(.S(n_442068004), .A(n_30924), .B(regs_10[0]), .Z(n_22841
		));
	notech_and4 i_212441256(.A(n_2613), .B(n_2612), .C(n_2610), .D(n_260960492
		), .Z(n_2615));
	notech_reg regs_reg_10_1(.CP(n_63588), .D(n_22847), .CD(n_62475), .Q(regs_10
		[1]));
	notech_mux2 i_4811(.S(n_442068004), .A(n_18530), .B(regs_10[1]), .Z(n_22847
		));
	notech_reg regs_reg_10_2(.CP(n_63588), .D(n_22853), .CD(n_62475), .Q(regs_10
		[2]));
	notech_mux2 i_4819(.S(n_442068004), .A(n_4356), .B(regs_10[2]), .Z(n_22853
		));
	notech_ao4 i_211841262(.A(n_57512), .B(n_31836), .C(n_58550), .D(n_31804
		), .Z(n_2613));
	notech_reg regs_reg_10_3(.CP(n_63588), .D(n_22859), .CD(n_62474), .Q(regs_10
		[3]));
	notech_mux2 i_4827(.S(n_442068004), .A(n_18542), .B(regs_10[3]), .Z(n_22859
		));
	notech_ao4 i_211941261(.A(n_57500), .B(n_31772), .C(n_57489), .D(n_31740
		), .Z(n_2612));
	notech_reg regs_reg_10_4(.CP(n_63508), .D(n_22865), .CD(n_62475), .Q(regs_10
		[4]));
	notech_mux2 i_4835(.S(n_442068004), .A(n_383964370), .B(regs_10[4]), .Z(n_22865
		));
	notech_reg regs_reg_10_5(.CP(n_63588), .D(n_22871), .CD(n_62474), .Q(regs_10
		[5]));
	notech_mux2 i_4843(.S(n_442068004), .A(n_4369), .B(regs_10[5]), .Z(n_22871
		));
	notech_ao4 i_212141259(.A(n_57622), .B(n_31368), .C(n_57480), .D(n_31708
		), .Z(n_2610));
	notech_reg regs_reg_10_6(.CP(n_63594), .D(n_22877), .CD(n_62471), .Q(regs_10
		[6]));
	notech_mux2 i_4851(.S(n_442068004), .A(n_18560), .B(regs_10[6]), .Z(n_22877
		));
	notech_ao4 i_212241258(.A(n_57467), .B(n_31676), .C(n_57456), .D(n_31644
		), .Z(n_260960492));
	notech_reg regs_reg_10_7(.CP(n_63510), .D(n_22883), .CD(n_62474), .Q(regs_10
		[7]));
	notech_mux2 i_4859(.S(n_442068004), .A(n_4355), .B(regs_10[7]), .Z(n_22883
		));
	notech_reg regs_reg_10_8(.CP(n_63510), .D(n_22889), .CD(n_62471), .Q(regs_10
		[8]));
	notech_mux2 i_4867(.S(n_442068004), .A(n_18572), .B(regs_10[8]), .Z(n_22889
		));
	notech_reg regs_reg_10_9(.CP(n_63510), .D(n_22895), .CD(n_62471), .Q(regs_10
		[9]));
	notech_mux2 i_4875(.S(n_442068004), .A(n_4354), .B(regs_10[9]), .Z(n_22895
		));
	notech_ao4 i_215641224(.A(n_58596), .B(n_31998), .C(n_58565), .D(n_31966
		), .Z(n_2606));
	notech_reg regs_reg_10_10(.CP(n_63510), .D(n_22901), .CD(n_62474), .Q(regs_10
		[10]));
	notech_mux2 i_4883(.S(n_442068004), .A(n_383864369), .B(regs_10[10]), .Z
		(n_22901));
	notech_ao4 i_215741223(.A(n_58574), .B(n_31410), .C(n_57524), .D(n_33129
		), .Z(n_2605));
	notech_reg regs_reg_10_11(.CP(n_63510), .D(n_22907), .CD(n_62474), .Q(regs_10
		[11]));
	notech_mux2 i_4891(.S(n_442068004), .A(n_437467958), .B(regs_10[11]), .Z
		(n_22907));
	notech_and2 i_216141219(.A(n_2603), .B(n_2602), .Z(n_2604));
	notech_reg regs_reg_10_12(.CP(n_63510), .D(n_22913), .CD(n_62474), .Q(regs_10
		[12]));
	notech_mux2 i_4899(.S(n_442068004), .A(n_437367957), .B(regs_10[12]), .Z
		(n_22913));
	notech_ao4 i_215941221(.A(n_57444), .B(n_31574), .C(n_57429), .D(n_31933
		), .Z(n_2603));
	notech_reg regs_reg_10_13(.CP(n_63510), .D(n_22919), .CD(n_62474), .Q(regs_10
		[13]));
	notech_mux2 i_4907(.S(n_442068004), .A(n_377464305), .B(regs_10[13]), .Z
		(n_22919));
	notech_ao4 i_216041220(.A(n_57412), .B(n_31901), .C(n_57406), .D(n_31869
		), .Z(n_2602));
	notech_reg regs_reg_10_14(.CP(n_63510), .D(n_22925), .CD(n_62474), .Q(regs_10
		[14]));
	notech_mux2 i_4915(.S(n_442068004), .A(n_18608), .B(regs_10[14]), .Z(n_22925
		));
	notech_and4 i_216941211(.A(n_2599), .B(n_2598), .C(n_259660491), .D(n_2595
		), .Z(n_2601));
	notech_reg regs_reg_10_15(.CP(n_63510), .D(n_22931), .CD(n_62476), .Q(regs_10
		[15]));
	notech_mux2 i_4923(.S(n_442068004), .A(n_437267956), .B(regs_10[15]), .Z
		(n_22931));
	notech_reg regs_reg_10_16(.CP(n_63510), .D(n_22937), .CD(n_62476), .Q(regs_10
		[16]));
	notech_mux2 i_4931(.S(n_55862), .A(n_18620), .B(regs_10[16]), .Z(n_22937
		));
	notech_ao4 i_216341217(.A(n_57512), .B(n_31837), .C(n_58550), .D(n_31805
		), .Z(n_2599));
	notech_reg regs_reg_10_17(.CP(n_63596), .D(n_22943), .CD(n_62475), .Q(regs_10
		[17]));
	notech_mux2 i_4939(.S(n_55862), .A(n_18626), .B(regs_10[17]), .Z(n_22943
		));
	notech_ao4 i_216441216(.A(n_57500), .B(n_31773), .C(n_57489), .D(n_31741
		), .Z(n_2598));
	notech_reg regs_reg_10_18(.CP(n_63596), .D(n_22949), .CD(n_62476), .Q(regs_10
		[18]));
	notech_mux2 i_4947(.S(n_55862), .A(n_18632), .B(regs_10[18]), .Z(n_22949
		));
	notech_reg regs_reg_10_19(.CP(n_63596), .D(n_22955), .CD(n_62476), .Q(regs_10
		[19]));
	notech_mux2 i_4955(.S(n_55862), .A(n_18638), .B(regs_10[19]), .Z(n_22955
		));
	notech_ao4 i_216641214(.A(n_57622), .B(n_33130), .C(n_57480), .D(n_31709
		), .Z(n_259660491));
	notech_reg regs_reg_10_20(.CP(n_63596), .D(n_22961), .CD(n_62476), .Q(regs_10
		[20]));
	notech_mux2 i_4963(.S(n_55862), .A(n_18644), .B(regs_10[20]), .Z(n_22961
		));
	notech_ao4 i_216741213(.A(n_57471), .B(n_31677), .C(n_57456), .D(n_31645
		), .Z(n_2595));
	notech_reg regs_reg_10_21(.CP(n_63596), .D(n_22969), .CD(n_62476), .Q(regs_10
		[21]));
	notech_mux2 i_4971(.S(n_55862), .A(n_18650), .B(regs_10[21]), .Z(n_22969
		));
	notech_reg regs_reg_10_22(.CP(n_63596), .D(n_22975), .CD(n_62476), .Q(regs_10
		[22]));
	notech_mux2 i_4979(.S(n_55862), .A(n_18656), .B(regs_10[22]), .Z(n_22975
		));
	notech_reg regs_reg_10_23(.CP(n_63596), .D(n_22987), .CD(n_62476), .Q(regs_10
		[23]));
	notech_mux2 i_4987(.S(n_55862), .A(n_18662), .B(regs_10[23]), .Z(n_22987
		));
	notech_ao4 i_217041210(.A(n_58596), .B(n_31996), .C(n_58565), .D(n_31964
		), .Z(n_2592));
	notech_reg regs_reg_10_24(.CP(n_63596), .D(n_22994), .CD(n_62475), .Q(regs_10
		[24]));
	notech_mux2 i_4995(.S(n_55862), .A(n_335281823), .B(regs_10[24]), .Z(n_22994
		));
	notech_ao4 i_217141209(.A(n_58574), .B(n_31408), .C(n_57524), .D(n_33134
		), .Z(n_2591));
	notech_reg regs_reg_10_25(.CP(n_63596), .D(n_23000), .CD(n_62475), .Q(regs_10
		[25]));
	notech_mux2 i_5003(.S(n_55862), .A(n_18674), .B(regs_10[25]), .Z(n_23000
		));
	notech_and2 i_217541205(.A(n_2589), .B(n_2588), .Z(n_2590));
	notech_reg regs_reg_10_26(.CP(n_63596), .D(n_23006), .CD(n_62475), .Q(regs_10
		[26]));
	notech_mux2 i_5011(.S(n_55862), .A(n_18680), .B(regs_10[26]), .Z(n_23006
		));
	notech_ao4 i_217341207(.A(n_57444), .B(n_31572), .C(n_57429), .D(n_31931
		), .Z(n_2589));
	notech_reg regs_reg_10_27(.CP(n_63596), .D(n_23012), .CD(n_62475), .Q(regs_10
		[27]));
	notech_mux2 i_5019(.S(n_55862), .A(n_18686), .B(regs_10[27]), .Z(n_23012
		));
	notech_ao4 i_217441206(.A(n_57412), .B(n_31899), .C(n_57406), .D(n_31867
		), .Z(n_2588));
	notech_reg regs_reg_10_28(.CP(n_63596), .D(n_23018), .CD(n_62475), .Q(regs_10
		[28]));
	notech_mux2 i_5027(.S(n_55862), .A(n_18692), .B(regs_10[28]), .Z(n_23018
		));
	notech_and4 i_218341197(.A(n_2585), .B(n_2584), .C(n_2582), .D(n_2581), 
		.Z(n_2587));
	notech_reg regs_reg_10_29(.CP(n_63596), .D(n_23026), .CD(n_62475), .Q(regs_10
		[29]));
	notech_mux2 i_5035(.S(n_55862), .A(n_4391), .B(regs_10[29]), .Z(n_23026)
		);
	notech_reg regs_reg_10_30(.CP(n_63596), .D(n_23032), .CD(n_62475), .Q(regs_10
		[30]));
	notech_mux2 i_5043(.S(n_55862), .A(n_18704), .B(regs_10[30]), .Z(n_23032
		));
	notech_ao4 i_217741203(.A(n_57512), .B(n_31835), .C(n_58550), .D(n_31803
		), .Z(n_2585));
	notech_reg regs_reg_10_31(.CP(n_63596), .D(n_23039), .CD(n_62475), .Q(regs_10
		[31]));
	notech_mux2 i_5051(.S(n_55862), .A(n_18710), .B(regs_10[31]), .Z(n_23039
		));
	notech_ao4 i_217841202(.A(n_57500), .B(n_31771), .C(n_57489), .D(n_31739
		), .Z(n_2584));
	notech_reg regs_reg_9_0(.CP(n_63596), .D(n_23045), .CD(n_62475), .Q(cs[0
		]));
	notech_mux2 i_5059(.S(n_157062602), .A(n_30925), .B(cs[0]), .Z(n_23045)
		);
	notech_reg regs_reg_9_1(.CP(n_63596), .D(n_23051), .CD(n_62475), .Q(cs[1
		]));
	notech_mux2 i_5067(.S(n_157062602), .A(n_16229), .B(cs[1]), .Z(n_23051)
		);
	notech_ao4 i_218041200(.A(n_57622), .B(n_31367), .C(n_57480), .D(n_31707
		), .Z(n_2582));
	notech_reg regs_reg_9_2(.CP(n_63596), .D(n_23057), .CD(n_62469), .Q(\nbus_14543[2] 
		));
	notech_mux2 i_5075(.S(n_157062602), .A(n_4359), .B(\nbus_14543[2] ), .Z(n_23057
		));
	notech_ao4 i_218141199(.A(n_57471), .B(n_31675), .C(n_57456), .D(n_31643
		), .Z(n_2581));
	notech_reg regs_reg_9_3(.CP(n_63596), .D(n_23063), .CD(n_62469), .Q(\nbus_14543[3] 
		));
	notech_mux2 i_5083(.S(n_157062602), .A(n_16241), .B(\nbus_14543[3] ), .Z
		(n_23063));
	notech_nand2 i_220441176(.A(n_61828), .B(n_61964), .Z(n_2580));
	notech_reg regs_reg_9_4(.CP(n_63664), .D(n_23069), .CD(n_62469), .Q(\nbus_14543[4] 
		));
	notech_mux2 i_5091(.S(n_157062602), .A(n_16247), .B(\nbus_14543[4] ), .Z
		(n_23069));
	notech_reg regs_reg_9_5(.CP(n_63594), .D(n_23075), .CD(n_62469), .Q(\nbus_14543[5] 
		));
	notech_mux2 i_5099(.S(n_157062602), .A(n_4370), .B(\nbus_14543[5] ), .Z(n_23075
		));
	notech_reg regs_reg_9_6(.CP(n_63664), .D(n_23081), .CD(n_62469), .Q(\nbus_14543[6] 
		));
	notech_mux2 i_5107(.S(n_157062602), .A(n_16259), .B(\nbus_14543[6] ), .Z
		(n_23081));
	notech_nand2 i_140243283(.A(n_61828), .B(n_61757), .Z(n_2577));
	notech_reg regs_reg_9_7(.CP(n_63664), .D(n_23087), .CD(n_62470), .Q(\nbus_14543[7] 
		));
	notech_mux2 i_5115(.S(n_157062602), .A(n_4358), .B(\nbus_14543[7] ), .Z(n_23087
		));
	notech_reg regs_reg_9_8(.CP(n_63664), .D(n_23093), .CD(n_62470), .Q(\nbus_14543[8] 
		));
	notech_mux2 i_5123(.S(n_157062602), .A(n_16271), .B(\nbus_14543[8] ), .Z
		(n_23093));
	notech_reg regs_reg_9_9(.CP(n_63664), .D(n_23099), .CD(n_62470), .Q(\nbus_14543[9] 
		));
	notech_mux2 i_5131(.S(n_157062602), .A(n_4357), .B(\nbus_14543[9] ), .Z(n_23099
		));
	notech_reg regs_reg_9_10(.CP(n_63664), .D(n_23105), .CD(n_62470), .Q(\nbus_14543[10] 
		));
	notech_mux2 i_5139(.S(n_157062602), .A(n_377564306), .B(\nbus_14543[10] 
		), .Z(n_23105));
	notech_reg regs_reg_9_11(.CP(n_63664), .D(n_23111), .CD(n_62469), .Q(\nbus_14543[11] 
		));
	notech_mux2 i_5147(.S(n_157062602), .A(n_437767961), .B(\nbus_14543[11] 
		), .Z(n_23111));
	notech_reg regs_reg_9_12(.CP(n_63664), .D(n_23117), .CD(n_62469), .Q(\nbus_14543[12] 
		));
	notech_mux2 i_5155(.S(n_157062602), .A(n_437667960), .B(\nbus_14543[12] 
		), .Z(n_23117));
	notech_reg regs_reg_9_13(.CP(n_63664), .D(n_23123), .CD(n_62469), .Q(\nbus_14543[13] 
		));
	notech_mux2 i_5163(.S(n_157062602), .A(n_16301), .B(\nbus_14543[13] ), .Z
		(n_23123));
	notech_reg regs_reg_9_14(.CP(n_63664), .D(n_23129), .CD(n_62468), .Q(\nbus_14543[14] 
		));
	notech_mux2 i_5171(.S(n_157062602), .A(n_16307), .B(\nbus_14543[14] ), .Z
		(n_23129));
	notech_reg regs_reg_9_15(.CP(n_63664), .D(n_23135), .CD(n_62468), .Q(\nbus_14543[15] 
		));
	notech_mux2 i_5179(.S(n_157062602), .A(n_437567959), .B(\nbus_14543[15] 
		), .Z(n_23135));
	notech_reg regs_reg_9_16(.CP(n_63664), .D(n_23141), .CD(n_62469), .Q(\nbus_14543[16] 
		));
	notech_mux2 i_5187(.S(n_57575), .A(n_16319), .B(\nbus_14543[16] ), .Z(n_23141
		));
	notech_reg regs_reg_9_17(.CP(n_63664), .D(n_23147), .CD(n_62469), .Q(\nbus_14543[17] 
		));
	notech_mux2 i_5195(.S(n_57575), .A(n_16325), .B(\nbus_14543[17] ), .Z(n_23147
		));
	notech_reg regs_reg_9_18(.CP(n_63664), .D(n_23153), .CD(n_62469), .Q(\nbus_14543[18] 
		));
	notech_mux2 i_5203(.S(n_57575), .A(n_16331), .B(\nbus_14543[18] ), .Z(n_23153
		));
	notech_reg regs_reg_9_19(.CP(n_63664), .D(n_23159), .CD(n_62469), .Q(\nbus_14543[19] 
		));
	notech_mux2 i_5211(.S(n_57575), .A(n_16337), .B(\nbus_14543[19] ), .Z(n_23159
		));
	notech_reg regs_reg_9_20(.CP(n_63664), .D(n_23165), .CD(n_62469), .Q(\nbus_14543[20] 
		));
	notech_mux2 i_5219(.S(n_57575), .A(n_16343), .B(\nbus_14543[20] ), .Z(n_23165
		));
	notech_reg regs_reg_9_21(.CP(n_63664), .D(n_23171), .CD(n_62471), .Q(\nbus_14543[21] 
		));
	notech_mux2 i_5227(.S(n_57575), .A(n_16349), .B(\nbus_14543[21] ), .Z(n_23171
		));
	notech_reg regs_reg_9_22(.CP(n_63664), .D(n_23177), .CD(n_62471), .Q(\nbus_14543[22] 
		));
	notech_mux2 i_5235(.S(n_57575), .A(n_16355), .B(\nbus_14543[22] ), .Z(n_23177
		));
	notech_reg regs_reg_9_23(.CP(n_63664), .D(n_23183), .CD(n_62471), .Q(\nbus_14543[23] 
		));
	notech_mux2 i_5243(.S(n_57575), .A(n_16361), .B(\nbus_14543[23] ), .Z(n_23183
		));
	notech_reg regs_reg_9_24(.CP(n_63594), .D(n_23189), .CD(n_62471), .Q(\nbus_14543[24] 
		));
	notech_mux2 i_5251(.S(n_57575), .A(n_16367), .B(\nbus_14543[24] ), .Z(n_23189
		));
	notech_reg regs_reg_9_25(.CP(n_63594), .D(n_23195), .CD(n_62471), .Q(\nbus_14543[25] 
		));
	notech_mux2 i_5259(.S(n_57575), .A(n_16373), .B(\nbus_14543[25] ), .Z(n_23195
		));
	notech_reg regs_reg_9_26(.CP(n_63594), .D(n_23201), .CD(n_62471), .Q(\nbus_14543[26] 
		));
	notech_mux2 i_5267(.S(n_57575), .A(n_16379), .B(\nbus_14543[26] ), .Z(n_23201
		));
	notech_reg regs_reg_9_27(.CP(n_63594), .D(n_23207), .CD(n_62471), .Q(\nbus_14543[27] 
		));
	notech_mux2 i_5275(.S(n_57575), .A(n_16385), .B(\nbus_14543[27] ), .Z(n_23207
		));
	notech_reg regs_reg_9_28(.CP(n_63594), .D(n_23213), .CD(n_62471), .Q(\nbus_14543[28] 
		));
	notech_mux2 i_5283(.S(n_57575), .A(n_16391), .B(\nbus_14543[28] ), .Z(n_23213
		));
	notech_reg regs_reg_9_29(.CP(n_63594), .D(n_23219), .CD(n_62471), .Q(\nbus_14543[29] 
		));
	notech_mux2 i_5291(.S(n_57575), .A(n_30927), .B(\nbus_14543[29] ), .Z(n_23219
		));
	notech_reg regs_reg_9_30(.CP(n_63594), .D(n_23225), .CD(n_62471), .Q(\nbus_14543[30] 
		));
	notech_mux2 i_5299(.S(n_57575), .A(n_16403), .B(\nbus_14543[30] ), .Z(n_23225
		));
	notech_reg regs_reg_9_31(.CP(n_63594), .D(n_23231), .CD(n_62470), .Q(\nbus_14543[31] 
		));
	notech_mux2 i_5307(.S(n_57575), .A(n_16409), .B(\nbus_14543[31] ), .Z(n_23231
		));
	notech_reg regs_reg_8_0(.CP(n_63594), .D(n_23237), .CD(n_62470), .Q(regs_8
		[0]));
	notech_mux2 i_5315(.S(n_389964430), .A(n_30660), .B(regs_8[0]), .Z(n_23237
		));
	notech_reg regs_reg_8_1(.CP(n_63594), .D(n_23243), .CD(n_62470), .Q(regs_8
		[1]));
	notech_mux2 i_5323(.S(n_389964430), .A(n_379964330), .B(regs_8[1]), .Z(n_23243
		));
	notech_reg regs_reg_8_2(.CP(n_63510), .D(n_23249), .CD(n_62470), .Q(regs_8
		[2]));
	notech_mux2 i_5331(.S(n_389964430), .A(n_178662814), .B(regs_8[2]), .Z(n_23249
		));
	notech_reg regs_reg_8_3(.CP(n_63510), .D(n_23255), .CD(n_62470), .Q(regs_8
		[3]));
	notech_mux2 i_5339(.S(n_389964430), .A(n_388564416), .B(regs_8[3]), .Z(n_23255
		));
	notech_reg regs_reg_8_4(.CP(n_63598), .D(n_23261), .CD(n_62470), .Q(regs_8
		[4]));
	notech_mux2 i_5347(.S(n_389964430), .A(n_384164372), .B(regs_8[4]), .Z(n_23261
		));
	notech_reg regs_reg_8_5(.CP(n_63512), .D(n_23267), .CD(n_62470), .Q(regs_8
		[5]));
	notech_mux2 i_5355(.S(n_389964430), .A(n_379864329), .B(regs_8[5]), .Z(n_23267
		));
	notech_reg regs_reg_8_6(.CP(n_63512), .D(n_23273), .CD(n_62470), .Q(regs_8
		[6]));
	notech_mux2 i_5363(.S(n_389964430), .A(n_177262800), .B(regs_8[6]), .Z(n_23273
		));
	notech_reg regs_reg_8_7(.CP(n_63512), .D(n_23279), .CD(n_62470), .Q(regs_8
		[7]));
	notech_mux2 i_5371(.S(n_389964430), .A(n_175962787), .B(regs_8[7]), .Z(n_23279
		));
	notech_reg regs_reg_8_8(.CP(n_63512), .D(n_23285), .CD(n_62481), .Q(regs_8
		[8]));
	notech_mux2 i_5379(.S(n_389964430), .A(n_13388), .B(regs_8[8]), .Z(n_23285
		));
	notech_reg regs_reg_8_9(.CP(n_63512), .D(n_23291), .CD(n_62481), .Q(regs_8
		[9]));
	notech_mux2 i_5387(.S(n_389964430), .A(n_210666516), .B(regs_8[9]), .Z(n_23291
		));
	notech_reg regs_reg_8_10(.CP(n_63512), .D(n_23297), .CD(n_62481), .Q(regs_8
		[10]));
	notech_mux2 i_5395(.S(n_389964430), .A(n_384064371), .B(regs_8[10]), .Z(n_23297
		));
	notech_reg regs_reg_8_11(.CP(n_63512), .D(n_23303), .CD(n_62481), .Q(regs_8
		[11]));
	notech_mux2 i_5403(.S(n_389964430), .A(n_209366505), .B(regs_8[11]), .Z(n_23303
		));
	notech_reg regs_reg_8_12(.CP(n_63512), .D(n_23309), .CD(n_62481), .Q(regs_8
		[12]));
	notech_mux2 i_5411(.S(n_389964430), .A(n_208066494), .B(regs_8[12]), .Z(n_23309
		));
	notech_reg regs_reg_8_13(.CP(n_63512), .D(n_23315), .CD(n_62481), .Q(regs_8
		[13]));
	notech_mux2 i_5419(.S(n_389964430), .A(n_174662774), .B(regs_8[13]), .Z(n_23315
		));
	notech_reg regs_reg_8_14(.CP(n_63512), .D(n_23321), .CD(n_62481), .Q(regs_8
		[14]));
	notech_mux2 i_5427(.S(n_389964430), .A(n_173562763), .B(regs_8[14]), .Z(n_23321
		));
	notech_reg regs_reg_8_15(.CP(n_63598), .D(n_23328), .CD(n_62481), .Q(regs_8
		[15]));
	notech_mux2 i_5435(.S(n_389964430), .A(n_206566483), .B(regs_8[15]), .Z(n_23328
		));
	notech_reg regs_reg_8_16(.CP(n_63598), .D(n_23337), .CD(n_62481), .Q(regs_8
		[16]));
	notech_mux2 i_5443(.S(n_55873), .A(n_13436), .B(regs_8[16]), .Z(n_23337)
		);
	notech_reg regs_reg_8_17(.CP(n_63598), .D(n_23344), .CD(n_62480), .Q(regs_8
		[17]));
	notech_mux2 i_5451(.S(n_55873), .A(n_13442), .B(regs_8[17]), .Z(n_23344)
		);
	notech_reg regs_reg_8_18(.CP(n_63598), .D(n_23354), .CD(n_62480), .Q(regs_8
		[18]));
	notech_mux2 i_5459(.S(n_55873), .A(n_13448), .B(regs_8[18]), .Z(n_23354)
		);
	notech_reg regs_reg_8_19(.CP(n_63598), .D(n_23361), .CD(n_62480), .Q(regs_8
		[19]));
	notech_mux2 i_5468(.S(n_55873), .A(n_388464415), .B(regs_8[19]), .Z(n_23361
		));
	notech_reg regs_reg_8_20(.CP(n_63598), .D(n_23368), .CD(n_62480), .Q(regs_8
		[20]));
	notech_mux2 i_5476(.S(n_55873), .A(n_3013), .B(regs_8[20]), .Z(n_23368)
		);
	notech_reg regs_reg_8_21(.CP(n_63598), .D(n_23376), .CD(n_62480), .Q(regs_8
		[21]));
	notech_mux2 i_5484(.S(n_55873), .A(n_3004), .B(regs_8[21]), .Z(n_23376)
		);
	notech_reg regs_reg_8_22(.CP(n_63598), .D(n_23384), .CD(n_62480), .Q(regs_8
		[22]));
	notech_mux2 i_5492(.S(n_55873), .A(n_2995), .B(regs_8[22]), .Z(n_23384)
		);
	notech_reg regs_reg_8_23(.CP(n_63598), .D(n_23392), .CD(n_62480), .Q(regs_8
		[23]));
	notech_mux2 i_5500(.S(n_55873), .A(n_298663884), .B(regs_8[23]), .Z(n_23392
		));
	notech_reg regs_reg_8_24(.CP(n_63598), .D(n_23398), .CD(n_62480), .Q(regs_8
		[24]));
	notech_mux2 i_5508(.S(n_55873), .A(n_297763875), .B(regs_8[24]), .Z(n_23398
		));
	notech_reg regs_reg_8_25(.CP(n_63598), .D(n_23404), .CD(n_62480), .Q(regs_8
		[25]));
	notech_mux2 i_5516(.S(n_55873), .A(n_296863866), .B(regs_8[25]), .Z(n_23404
		));
	notech_reg regs_reg_8_26(.CP(n_63598), .D(n_23410), .CD(n_62480), .Q(regs_8
		[26]));
	notech_mux2 i_5524(.S(n_55873), .A(n_13496), .B(regs_8[26]), .Z(n_23410)
		);
	notech_reg regs_reg_8_27(.CP(n_63598), .D(n_23416), .CD(n_62482), .Q(regs_8
		[27]));
	notech_mux2 i_5532(.S(n_55873), .A(n_13502), .B(regs_8[27]), .Z(n_23416)
		);
	notech_reg regs_reg_8_28(.CP(n_63598), .D(n_23422), .CD(n_62482), .Q(regs_8
		[28]));
	notech_mux2 i_5540(.S(n_55873), .A(n_13508), .B(regs_8[28]), .Z(n_23422)
		);
	notech_reg regs_reg_8_29(.CP(n_63598), .D(n_23428), .CD(n_62482), .Q(regs_8
		[29]));
	notech_mux2 i_5548(.S(n_55873), .A(n_30405), .B(regs_8[29]), .Z(n_23428)
		);
	notech_reg regs_reg_8_30(.CP(n_63598), .D(n_23434), .CD(n_62482), .Q(regs_8
		[30]));
	notech_mux2 i_5556(.S(n_55873), .A(n_13520), .B(regs_8[30]), .Z(n_23434)
		);
	notech_reg regs_reg_8_31(.CP(n_63598), .D(n_23440), .CD(n_62482), .Q(regs_8
		[31]));
	notech_mux2 i_5564(.S(n_55873), .A(n_13526), .B(regs_8[31]), .Z(n_23440)
		);
	notech_reg regs_reg_7_0(.CP(n_63598), .D(n_23446), .CD(n_62482), .Q(regs_7
		[0]));
	notech_mux2 i_5572(.S(n_30918), .A(n_30928), .B(regs_7[0]), .Z(n_23446)
		);
	notech_reg regs_reg_7_1(.CP(n_63512), .D(n_23452), .CD(n_62482), .Q(regs_7
		[1]));
	notech_mux2 i_5580(.S(n_30918), .A(n_30929), .B(regs_7[1]), .Z(n_23452)
		);
	notech_reg regs_reg_7_2(.CP(n_63512), .D(n_23458), .CD(n_62482), .Q(regs_7
		[2]));
	notech_mux2 i_5588(.S(n_30918), .A(n_30445), .B(regs_7[2]), .Z(n_23458)
		);
	notech_reg regs_reg_7_3(.CP(n_63514), .D(n_23464), .CD(n_62482), .Q(regs_7
		[3]));
	notech_mux2 i_5596(.S(n_30918), .A(n_30411), .B(regs_7[3]), .Z(n_23464)
		);
	notech_reg regs_reg_7_4(.CP(n_63514), .D(n_23470), .CD(n_62482), .Q(regs_7
		[4]));
	notech_mux2 i_5604(.S(n_30918), .A(n_30930), .B(regs_7[4]), .Z(n_23470)
		);
	notech_reg regs_reg_7_5(.CP(n_63514), .D(n_23476), .CD(n_62481), .Q(regs_7
		[5]));
	notech_mux2 i_5612(.S(n_30918), .A(n_30931), .B(regs_7[5]), .Z(n_23476)
		);
	notech_reg regs_reg_7_6(.CP(n_63514), .D(n_23482), .CD(n_62481), .Q(regs_7
		[6]));
	notech_mux2 i_5620(.S(n_30918), .A(n_30932), .B(regs_7[6]), .Z(n_23482)
		);
	notech_reg regs_reg_7_7(.CP(n_63514), .D(n_23488), .CD(n_62481), .Q(regs_7
		[7]));
	notech_mux2 i_5628(.S(n_30918), .A(n_30933), .B(regs_7[7]), .Z(n_23488)
		);
	notech_reg regs_reg_7_8(.CP(n_63514), .D(n_23494), .CD(n_62481), .Q(regs_7
		[8]));
	notech_mux2 i_5636(.S(n_30918), .A(n_15922), .B(regs_7[8]), .Z(n_23494)
		);
	notech_reg regs_reg_7_9(.CP(n_63514), .D(n_23500), .CD(n_62481), .Q(regs_7
		[9]));
	notech_mux2 i_5644(.S(n_30918), .A(n_4360), .B(regs_7[9]), .Z(n_23500)
		);
	notech_reg regs_reg_7_10(.CP(n_63514), .D(n_23506), .CD(n_62482), .Q(regs_7
		[10]));
	notech_mux2 i_5652(.S(n_30918), .A(n_377764308), .B(regs_7[10]), .Z(n_23506
		));
	notech_reg regs_reg_7_11(.CP(n_63514), .D(n_23516), .CD(n_62482), .Q(regs_7
		[11]));
	notech_mux2 i_5660(.S(n_30918), .A(n_438067964), .B(regs_7[11]), .Z(n_23516
		));
	notech_reg regs_reg_7_12(.CP(n_63514), .D(n_23525), .CD(n_62482), .Q(regs_7
		[12]));
	notech_mux2 i_5668(.S(n_30918), .A(n_437967963), .B(regs_7[12]), .Z(n_23525
		));
	notech_reg regs_reg_7_13(.CP(n_63514), .D(n_23531), .CD(n_62482), .Q(regs_7
		[13]));
	notech_mux2 i_5676(.S(n_30918), .A(n_377664307), .B(regs_7[13]), .Z(n_23531
		));
	notech_reg regs_reg_7_14(.CP(n_63514), .D(n_23537), .CD(n_62477), .Q(regs_7
		[14]));
	notech_mux2 i_5684(.S(n_30918), .A(n_30934), .B(regs_7[14]), .Z(n_23537)
		);
	notech_reg regs_reg_7_15(.CP(n_63514), .D(n_23543), .CD(n_62477), .Q(regs_7
		[15]));
	notech_mux2 i_5692(.S(n_30918), .A(n_437867962), .B(regs_7[15]), .Z(n_23543
		));
	notech_reg regs_reg_7_16(.CP(n_63514), .D(n_23549), .CD(n_62477), .Q(regs_7
		[16]));
	notech_mux2 i_5700(.S(n_55893), .A(n_15970), .B(regs_7[16]), .Z(n_23549)
		);
	notech_reg regs_reg_7_17(.CP(n_63514), .D(n_23555), .CD(n_62477), .Q(regs_7
		[17]));
	notech_mux2 i_5708(.S(n_55893), .A(n_15976), .B(regs_7[17]), .Z(n_23555)
		);
	notech_reg regs_reg_7_18(.CP(n_63514), .D(n_23561), .CD(n_62477), .Q(regs_7
		[18]));
	notech_mux2 i_5716(.S(n_55893), .A(n_15982), .B(regs_7[18]), .Z(n_23561)
		);
	notech_reg regs_reg_7_19(.CP(n_63514), .D(n_23567), .CD(n_62477), .Q(regs_7
		[19]));
	notech_mux2 i_5724(.S(n_55893), .A(n_15988), .B(regs_7[19]), .Z(n_23567)
		);
	notech_reg regs_reg_7_20(.CP(n_63514), .D(n_23573), .CD(n_62477), .Q(regs_7
		[20]));
	notech_mux2 i_5732(.S(n_55893), .A(n_15994), .B(regs_7[20]), .Z(n_23573)
		);
	notech_reg regs_reg_7_21(.CP(n_63514), .D(n_23579), .CD(n_62477), .Q(regs_7
		[21]));
	notech_mux2 i_5740(.S(n_55893), .A(n_16000), .B(regs_7[21]), .Z(n_23579)
		);
	notech_reg regs_reg_7_22(.CP(n_63458), .D(n_23585), .CD(n_62477), .Q(regs_7
		[22]));
	notech_mux2 i_5748(.S(n_55893), .A(n_16006), .B(regs_7[22]), .Z(n_23585)
		);
	notech_reg regs_reg_7_23(.CP(n_63458), .D(n_23591), .CD(n_62477), .Q(regs_7
		[23]));
	notech_mux2 i_5756(.S(n_55893), .A(n_1923), .B(regs_7[23]), .Z(n_23591)
		);
	notech_reg regs_reg_7_24(.CP(n_63458), .D(n_23597), .CD(n_62476), .Q(regs_7
		[24]));
	notech_mux2 i_5764(.S(n_55893), .A(n_351567679), .B(regs_7[24]), .Z(n_23597
		));
	notech_reg regs_reg_7_25(.CP(n_63458), .D(n_23603), .CD(n_62476), .Q(regs_7
		[25]));
	notech_mux2 i_5772(.S(n_55893), .A(n_350167666), .B(regs_7[25]), .Z(n_23603
		));
	notech_reg regs_reg_7_26(.CP(n_63458), .D(n_23609), .CD(n_62476), .Q(regs_7
		[26]));
	notech_mux2 i_5780(.S(n_55893), .A(n_16030), .B(regs_7[26]), .Z(n_23609)
		);
	notech_reg regs_reg_7_27(.CP(n_63458), .D(n_23619), .CD(n_62476), .Q(regs_7
		[27]));
	notech_mux2 i_5788(.S(n_55893), .A(n_16036), .B(regs_7[27]), .Z(n_23619)
		);
	notech_reg regs_reg_7_28(.CP(n_63458), .D(n_23625), .CD(n_62476), .Q(regs_7
		[28]));
	notech_mux2 i_5796(.S(n_55893), .A(n_16042), .B(regs_7[28]), .Z(n_23625)
		);
	notech_reg regs_reg_7_29(.CP(n_63458), .D(n_23631), .CD(n_62477), .Q(regs_7
		[29]));
	notech_mux2 i_5804(.S(n_55893), .A(n_4393), .B(regs_7[29]), .Z(n_23631)
		);
	notech_reg regs_reg_7_30(.CP(n_63458), .D(n_23637), .CD(n_62477), .Q(regs_7
		[30]));
	notech_mux2 i_5813(.S(n_55893), .A(n_16054), .B(regs_7[30]), .Z(n_23637)
		);
	notech_reg regs_reg_7_31(.CP(n_63458), .D(n_23643), .CD(n_62476), .Q(regs_7
		[31]));
	notech_mux2 i_5821(.S(n_55893), .A(n_16060), .B(regs_7[31]), .Z(n_23643)
		);
	notech_reg pipe_mul_reg_0(.CP(n_63508), .D(n_23649), .CD(n_62477), .Q(pipe_mul
		[0]));
	notech_mux2 i_5829(.S(\nbus_11285[0] ), .A(pipe_mul[0]), .B(n_315492473)
		, .Z(n_23649));
	notech_reg pipe_mul_reg_1(.CP(n_63498), .D(n_23655), .CD(n_62479), .Q(pipe_mul
		[1]));
	notech_mux2 i_5837(.S(\nbus_11285[0] ), .A(pipe_mul[1]), .B(n_315592474)
		, .Z(n_23655));
	notech_reg CFOF_mul_reg(.CP(n_63498), .D(n_23661), .CD(n_62479), .Q(CFOF_mul
		));
	notech_mux2 i_5845(.S(n_365728697), .A(CFOF_mul), .B(n_8438), .Z(n_23661
		));
	notech_reg eval_flag_reg(.CP(n_63498), .D(n_23667), .CD(n_62479), .Q(eval_flag
		));
	notech_mux2 i_5853(.S(n_11366), .A(eval_flag), .B(n_230691660), .Z(n_23667
		));
	notech_reg rep_en1_reg(.CP(n_63498), .D(n_23673), .CD(n_62479), .Q(rep_en1
		));
	notech_mux2 i_5861(.S(n_8771), .A(rep_en1), .B(n_61661), .Z(n_23673));
	notech_reg rep_en2_reg(.CP(n_63498), .D(n_23679), .CD(n_62479), .Q(rep_en2
		));
	notech_mux2 i_5870(.S(n_8589), .A(rep_en2), .B(n_61661), .Z(n_23679));
	notech_reg rep_en3_reg(.CP(n_63498), .D(n_23685), .CD(n_62480), .Q(rep_en3
		));
	notech_mux2 i_5881(.S(n_10054), .A(rep_en3), .B(n_61665), .Z(n_23685));
	notech_reg rep_en4_reg(.CP(n_63498), .D(n_23691), .CD(n_62480), .Q(rep_en4
		));
	notech_mux2 i_5889(.S(n_14525), .A(rep_en4), .B(n_61661), .Z(n_23691));
	notech_reg rep_en5_reg(.CP(n_63498), .D(n_23697), .CD(n_62480), .Q(rep_en5
		));
	notech_mux2 i_5897(.S(n_10088), .A(rep_en5), .B(n_61661), .Z(n_23697));
	notech_reg nCF_reg(.CP(n_63498), .D(n_23703), .CD(n_62480), .Q(nCF));
	notech_mux2 i_5905(.S(n_30940), .A(nCF), .B(n_7418), .Z(n_23703));
	notech_reg nPF_reg(.CP(n_63498), .D(n_23709), .CD(n_62479), .Q(nPF));
	notech_mux2 i_5914(.S(n_30941), .A(nPF), .B(n_302392361), .Z(n_23709));
	notech_reg nAF_reg(.CP(n_63498), .D(n_23715), .CD(n_62479), .Q(nAF));
	notech_mux2 i_5922(.S(n_30944), .A(nAF), .B(nAF_arithbox), .Z(n_23715)
		);
	notech_reg nSF_reg(.CP(n_63498), .D(n_23721), .CD(n_62479), .Q(nSF));
	notech_mux2 i_5930(.S(n_223991593), .A(n_30424), .B(nSF), .Z(n_23721));
	notech_reg opas_reg(.CP(n_63574), .D(n_23727), .CD(n_62477), .Q(opas));
	notech_mux2 i_5938(.S(n_30944), .A(opas), .B(opas_arithbox), .Z(n_23727)
		);
	notech_reg opbs_reg(.CP(n_63574), .D(n_23733), .CD(n_62479), .Q(opbs));
	notech_mux2 i_5946(.S(n_30944), .A(opbs), .B(opbs_arithbox), .Z(n_23733)
		);
	notech_reg nOF_reg(.CP(n_63574), .D(n_23739), .CD(n_62479), .Q(nOF));
	notech_mux2 i_5954(.S(n_30946), .A(nOF), .B(n_30945), .Z(n_23739));
	notech_reg regs_reg_15_0(.CP(n_63574), .D(n_23748), .CD(n_62479), .Q(\eflags[0] 
		));
	notech_mux2 i_5962(.S(\nbus_11352[0] ), .A(\eflags[0] ), .B(n_30947), .Z
		(n_23748));
	notech_reg regs_reg_15_1(.CP(n_63574), .D(n_23756), .CD(n_62479), .Q(\eflags[1] 
		));
	notech_mux2 i_5970(.S(\nbus_11352[1] ), .A(\eflags[1] ), .B(n_20390), .Z
		(n_23756));
	notech_reg regs_reg_15_2(.CP(n_63574), .D(n_23766), .CD(n_62479), .Q(\eflags[2] 
		));
	notech_mux2 i_5978(.S(\nbus_11352[2] ), .A(\eflags[2] ), .B(n_20396), .Z
		(n_23766));
	notech_reg regs_reg_15_3(.CP(n_63574), .D(n_23772), .CD(n_62479), .Q(\eflags[3] 
		));
	notech_mux2 i_5986(.S(\nbus_11352[1] ), .A(\eflags[3] ), .B(n_20402), .Z
		(n_23772));
	notech_reg regs_reg_15_4(.CP(n_63574), .D(n_23778), .CD(n_62458), .Q(\eflags[4] 
		));
	notech_mux2 i_5994(.S(\nbus_11352[0] ), .A(\eflags[4] ), .B(n_20408), .Z
		(n_23778));
	notech_reg regs_reg_15_5(.CP(n_63574), .D(n_23784), .CD(n_62458), .Q(\eflags[5] 
		));
	notech_mux2 i_6002(.S(\nbus_11352[1] ), .A(\eflags[5] ), .B(n_4379), .Z(n_23784
		));
	notech_reg regs_reg_15_6(.CP(n_63574), .D(n_23790), .CD(n_62457), .Q(\eflags[6] 
		));
	notech_mux2 i_6010(.S(\nbus_11352[6] ), .A(\eflags[6] ), .B(n_30948), .Z
		(n_23790));
	notech_reg regs_reg_15_7(.CP(n_63574), .D(n_23796), .CD(n_62457), .Q(\eflags[7] 
		));
	notech_mux2 i_6018(.S(\nbus_11352[6] ), .A(\eflags[7] ), .B(n_30396), .Z
		(n_23796));
	notech_reg regs_reg_15_8(.CP(n_63574), .D(n_23802), .CD(n_62458), .Q(\eflags[8] 
		));
	notech_mux2 i_6026(.S(\nbus_11352[8] ), .A(\eflags[8] ), .B(n_20432), .Z
		(n_23802));
	notech_reg regs_reg_15_9(.CP(n_63574), .D(n_23808), .CD(n_62458), .Q(ie)
		);
	notech_mux2 i_6034(.S(n_30949), .A(ie), .B(n_20438), .Z(n_23808));
	notech_reg regs_reg_15_10(.CP(n_63574), .D(n_23814), .CD(n_62458), .Q(\eflags[10] 
		));
	notech_mux2 i_6042(.S(\nbus_11352[10] ), .A(\eflags[10] ), .B(n_377964310
		), .Z(n_23814));
	notech_reg regs_reg_15_11(.CP(n_63574), .D(n_23820), .CD(n_62458), .Q(\eflags[11] 
		));
	notech_mux2 i_6050(.S(\nbus_11352[6] ), .A(\eflags[11] ), .B(n_447168055
		), .Z(n_23820));
	notech_reg regs_reg_15_12(.CP(n_63574), .D(n_23826), .CD(n_62458), .Q(\eflags[12] 
		));
	notech_mux2 i_6058(.S(n_179766229), .A(n_30443), .B(\eflags[12] ), .Z(n_23826
		));
	notech_reg regs_reg_15_13(.CP(n_63574), .D(n_23832), .CD(n_62457), .Q(\eflags[13] 
		));
	notech_mux2 i_6066(.S(n_179766229), .A(n_30659), .B(\eflags[13] ), .Z(n_23832
		));
	notech_reg regs_reg_15_14(.CP(n_63574), .D(n_23840), .CD(n_62457), .Q(\eflags[14] 
		));
	notech_mux2 i_6074(.S(n_179766229), .A(n_20468), .B(\eflags[14] ), .Z(n_23840
		));
	notech_reg regs_reg_15_15(.CP(n_63574), .D(n_23849), .CD(n_62457), .Q(\eflags[15] 
		));
	notech_mux2 i_6082(.S(\nbus_11352[1] ), .A(\eflags[15] ), .B(n_30444), .Z
		(n_23849));
	notech_reg regs_reg_15_16(.CP(n_63572), .D(n_23855), .CD(n_62457), .Q(\eflags[16] 
		));
	notech_mux2 i_6090(.S(n_179766229), .A(n_20480), .B(\eflags[16] ), .Z(n_23855
		));
	notech_reg regs_reg_15_17(.CP(n_63572), .D(n_23861), .CD(n_62457), .Q(\eflags[17] 
		));
	notech_mux2 i_6098(.S(n_179766229), .A(n_20486), .B(\eflags[17] ), .Z(n_23861
		));
	notech_reg regs_reg_15_18(.CP(n_63648), .D(n_23867), .CD(n_62457), .Q(\eflags[18] 
		));
	notech_mux2 i_6106(.S(n_179766229), .A(n_20492), .B(\eflags[18] ), .Z(n_23867
		));
	notech_reg regs_reg_15_19(.CP(n_63648), .D(n_23874), .CD(n_62457), .Q(\eflags[19] 
		));
	notech_mux2 i_6114(.S(n_179766229), .A(n_20498), .B(\eflags[19] ), .Z(n_23874
		));
	notech_reg regs_reg_15_20(.CP(n_63648), .D(n_23880), .CD(n_62457), .Q(\eflags[20] 
		));
	notech_mux2 i_6122(.S(n_179766229), .A(n_20504), .B(\eflags[20] ), .Z(n_23880
		));
	notech_reg regs_reg_15_21(.CP(n_63648), .D(n_23886), .CD(n_62457), .Q(\eflags[21] 
		));
	notech_mux2 i_6130(.S(n_179766229), .A(n_20510), .B(\eflags[21] ), .Z(n_23886
		));
	notech_reg regs_reg_15_22(.CP(n_63648), .D(n_23892), .CD(n_62457), .Q(\eflags[22] 
		));
	notech_mux2 i_6138(.S(n_179766229), .A(n_20516), .B(\eflags[22] ), .Z(n_23892
		));
	notech_reg regs_reg_15_23(.CP(n_63648), .D(n_23898), .CD(n_62459), .Q(\eflags[23] 
		));
	notech_mux2 i_6146(.S(n_179766229), .A(n_20522), .B(\eflags[23] ), .Z(n_23898
		));
	notech_reg regs_reg_15_24(.CP(n_63648), .D(n_23904), .CD(n_62459), .Q(\eflags[24] 
		));
	notech_mux2 i_6154(.S(n_179766229), .A(n_20528), .B(\eflags[24] ), .Z(n_23904
		));
	notech_reg regs_reg_15_25(.CP(n_63648), .D(n_23910), .CD(n_62459), .Q(\eflags[25] 
		));
	notech_mux2 i_6162(.S(n_179766229), .A(n_20534), .B(\eflags[25] ), .Z(n_23910
		));
	notech_reg regs_reg_15_26(.CP(n_63648), .D(n_23916), .CD(n_62459), .Q(\eflags[26] 
		));
	notech_mux2 i_6170(.S(n_179766229), .A(n_20540), .B(\eflags[26] ), .Z(n_23916
		));
	notech_reg regs_reg_15_27(.CP(n_63648), .D(n_23922), .CD(n_62459), .Q(\eflags[27] 
		));
	notech_mux2 i_6178(.S(n_179766229), .A(n_20546), .B(\eflags[27] ), .Z(n_23922
		));
	notech_reg regs_reg_15_28(.CP(n_63648), .D(n_23928), .CD(n_62459), .Q(\eflags[28] 
		));
	notech_mux2 i_6186(.S(n_179766229), .A(n_20552), .B(\eflags[28] ), .Z(n_23928
		));
	notech_reg regs_reg_15_29(.CP(n_63648), .D(n_23934), .CD(n_62459), .Q(\eflags[29] 
		));
	notech_mux2 i_6194(.S(n_179766229), .A(n_20558), .B(\eflags[29] ), .Z(n_23934
		));
	notech_reg regs_reg_15_30(.CP(n_63648), .D(n_23940), .CD(n_62459), .Q(\eflags[30] 
		));
	notech_mux2 i_6202(.S(n_179766229), .A(n_20564), .B(\eflags[30] ), .Z(n_23940
		));
	notech_reg regs_reg_15_31(.CP(n_63648), .D(n_23946), .CD(n_62459), .Q(\eflags[31] 
		));
	notech_mux2 i_6210(.S(n_179766229), .A(n_20570), .B(\eflags[31] ), .Z(n_23946
		));
	notech_reg regs_reg_6_0(.CP(n_63648), .D(n_23952), .CD(n_62459), .Q(regs_6
		[0]));
	notech_mux2 i_6218(.S(n_30961), .A(regs_6[0]), .B(n_30951), .Z(n_23952)
		);
	notech_reg regs_reg_6_1(.CP(n_63648), .D(n_23958), .CD(n_62458), .Q(regs_6
		[1]));
	notech_mux2 i_6226(.S(n_30961), .A(regs_6[1]), .B(n_30952), .Z(n_23958)
		);
	notech_reg regs_reg_6_2(.CP(n_63648), .D(n_23964), .CD(n_62458), .Q(regs_6
		[2]));
	notech_mux2 i_6234(.S(n_30961), .A(regs_6[2]), .B(n_30953), .Z(n_23964)
		);
	notech_reg regs_reg_6_3(.CP(n_63648), .D(n_23970), .CD(n_62458), .Q(regs_6
		[3]));
	notech_mux2 i_6242(.S(n_30961), .A(regs_6[3]), .B(n_30954), .Z(n_23970)
		);
	notech_reg regs_reg_6_4(.CP(n_63572), .D(n_23976), .CD(n_62458), .Q(regs_6
		[4]));
	notech_mux2 i_6250(.S(n_30961), .A(regs_6[4]), .B(n_30955), .Z(n_23976)
		);
	notech_reg regs_reg_6_5(.CP(n_63572), .D(n_23982), .CD(n_62458), .Q(regs_6
		[5]));
	notech_mux2 i_6258(.S(n_30961), .A(regs_6[5]), .B(n_30956), .Z(n_23982)
		);
	notech_reg regs_reg_6_6(.CP(n_63572), .D(n_23990), .CD(n_62459), .Q(regs_6
		[6]));
	notech_mux2 i_6266(.S(n_30961), .A(regs_6[6]), .B(n_30957), .Z(n_23990)
		);
	notech_reg regs_reg_6_7(.CP(n_63572), .D(n_23996), .CD(n_62459), .Q(regs_6
		[7]));
	notech_mux2 i_6274(.S(n_30961), .A(regs_6[7]), .B(n_30958), .Z(n_23996)
		);
	notech_reg regs_reg_6_8(.CP(n_63572), .D(n_24003), .CD(n_62458), .Q(regs_6
		[8]));
	notech_mux2 i_6282(.S(n_30961), .A(regs_6[8]), .B(n_15570), .Z(n_24003)
		);
	notech_reg regs_reg_6_9(.CP(n_63572), .D(n_24009), .CD(n_62459), .Q(regs_6
		[9]));
	notech_mux2 i_6291(.S(n_30961), .A(regs_6[9]), .B(n_15576), .Z(n_24009)
		);
	notech_reg regs_reg_6_10(.CP(n_63572), .D(n_24015), .CD(n_62454), .Q(regs_6
		[10]));
	notech_mux2 i_6299(.S(n_30961), .A(regs_6[10]), .B(n_378164312), .Z(n_24015
		));
	notech_reg regs_reg_6_11(.CP(n_63572), .D(n_24021), .CD(n_62454), .Q(regs_6
		[11]));
	notech_mux2 i_6307(.S(n_30961), .A(regs_6[11]), .B(n_438667970), .Z(n_24021
		));
	notech_reg regs_reg_6_12(.CP(n_63572), .D(n_24027), .CD(n_62453), .Q(regs_6
		[12]));
	notech_mux2 i_6315(.S(n_30961), .A(regs_6[12]), .B(n_438567969), .Z(n_24027
		));
	notech_reg regs_reg_6_13(.CP(n_63572), .D(n_24033), .CD(n_62454), .Q(regs_6
		[13]));
	notech_mux2 i_6323(.S(n_30961), .A(regs_6[13]), .B(n_378064311), .Z(n_24033
		));
	notech_reg regs_reg_6_14(.CP(n_63648), .D(n_24039), .CD(n_62454), .Q(regs_6
		[14]));
	notech_mux2 i_6331(.S(n_30961), .A(regs_6[14]), .B(n_30959), .Z(n_24039)
		);
	notech_reg regs_reg_6_15(.CP(n_63570), .D(n_24045), .CD(n_62454), .Q(regs_6
		[15]));
	notech_mux2 i_6339(.S(n_30961), .A(regs_6[15]), .B(n_438467968), .Z(n_24045
		));
	notech_reg regs_reg_6_16(.CP(n_63570), .D(n_24051), .CD(n_62454), .Q(regs_6
		[16]));
	notech_mux2 i_6348(.S(n_55924), .A(regs_6[16]), .B(n_15618), .Z(n_24051)
		);
	notech_reg regs_reg_6_17(.CP(n_63644), .D(n_24057), .CD(n_62454), .Q(regs_6
		[17]));
	notech_mux2 i_6356(.S(n_55924), .A(regs_6[17]), .B(n_15624), .Z(n_24057)
		);
	notech_reg regs_reg_6_18(.CP(n_63644), .D(n_24063), .CD(n_62454), .Q(regs_6
		[18]));
	notech_mux2 i_6364(.S(n_55924), .A(regs_6[18]), .B(n_15630), .Z(n_24063)
		);
	notech_reg regs_reg_6_19(.CP(n_63644), .D(n_24069), .CD(n_62453), .Q(regs_6
		[19]));
	notech_mux2 i_6372(.S(n_55924), .A(regs_6[19]), .B(n_15636), .Z(n_24069)
		);
	notech_reg regs_reg_6_20(.CP(n_63644), .D(n_24075), .CD(n_62453), .Q(regs_6
		[20]));
	notech_mux2 i_6380(.S(n_55924), .A(regs_6[20]), .B(n_15642), .Z(n_24075)
		);
	notech_reg regs_reg_6_21(.CP(n_63644), .D(n_24081), .CD(n_62453), .Q(regs_6
		[21]));
	notech_mux2 i_6388(.S(n_55924), .A(regs_6[21]), .B(n_15648), .Z(n_24081)
		);
	notech_reg regs_reg_6_22(.CP(n_63644), .D(n_24087), .CD(n_62453), .Q(regs_6
		[22]));
	notech_mux2 i_6396(.S(n_55924), .A(regs_6[22]), .B(n_15654), .Z(n_24087)
		);
	notech_reg regs_reg_6_23(.CP(n_63644), .D(n_24093), .CD(n_62453), .Q(regs_6
		[23]));
	notech_mux2 i_6404(.S(n_55924), .A(regs_6[23]), .B(n_15660), .Z(n_24093)
		);
	notech_reg regs_reg_6_24(.CP(n_63644), .D(n_24099), .CD(n_62453), .Q(regs_6
		[24]));
	notech_mux2 i_6413(.S(n_55924), .A(regs_6[24]), .B(n_1936), .Z(n_24099)
		);
	notech_reg regs_reg_6_25(.CP(n_63644), .D(n_24105), .CD(n_62453), .Q(regs_6
		[25]));
	notech_mux2 i_6421(.S(n_55924), .A(regs_6[25]), .B(n_15672), .Z(n_24105)
		);
	notech_reg regs_reg_6_26(.CP(n_63644), .D(n_24111), .CD(n_62453), .Q(regs_6
		[26]));
	notech_mux2 i_6429(.S(n_55924), .A(regs_6[26]), .B(n_15678), .Z(n_24111)
		);
	notech_reg regs_reg_6_27(.CP(n_63686), .D(n_24117), .CD(n_62453), .Q(regs_6
		[27]));
	notech_mux2 i_6437(.S(n_55924), .A(regs_6[27]), .B(n_15684), .Z(n_24117)
		);
	notech_reg regs_reg_6_28(.CP(n_63686), .D(n_24123), .CD(n_62453), .Q(regs_6
		[28]));
	notech_mux2 i_6445(.S(n_55924), .A(regs_6[28]), .B(n_15690), .Z(n_24123)
		);
	notech_reg regs_reg_6_29(.CP(n_63686), .D(n_24130), .CD(n_62455), .Q(regs_6
		[29]));
	notech_mux2 i_6453(.S(n_55924), .A(regs_6[29]), .B(n_15696), .Z(n_24130)
		);
	notech_reg regs_reg_6_30(.CP(n_63686), .D(n_24139), .CD(n_62455), .Q(regs_6
		[30]));
	notech_mux2 i_6461(.S(n_55924), .A(regs_6[30]), .B(n_15702), .Z(n_24139)
		);
	notech_reg regs_reg_6_31(.CP(n_63686), .D(n_24150), .CD(n_62455), .Q(regs_6
		[31]));
	notech_mux2 i_6469(.S(n_55924), .A(regs_6[31]), .B(n_15708), .Z(n_24150)
		);
	notech_reg regs_reg_5_0(.CP(n_63686), .D(n_24156), .CD(n_62455), .Q(regs_5
		[0]));
	notech_mux2 i_6477(.S(n_164362675), .A(n_1567), .B(regs_5[0]), .Z(n_24156
		));
	notech_reg regs_reg_5_1(.CP(n_63686), .D(n_24162), .CD(n_62455), .Q(regs_5
		[1]));
	notech_mux2 i_6485(.S(n_164362675), .A(n_380264333), .B(regs_5[1]), .Z(n_24162
		));
	notech_reg regs_reg_5_2(.CP(n_63686), .D(n_24168), .CD(n_62455), .Q(regs_5
		[2]));
	notech_mux2 i_6493(.S(n_164362675), .A(n_187262899), .B(regs_5[2]), .Z(n_24168
		));
	notech_reg regs_reg_5_3(.CP(n_63686), .D(n_24174), .CD(n_62457), .Q(regs_5
		[3]));
	notech_mux2 i_6501(.S(n_164362675), .A(n_389064421), .B(regs_5[3]), .Z(n_24174
		));
	notech_reg regs_reg_5_4(.CP(n_63686), .D(n_24180), .CD(n_62455), .Q(regs_5
		[4]));
	notech_mux2 i_6509(.S(n_164362675), .A(n_384264373), .B(regs_5[4]), .Z(n_24180
		));
	notech_reg regs_reg_5_5(.CP(n_63686), .D(n_24186), .CD(n_62455), .Q(regs_5
		[5]));
	notech_mux2 i_6517(.S(n_164362675), .A(n_380164332), .B(regs_5[5]), .Z(n_24186
		));
	notech_reg regs_reg_5_6(.CP(n_63686), .D(n_24192), .CD(n_62455), .Q(regs_5
		[6]));
	notech_mux2 i_6525(.S(n_164362675), .A(n_185862885), .B(regs_5[6]), .Z(n_24192
		));
	notech_reg regs_reg_5_7(.CP(n_63686), .D(n_24198), .CD(n_62454), .Q(regs_5
		[7]));
	notech_mux2 i_6533(.S(n_164362675), .A(n_184462872), .B(regs_5[7]), .Z(n_24198
		));
	notech_reg regs_reg_5_8(.CP(n_63686), .D(n_24204), .CD(n_62454), .Q(regs_5
		[8]));
	notech_mux2 i_6541(.S(n_164362675), .A(n_13040), .B(regs_5[8]), .Z(n_24204
		));
	notech_reg regs_reg_5_9(.CP(n_63686), .D(n_24210), .CD(n_62454), .Q(regs_5
		[9]));
	notech_mux2 i_6549(.S(n_164362675), .A(n_1556), .B(regs_5[9]), .Z(n_24210
		));
	notech_reg regs_reg_5_10(.CP(n_63686), .D(n_24217), .CD(n_62454), .Q(regs_5
		[10]));
	notech_mux2 i_6557(.S(n_164362675), .A(n_183162859), .B(regs_5[10]), .Z(n_24217
		));
	notech_reg regs_reg_5_11(.CP(n_63686), .D(n_24223), .CD(n_62454), .Q(regs_5
		[11]));
	notech_mux2 i_6565(.S(n_164362675), .A(n_213966549), .B(regs_5[11]), .Z(n_24223
		));
	notech_reg regs_reg_5_12(.CP(n_63686), .D(n_24231), .CD(n_62455), .Q(regs_5
		[12]));
	notech_mux2 i_6573(.S(n_164362675), .A(n_212866538), .B(regs_5[12]), .Z(n_24231
		));
	notech_reg regs_reg_5_13(.CP(n_63644), .D(n_24237), .CD(n_62455), .Q(regs_5
		[13]));
	notech_mux2 i_6581(.S(n_164362675), .A(n_182062848), .B(regs_5[13]), .Z(n_24237
		));
	notech_reg regs_reg_5_14(.CP(n_63686), .D(n_24243), .CD(n_62455), .Q(regs_5
		[14]));
	notech_mux2 i_6589(.S(n_164362675), .A(n_180962837), .B(regs_5[14]), .Z(n_24243
		));
	notech_reg regs_reg_5_15(.CP(n_63646), .D(n_24249), .CD(n_62455), .Q(regs_5
		[15]));
	notech_mux2 i_6597(.S(n_164362675), .A(n_211766527), .B(regs_5[15]), .Z(n_24249
		));
	notech_reg regs_reg_5_16(.CP(n_63646), .D(n_24255), .CD(n_62465), .Q(regs_5
		[16]));
	notech_mux2 i_6605(.S(n_55935), .A(n_388964420), .B(regs_5[16]), .Z(n_24255
		));
	notech_reg regs_reg_5_17(.CP(n_63646), .D(n_24261), .CD(n_62465), .Q(regs_5
		[17]));
	notech_mux2 i_6613(.S(n_55935), .A(n_388864419), .B(regs_5[17]), .Z(n_24261
		));
	notech_reg regs_reg_5_18(.CP(n_63646), .D(n_24267), .CD(n_62465), .Q(regs_5
		[18]));
	notech_mux2 i_6621(.S(n_55935), .A(n_388764418), .B(regs_5[18]), .Z(n_24267
		));
	notech_reg regs_reg_5_19(.CP(n_63646), .D(n_24273), .CD(n_62465), .Q(regs_5
		[19]));
	notech_mux2 i_6629(.S(n_55935), .A(n_388664417), .B(regs_5[19]), .Z(n_24273
		));
	notech_reg regs_reg_5_20(.CP(n_63646), .D(n_24279), .CD(n_62466), .Q(regs_5
		[20]));
	notech_mux2 i_6637(.S(n_55935), .A(n_13112), .B(regs_5[20]), .Z(n_24279)
		);
	notech_reg regs_reg_5_21(.CP(n_63646), .D(n_24285), .CD(n_62466), .Q(regs_5
		[21]));
	notech_mux2 i_6645(.S(n_55935), .A(n_13118), .B(regs_5[21]), .Z(n_24285)
		);
	notech_reg regs_reg_5_22(.CP(n_63646), .D(n_24291), .CD(n_62466), .Q(regs_5
		[22]));
	notech_mux2 i_6653(.S(n_55935), .A(n_13124), .B(regs_5[22]), .Z(n_24291)
		);
	notech_reg regs_reg_5_23(.CP(n_63646), .D(n_24297), .CD(n_62466), .Q(regs_5
		[23]));
	notech_mux2 i_6661(.S(n_55935), .A(n_13130), .B(regs_5[23]), .Z(n_24297)
		);
	notech_reg regs_reg_5_24(.CP(n_63646), .D(n_24306), .CD(n_62466), .Q(regs_5
		[24]));
	notech_mux2 i_6669(.S(n_55935), .A(n_13136), .B(regs_5[24]), .Z(n_24306)
		);
	notech_or2 i_181243276(.A(n_61828), .B(n_32160), .Z(n_2383));
	notech_reg regs_reg_5_25(.CP(n_63646), .D(n_24312), .CD(n_62465), .Q(regs_5
		[25]));
	notech_mux2 i_6677(.S(n_55935), .A(n_3022), .B(regs_5[25]), .Z(n_24312)
		);
	notech_nand2 i_152543280(.A(n_61786), .B(n_61944), .Z(n_2382));
	notech_reg regs_reg_5_26(.CP(n_63646), .D(n_24318), .CD(n_62465), .Q(regs_5
		[26]));
	notech_mux2 i_6685(.S(n_55935), .A(n_387464405), .B(regs_5[26]), .Z(n_24318
		));
	notech_reg regs_reg_5_27(.CP(n_63646), .D(n_24324), .CD(n_62465), .Q(regs_5
		[27]));
	notech_mux2 i_6693(.S(n_55935), .A(n_387364404), .B(regs_5[27]), .Z(n_24324
		));
	notech_reg regs_reg_5_28(.CP(n_63646), .D(n_24330), .CD(n_62464), .Q(regs_5
		[28]));
	notech_mux2 i_6701(.S(n_55935), .A(n_387264403), .B(regs_5[28]), .Z(n_24330
		));
	notech_ao4 i_203544479(.A(n_57117), .B(n_31780), .C(n_57609), .D(n_33132
		), .Z(n_2379));
	notech_reg regs_reg_5_29(.CP(n_63646), .D(n_24336), .CD(n_62465), .Q(regs_5
		[29]));
	notech_mux2 i_6709(.S(n_55935), .A(n_30641), .B(regs_5[29]), .Z(n_24336)
		);
	notech_ao4 i_203644478(.A(n_57136), .B(n_31748), .C(n_57157), .D(n_33131
		), .Z(n_2378));
	notech_reg regs_reg_5_30(.CP(n_63646), .D(n_24342), .CD(n_62465), .Q(regs_5
		[30]));
	notech_mux2 i_6717(.S(n_55935), .A(n_380064331), .B(regs_5[30]), .Z(n_24342
		));
	notech_and2 i_204044474(.A(n_2376), .B(n_2375), .Z(n_2377));
	notech_reg regs_reg_5_31(.CP(n_63646), .D(n_24348), .CD(n_62465), .Q(regs_5
		[31]));
	notech_mux2 i_6725(.S(n_55935), .A(n_389564426), .B(regs_5[31]), .Z(n_24348
		));
	notech_ao4 i_203844476(.A(n_57163), .B(n_31844), .C(n_57178), .D(n_32005
		), .Z(n_2376));
	notech_reg sav_cs_reg_0(.CP(n_63646), .D(n_24354), .CD(n_62465), .Q(sav_cs
		[0]));
	notech_mux2 i_6733(.S(n_59599), .A(cs[0]), .B(sav_cs[0]), .Z(n_24354));
	notech_ao4 i_203944475(.A(n_57189), .B(n_31716), .C(n_57199), .D(n_31940
		), .Z(n_2375));
	notech_reg sav_cs_reg_1(.CP(n_63646), .D(n_24360), .CD(n_62465), .Q(sav_cs
		[1]));
	notech_mux2 i_6741(.S(n_59599), .A(cs[1]), .B(sav_cs[1]), .Z(n_24360));
	notech_and4 i_204844466(.A(n_2372), .B(n_2371), .C(n_2369), .D(n_2368), 
		.Z(n_2374));
	notech_reg tss_esp0_reg(.CP(n_63570), .D(n_24366), .CD(n_62465), .Q(tss_esp0
		));
	notech_mux2 i_6749(.S(n_14184), .A(tss_esp0), .B(n_61661), .Z(n_24366)
		);
	notech_reg_set temp_sp_reg_0(.CP(n_63570), .D(n_24372), .SD(1'b1), .Q(temp_sp
		[0]));
	notech_mux2 i_6757(.S(\nbus_11320[0] ), .A(temp_sp[0]), .B(n_30966), .Z(n_24372
		));
	notech_ao4 i_204244472(.A(n_57059), .B(n_31684), .C(n_57072), .D(n_31812
		), .Z(n_2372));
	notech_reg_set temp_sp_reg_1(.CP(n_63570), .D(n_24378), .SD(1'b1), .Q(temp_sp
		[1]));
	notech_mux2 i_6765(.S(\nbus_11320[0] ), .A(temp_sp[1]), .B(n_30968), .Z(n_24378
		));
	notech_ao4 i_204344471(.A(n_57086), .B(n_31876), .C(n_57097), .D(n_31581
		), .Z(n_2371));
	notech_reg_set temp_sp_reg_2(.CP(n_63570), .D(n_24384), .SD(1'b1), .Q(temp_sp
		[2]));
	notech_mux2 i_6773(.S(\nbus_11320[0] ), .A(temp_sp[2]), .B(n_30970), .Z(n_24384
		));
	notech_reg_set temp_sp_reg_3(.CP(n_63570), .D(n_24390), .SD(1'b1), .Q(temp_sp
		[3]));
	notech_mux2 i_6781(.S(\nbus_11320[0] ), .A(temp_sp[3]), .B(n_30972), .Z(n_24390
		));
	notech_ao4 i_204544469(.A(n_58696), .B(n_31973), .C(n_59095), .D(n_31908
		), .Z(n_2369));
	notech_reg_set temp_sp_reg_4(.CP(n_63570), .D(n_24396), .SD(1'b1), .Q(temp_sp
		[4]));
	notech_mux2 i_6789(.S(\nbus_11320[0] ), .A(temp_sp[4]), .B(n_30974), .Z(n_24396
		));
	notech_ao4 i_204644468(.A(n_57211), .B(n_31417), .C(n_57225), .D(n_31652
		), .Z(n_2368));
	notech_reg_set temp_sp_reg_5(.CP(n_63570), .D(n_24402), .SD(1'b1), .Q(temp_sp
		[5]));
	notech_mux2 i_6797(.S(\nbus_11320[0] ), .A(temp_sp[5]), .B(n_30976), .Z(n_24402
		));
	notech_reg_set temp_sp_reg_6(.CP(n_63570), .D(n_24408), .SD(1'b1), .Q(temp_sp
		[6]));
	notech_mux2 i_6805(.S(\nbus_11320[0] ), .A(temp_sp[6]), .B(n_30978), .Z(n_24408
		));
	notech_reg_set temp_sp_reg_7(.CP(n_63570), .D(n_24414), .SD(1'b1), .Q(temp_sp
		[7]));
	notech_mux2 i_6813(.S(\nbus_11320[0] ), .A(temp_sp[7]), .B(n_30980), .Z(n_24414
		));
	notech_ao4 i_205044464(.A(n_57117), .B(n_31772), .C(n_57609), .D(n_31368
		), .Z(n_2365));
	notech_reg_set temp_sp_reg_8(.CP(n_63570), .D(n_24420), .SD(1'b1), .Q(temp_sp
		[8]));
	notech_mux2 i_6821(.S(\nbus_11320[0] ), .A(temp_sp[8]), .B(n_30982), .Z(n_24420
		));
	notech_ao4 i_205144463(.A(n_57136), .B(n_31740), .C(n_57157), .D(n_33133
		), .Z(n_2364));
	notech_reg_set temp_sp_reg_9(.CP(n_63644), .D(n_24433), .SD(1'b1), .Q(temp_sp
		[9]));
	notech_mux2 i_6829(.S(\nbus_11320[0] ), .A(temp_sp[9]), .B(n_30984), .Z(n_24433
		));
	notech_and2 i_205544459(.A(n_2362), .B(n_2361), .Z(n_2363));
	notech_reg_set temp_sp_reg_10(.CP(n_63638), .D(n_24439), .SD(1'b1), .Q(temp_sp
		[10]));
	notech_mux2 i_6837(.S(\nbus_11320[0] ), .A(temp_sp[10]), .B(n_30986), .Z
		(n_24439));
	notech_ao4 i_205344461(.A(n_57163), .B(n_31836), .C(n_57178), .D(n_31997
		), .Z(n_2362));
	notech_reg_set temp_sp_reg_11(.CP(n_63638), .D(n_24445), .SD(1'b1), .Q(temp_sp
		[11]));
	notech_mux2 i_6845(.S(\nbus_11320[0] ), .A(temp_sp[11]), .B(n_30988), .Z
		(n_24445));
	notech_ao4 i_205444460(.A(n_57189), .B(n_31708), .C(n_57199), .D(n_31932
		), .Z(n_2361));
	notech_reg_set temp_sp_reg_12(.CP(n_63638), .D(n_24451), .SD(1'b1), .Q(temp_sp
		[12]));
	notech_mux2 i_6853(.S(\nbus_11320[0] ), .A(temp_sp[12]), .B(n_30990), .Z
		(n_24451));
	notech_and4 i_206344451(.A(n_2358), .B(n_2357), .C(n_2355), .D(n_2354), 
		.Z(n_2360));
	notech_reg_set temp_sp_reg_13(.CP(n_63638), .D(n_24457), .SD(1'b1), .Q(temp_sp
		[13]));
	notech_mux2 i_6861(.S(\nbus_11320[0] ), .A(temp_sp[13]), .B(n_30992), .Z
		(n_24457));
	notech_reg_set temp_sp_reg_14(.CP(n_63638), .D(n_24463), .SD(1'b1), .Q(temp_sp
		[14]));
	notech_mux2 i_6869(.S(\nbus_11320[0] ), .A(temp_sp[14]), .B(n_30994), .Z
		(n_24463));
	notech_ao4 i_205744457(.A(n_57059), .B(n_31676), .C(n_57072), .D(n_31804
		), .Z(n_2358));
	notech_reg_set temp_sp_reg_15(.CP(n_63638), .D(n_24469), .SD(1'b1), .Q(temp_sp
		[15]));
	notech_mux2 i_6877(.S(\nbus_11320[0] ), .A(temp_sp[15]), .B(n_30996), .Z
		(n_24469));
	notech_ao4 i_205844456(.A(n_57086), .B(n_31868), .C(n_57097), .D(n_31573
		), .Z(n_2357));
	notech_reg_set temp_sp_reg_16(.CP(n_63638), .D(n_24475), .SD(1'b1), .Q(temp_sp
		[16]));
	notech_mux2 i_6885(.S(n_55599), .A(temp_sp[16]), .B(n_30998), .Z(n_24475
		));
	notech_reg_set temp_sp_reg_17(.CP(n_63638), .D(n_24481), .SD(1'b1), .Q(temp_sp
		[17]));
	notech_mux2 i_6893(.S(n_55599), .A(temp_sp[17]), .B(n_31001), .Z(n_24481
		));
	notech_ao4 i_206044454(.A(n_58701), .B(n_31965), .C(n_59095), .D(n_31900
		), .Z(n_2355));
	notech_reg_set temp_sp_reg_18(.CP(n_63638), .D(n_24487), .SD(1'b1), .Q(temp_sp
		[18]));
	notech_mux2 i_6901(.S(n_55599), .A(temp_sp[18]), .B(n_31003), .Z(n_24487
		));
	notech_ao4 i_206144453(.A(n_57211), .B(n_31409), .C(n_57225), .D(n_31644
		), .Z(n_2354));
	notech_reg_set temp_sp_reg_19(.CP(n_63638), .D(n_24493), .SD(1'b1), .Q(temp_sp
		[19]));
	notech_mux2 i_6909(.S(n_55599), .A(temp_sp[19]), .B(n_31005), .Z(n_24493
		));
	notech_reg_set temp_sp_reg_20(.CP(n_63638), .D(n_24499), .SD(1'b1), .Q(temp_sp
		[20]));
	notech_mux2 i_6917(.S(n_55599), .A(temp_sp[20]), .B(n_31007), .Z(n_24499
		));
	notech_reg_set temp_sp_reg_21(.CP(n_63638), .D(n_24505), .SD(1'b1), .Q(temp_sp
		[21]));
	notech_mux2 i_6925(.S(n_55599), .A(temp_sp[21]), .B(n_31009), .Z(n_24505
		));
	notech_ao4 i_206444450(.A(n_57117), .B(n_31771), .C(n_57609), .D(n_31367
		), .Z(n_2351));
	notech_reg_set temp_sp_reg_22(.CP(n_63682), .D(n_24511), .SD(1'b1), .Q(temp_sp
		[22]));
	notech_mux2 i_6933(.S(n_55599), .A(temp_sp[22]), .B(n_31011), .Z(n_24511
		));
	notech_ao4 i_206544449(.A(n_57136), .B(n_31739), .C(n_57152), .D(n_33134
		), .Z(n_2350));
	notech_reg_set temp_sp_reg_23(.CP(n_63682), .D(n_24517), .SD(1'b1), .Q(temp_sp
		[23]));
	notech_mux2 i_6941(.S(n_55599), .A(temp_sp[23]), .B(n_31013), .Z(n_24517
		));
	notech_and2 i_206944445(.A(n_2348), .B(n_2347), .Z(n_2349));
	notech_reg_set temp_sp_reg_24(.CP(n_63682), .D(n_24523), .SD(1'b1), .Q(temp_sp
		[24]));
	notech_mux2 i_6949(.S(n_55599), .A(temp_sp[24]), .B(n_31015), .Z(n_24523
		));
	notech_ao4 i_206744447(.A(n_57163), .B(n_31835), .C(n_57178), .D(n_31996
		), .Z(n_2348));
	notech_reg_set temp_sp_reg_25(.CP(n_63682), .D(n_24531), .SD(1'b1), .Q(temp_sp
		[25]));
	notech_mux2 i_6957(.S(n_55599), .A(temp_sp[25]), .B(n_31017), .Z(n_24531
		));
	notech_ao4 i_206844446(.A(n_57189), .B(n_31707), .C(n_57199), .D(n_31931
		), .Z(n_2347));
	notech_reg_set temp_sp_reg_26(.CP(n_63682), .D(n_24537), .SD(1'b1), .Q(temp_sp
		[26]));
	notech_mux2 i_6965(.S(n_55599), .A(temp_sp[26]), .B(n_31019), .Z(n_24537
		));
	notech_and4 i_207744437(.A(n_2344), .B(n_2343), .C(n_2341), .D(n_2340), 
		.Z(n_2346));
	notech_reg_set temp_sp_reg_27(.CP(n_63682), .D(n_24546), .SD(1'b1), .Q(temp_sp
		[27]));
	notech_mux2 i_6973(.S(n_55599), .A(temp_sp[27]), .B(n_31021), .Z(n_24546
		));
	notech_reg_set temp_sp_reg_28(.CP(n_63682), .D(n_24552), .SD(1'b1), .Q(temp_sp
		[28]));
	notech_mux2 i_6981(.S(n_55599), .A(temp_sp[28]), .B(n_31023), .Z(n_24552
		));
	notech_ao4 i_207144443(.A(n_57059), .B(n_31675), .C(n_57072), .D(n_31803
		), .Z(n_2344));
	notech_reg_set temp_sp_reg_29(.CP(n_63682), .D(n_24558), .SD(1'b1), .Q(temp_sp
		[29]));
	notech_mux2 i_6989(.S(n_55599), .A(temp_sp[29]), .B(n_31025), .Z(n_24558
		));
	notech_ao4 i_207244442(.A(n_57086), .B(n_31867), .C(n_57097), .D(n_31572
		), .Z(n_2343));
	notech_reg_set temp_sp_reg_30(.CP(n_63682), .D(n_24564), .SD(1'b1), .Q(temp_sp
		[30]));
	notech_mux2 i_6997(.S(n_55599), .A(temp_sp[30]), .B(n_31027), .Z(n_24564
		));
	notech_reg_set temp_sp_reg_31(.CP(n_63682), .D(n_24570), .SD(1'b1), .Q(temp_sp
		[31]));
	notech_mux2 i_7005(.S(n_55599), .A(temp_sp[31]), .B(n_31029), .Z(n_24570
		));
	notech_ao4 i_207444440(.A(n_58701), .B(n_31964), .C(n_59095), .D(n_31899
		), .Z(n_2341));
	notech_reg regs_reg_4_0(.CP(n_63682), .D(n_24576), .CD(n_62468), .Q(regs_4
		[0]));
	notech_mux2 i_7013(.S(n_445582455), .A(n_31031), .B(regs_4[0]), .Z(n_24576
		));
	notech_ao4 i_207544439(.A(n_57211), .B(n_31408), .C(n_57225), .D(n_31643
		), .Z(n_2340));
	notech_reg regs_reg_4_1(.CP(n_63682), .D(n_24582), .CD(n_62468), .Q(regs_4
		[1]));
	notech_mux2 i_7021(.S(n_445582455), .A(n_15176), .B(regs_4[1]), .Z(n_24582
		));
	notech_reg regs_reg_4_2(.CP(n_63682), .D(n_24588), .CD(n_62468), .Q(regs_4
		[2]));
	notech_mux2 i_7030(.S(n_445582455), .A(n_30442), .B(regs_4[2]), .Z(n_24588
		));
	notech_reg regs_reg_4_3(.CP(n_63682), .D(n_24594), .CD(n_62468), .Q(regs_4
		[3]));
	notech_mux2 i_7038(.S(n_445582455), .A(n_30905), .B(regs_4[3]), .Z(n_24594
		));
	notech_reg regs_reg_4_4(.CP(n_63682), .D(n_24600), .CD(n_62468), .Q(regs_4
		[4]));
	notech_mux2 i_7046(.S(n_445582455), .A(n_31032), .B(regs_4[4]), .Z(n_24600
		));
	notech_reg regs_reg_4_5(.CP(n_63682), .D(n_24606), .CD(n_62468), .Q(regs_4
		[5]));
	notech_mux2 i_7054(.S(n_445582455), .A(n_31033), .B(regs_4[5]), .Z(n_24606
		));
	notech_reg regs_reg_4_6(.CP(n_63682), .D(n_24612), .CD(n_62468), .Q(regs_4
		[6]));
	notech_mux2 i_7062(.S(n_445582455), .A(n_31034), .B(regs_4[6]), .Z(n_24612
		));
	notech_reg regs_reg_4_7(.CP(n_63682), .D(n_24618), .CD(n_62468), .Q(regs_4
		[7]));
	notech_mux2 i_7070(.S(n_445582455), .A(n_31035), .B(regs_4[7]), .Z(n_24618
		));
	notech_reg regs_reg_4_8(.CP(n_63682), .D(n_24624), .CD(n_62468), .Q(regs_4
		[8]));
	notech_mux2 i_7078(.S(n_445582455), .A(n_15218), .B(regs_4[8]), .Z(n_24624
		));
	notech_reg regs_reg_4_9(.CP(n_63694), .D(n_24630), .CD(n_62468), .Q(regs_4
		[9]));
	notech_mux2 i_7086(.S(n_445582455), .A(n_436282448), .B(regs_4[9]), .Z(n_24630
		));
	notech_reg regs_reg_4_10(.CP(n_63694), .D(n_24636), .CD(n_62466), .Q(regs_4
		[10]));
	notech_mux2 i_7094(.S(n_445582455), .A(n_378264313), .B(regs_4[10]), .Z(n_24636
		));
	notech_reg regs_reg_4_11(.CP(n_63694), .D(n_24642), .CD(n_62466), .Q(regs_4
		[11]));
	notech_mux2 i_7102(.S(n_445582455), .A(n_438967973), .B(regs_4[11]), .Z(n_24642
		));
	notech_reg regs_reg_4_12(.CP(n_63694), .D(n_24648), .CD(n_62466), .Q(regs_4
		[12]));
	notech_mux2 i_7110(.S(n_445582455), .A(n_438867972), .B(regs_4[12]), .Z(n_24648
		));
	notech_reg regs_reg_4_13(.CP(n_63694), .D(n_24654), .CD(n_62466), .Q(regs_4
		[13]));
	notech_mux2 i_7118(.S(n_445582455), .A(n_391564446), .B(regs_4[13]), .Z(n_24654
		));
	notech_reg regs_reg_4_14(.CP(n_63694), .D(n_24660), .CD(n_62466), .Q(regs_4
		[14]));
	notech_mux2 i_7126(.S(n_445582455), .A(n_15254), .B(regs_4[14]), .Z(n_24660
		));
	notech_reg regs_reg_4_15(.CP(n_63694), .D(n_24666), .CD(n_62466), .Q(regs_4
		[15]));
	notech_mux2 i_7134(.S(n_445582455), .A(n_438767971), .B(regs_4[15]), .Z(n_24666
		));
	notech_reg regs_reg_4_16(.CP(n_63694), .D(n_24672), .CD(n_62468), .Q(regs_4
		[16]));
	notech_mux2 i_7142(.S(n_55986), .A(n_4415), .B(regs_4[16]), .Z(n_24672)
		);
	notech_reg regs_reg_4_17(.CP(n_63694), .D(n_24678), .CD(n_62466), .Q(regs_4
		[17]));
	notech_mux2 i_7150(.S(n_55986), .A(n_4414), .B(regs_4[17]), .Z(n_24678)
		);
	notech_reg regs_reg_4_18(.CP(n_63694), .D(n_24684), .CD(n_62466), .Q(regs_4
		[18]));
	notech_mux2 i_7158(.S(n_55986), .A(n_4413), .B(regs_4[18]), .Z(n_24684)
		);
	notech_reg regs_reg_4_19(.CP(n_63694), .D(n_24690), .CD(n_62460), .Q(regs_4
		[19]));
	notech_mux2 i_7166(.S(n_55986), .A(n_4412), .B(regs_4[19]), .Z(n_24690)
		);
	notech_reg regs_reg_4_20(.CP(n_63694), .D(n_24696), .CD(n_62463), .Q(regs_4
		[20]));
	notech_mux2 i_7174(.S(n_55986), .A(n_15290), .B(regs_4[20]), .Z(n_24696)
		);
	notech_reg regs_reg_4_21(.CP(n_63694), .D(n_24702), .CD(n_62460), .Q(regs_4
		[21]));
	notech_mux2 i_7182(.S(n_55986), .A(n_15296), .B(regs_4[21]), .Z(n_24702)
		);
	notech_reg regs_reg_4_22(.CP(n_63694), .D(n_24708), .CD(n_62460), .Q(regs_4
		[22]));
	notech_mux2 i_7190(.S(n_55986), .A(n_15302), .B(regs_4[22]), .Z(n_24708)
		);
	notech_reg regs_reg_4_23(.CP(n_63694), .D(n_24714), .CD(n_62463), .Q(regs_4
		[23]));
	notech_mux2 i_7198(.S(n_55986), .A(n_15308), .B(regs_4[23]), .Z(n_24714)
		);
	notech_reg regs_reg_4_24(.CP(n_63694), .D(n_24722), .CD(n_62463), .Q(regs_4
		[24]));
	notech_mux2 i_7206(.S(n_55986), .A(n_352967693), .B(regs_4[24]), .Z(n_24722
		));
	notech_reg regs_reg_4_25(.CP(n_63694), .D(n_24730), .CD(n_62463), .Q(regs_4
		[25]));
	notech_mux2 i_7214(.S(n_55986), .A(n_1950), .B(regs_4[25]), .Z(n_24730)
		);
	notech_reg regs_reg_4_26(.CP(n_63694), .D(n_24739), .CD(n_62463), .Q(regs_4
		[26]));
	notech_mux2 i_7222(.S(n_55986), .A(n_4397), .B(regs_4[26]), .Z(n_24739)
		);
	notech_reg regs_reg_4_27(.CP(n_63694), .D(n_24745), .CD(n_62463), .Q(regs_4
		[27]));
	notech_mux2 i_7230(.S(n_55986), .A(n_4396), .B(regs_4[27]), .Z(n_24745)
		);
	notech_reg regs_reg_4_28(.CP(n_63694), .D(n_24751), .CD(n_62460), .Q(regs_4
		[28]));
	notech_mux2 i_7238(.S(n_55986), .A(n_4395), .B(regs_4[28]), .Z(n_24751)
		);
	notech_reg regs_reg_4_29(.CP(n_63680), .D(n_24757), .CD(n_62460), .Q(regs_4
		[29]));
	notech_mux2 i_7246(.S(n_55986), .A(n_4394), .B(regs_4[29]), .Z(n_24757)
		);
	notech_reg regs_reg_4_30(.CP(n_63680), .D(n_24763), .CD(n_62460), .Q(regs_4
		[30]));
	notech_mux2 i_7256(.S(n_55986), .A(n_4361), .B(regs_4[30]), .Z(n_24763)
		);
	notech_reg regs_reg_4_31(.CP(n_63680), .D(n_24769), .CD(n_62460), .Q(regs_4
		[31]));
	notech_mux2 i_7264(.S(n_55986), .A(n_4423), .B(regs_4[31]), .Z(n_24769)
		);
	notech_reg regs_reg_3_0(.CP(n_63680), .D(n_24775), .CD(n_62460), .Q(regs_3
		[0]));
	notech_mux2 i_7272(.S(n_159362625), .A(n_31037), .B(regs_3[0]), .Z(n_24775
		));
	notech_reg regs_reg_3_1(.CP(n_63680), .D(n_24781), .CD(n_62460), .Q(regs_3
		[1]));
	notech_mux2 i_7280(.S(n_159362625), .A(n_31038), .B(regs_3[1]), .Z(n_24781
		));
	notech_reg regs_reg_3_2(.CP(n_63680), .D(n_24787), .CD(n_62460), .Q(regs_3
		[2]));
	notech_mux2 i_7288(.S(n_159362625), .A(n_440167985), .B(regs_3[2]), .Z(n_24787
		));
	notech_reg regs_reg_3_3(.CP(n_63680), .D(n_24793), .CD(n_62460), .Q(regs_3
		[3]));
	notech_mux2 i_7296(.S(n_159362625), .A(n_12662), .B(regs_3[3]), .Z(n_24793
		));
	notech_reg regs_reg_3_4(.CP(n_63680), .D(n_24799), .CD(n_62460), .Q(regs_3
		[4]));
	notech_mux2 i_7304(.S(n_159362625), .A(n_12668), .B(regs_3[4]), .Z(n_24799
		));
	notech_reg regs_reg_3_5(.CP(n_63680), .D(n_24805), .CD(n_62460), .Q(regs_3
		[5]));
	notech_mux2 i_7312(.S(n_159362625), .A(n_437382449), .B(regs_3[5]), .Z(n_24805
		));
	notech_reg regs_reg_3_6(.CP(n_63680), .D(n_24811), .CD(n_62464), .Q(regs_3
		[6]));
	notech_mux2 i_7320(.S(n_159362625), .A(n_12680), .B(regs_3[6]), .Z(n_24811
		));
	notech_reg regs_reg_3_7(.CP(n_63680), .D(n_24817), .CD(n_62464), .Q(regs_3
		[7]));
	notech_mux2 i_7328(.S(n_159362625), .A(n_4372), .B(regs_3[7]), .Z(n_24817
		));
	notech_reg regs_reg_3_8(.CP(n_63680), .D(n_24823), .CD(n_62464), .Q(regs_3
		[8]));
	notech_mux2 i_7336(.S(n_159362625), .A(n_31039), .B(regs_3[8]), .Z(n_24823
		));
	notech_reg regs_reg_3_9(.CP(n_63680), .D(n_24829), .CD(n_62464), .Q(regs_3
		[9]));
	notech_mux2 i_7344(.S(n_159362625), .A(n_4371), .B(regs_3[9]), .Z(n_24829
		));
	notech_reg regs_reg_3_10(.CP(n_63684), .D(n_24835), .CD(n_62464), .Q(regs_3
		[10]));
	notech_mux2 i_7352(.S(n_159362625), .A(n_384364374), .B(regs_3[10]), .Z(n_24835
		));
	notech_reg regs_reg_3_11(.CP(n_63640), .D(n_24841), .CD(n_62464), .Q(regs_3
		[11]));
	notech_mux2 i_7360(.S(n_159362625), .A(n_440067984), .B(regs_3[11]), .Z(n_24841
		));
	notech_reg regs_reg_3_12(.CP(n_63640), .D(n_24847), .CD(n_62464), .Q(regs_3
		[12]));
	notech_mux2 i_7368(.S(n_159362625), .A(n_439267976), .B(regs_3[12]), .Z(n_24847
		));
	notech_reg regs_reg_3_13(.CP(n_63640), .D(n_24853), .CD(n_62464), .Q(regs_3
		[13]));
	notech_mux2 i_7376(.S(n_159362625), .A(n_30657), .B(regs_3[13]), .Z(n_24853
		));
	notech_reg regs_reg_3_14(.CP(n_63640), .D(n_24861), .CD(n_62464), .Q(regs_3
		[14]));
	notech_mux2 i_7384(.S(n_159362625), .A(n_31040), .B(regs_3[14]), .Z(n_24861
		));
	notech_reg regs_reg_3_15(.CP(n_63640), .D(n_24869), .CD(n_62464), .Q(regs_3
		[15]));
	notech_mux2 i_7392(.S(n_159362625), .A(n_439167975), .B(regs_3[15]), .Z(n_24869
		));
	notech_reg regs_reg_3_16(.CP(n_63640), .D(n_24875), .CD(n_62463), .Q(regs_3
		[16]));
	notech_mux2 i_7400(.S(n_56008), .A(n_12740), .B(regs_3[16]), .Z(n_24875)
		);
	notech_reg regs_reg_3_17(.CP(n_63640), .D(n_24881), .CD(n_62463), .Q(regs_3
		[17]));
	notech_mux2 i_7408(.S(n_56008), .A(n_31041), .B(regs_3[17]), .Z(n_24881)
		);
	notech_nand3 i_28478(.A(n_63698), .B(n_63764), .C(opb[1]), .Z(n_30920)
		);
	notech_reg regs_reg_3_18(.CP(n_63640), .D(n_24887), .CD(n_62463), .Q(regs_3
		[18]));
	notech_mux2 i_7416(.S(n_56008), .A(n_31042), .B(regs_3[18]), .Z(n_24887)
		);
	notech_nand3 i_28479(.A(n_63698), .B(n_63764), .C(opa[1]), .Z(n_30919)
		);
	notech_reg regs_reg_3_19(.CP(n_63640), .D(n_24893), .CD(n_62463), .Q(regs_3
		[19]));
	notech_mux2 i_7424(.S(n_56008), .A(n_31043), .B(regs_3[19]), .Z(n_24893)
		);
	notech_nand2 i_28482(.A(n_63792), .B(opc_10[1]), .Z(n_30916));
	notech_reg regs_reg_3_20(.CP(n_63640), .D(n_24899), .CD(n_62463), .Q(regs_3
		[20]));
	notech_mux2 i_7432(.S(n_56008), .A(n_12764), .B(regs_3[20]), .Z(n_24899)
		);
	notech_nand2 i_28484(.A(n_63772), .B(opc[1]), .Z(n_30914));
	notech_reg regs_reg_3_21(.CP(n_63684), .D(n_24905), .CD(n_62464), .Q(regs_3
		[21]));
	notech_mux2 i_7440(.S(n_56008), .A(n_12770), .B(regs_3[21]), .Z(n_24905)
		);
	notech_nao3 i_28502(.A(n_63772), .B(opa[1]), .C(n_63712), .Z(n_30896));
	notech_reg regs_reg_3_22(.CP(n_63684), .D(n_24911), .CD(n_62464), .Q(regs_3
		[22]));
	notech_mux2 i_7448(.S(n_56008), .A(n_31044), .B(regs_3[22]), .Z(n_24911)
		);
	notech_reg regs_reg_3_23(.CP(n_63684), .D(n_24917), .CD(n_62463), .Q(regs_3
		[23]));
	notech_mux2 i_7456(.S(n_56008), .A(n_12782), .B(regs_3[23]), .Z(n_24917)
		);
	notech_reg regs_reg_3_24(.CP(n_63684), .D(n_24923), .CD(n_62463), .Q(regs_3
		[24]));
	notech_mux2 i_7464(.S(n_56008), .A(n_12788), .B(regs_3[24]), .Z(n_24923)
		);
	notech_ao4 i_140848379(.A(n_55955), .B(n_30973), .C(n_55975), .D(n_32062
		), .Z(n_2289));
	notech_reg regs_reg_3_25(.CP(n_63684), .D(n_24929), .CD(n_62419), .Q(regs_3
		[25]));
	notech_mux2 i_7472(.S(n_56008), .A(n_12794), .B(regs_3[25]), .Z(n_24929)
		);
	notech_ao4 i_140948378(.A(n_55966), .B(n_33117), .C(n_28240), .D(n_58256
		), .Z(n_2288));
	notech_reg regs_reg_3_26(.CP(n_63684), .D(n_24935), .CD(n_62373), .Q(regs_3
		[26]));
	notech_mux2 i_7480(.S(n_56008), .A(n_31045), .B(regs_3[26]), .Z(n_24935)
		);
	notech_and3 i_141448373(.A(n_2284), .B(n_2286), .C(n_2045), .Z(n_2287)
		);
	notech_reg regs_reg_3_27(.CP(n_63684), .D(n_24941), .CD(n_62373), .Q(regs_3
		[27]));
	notech_mux2 i_7488(.S(n_56008), .A(n_12806), .B(regs_3[27]), .Z(n_24941)
		);
	notech_ao4 i_141148376(.A(n_331160939), .B(\nbus_11290[3] ), .C(n_332260950
		), .D(n_33118), .Z(n_2286));
	notech_reg regs_reg_3_28(.CP(n_63684), .D(n_24947), .CD(n_62373), .Q(regs_3
		[28]));
	notech_mux2 i_7496(.S(n_56008), .A(n_31046), .B(regs_3[28]), .Z(n_24947)
		);
	notech_reg regs_reg_3_29(.CP(n_63684), .D(n_24953), .CD(n_62373), .Q(regs_3
		[29]));
	notech_mux2 i_7504(.S(n_56008), .A(n_31049), .B(regs_3[29]), .Z(n_24953)
		);
	notech_ao4 i_141248375(.A(n_331460942), .B(n_58784), .C(n_55946), .D(n_31511
		), .Z(n_2284));
	notech_reg regs_reg_3_30(.CP(n_63684), .D(n_24959), .CD(n_62374), .Q(regs_3
		[30]));
	notech_mux2 i_7512(.S(n_56008), .A(n_31050), .B(regs_3[30]), .Z(n_24959)
		);
	notech_and4 i_142448363(.A(n_2052), .B(n_2279), .C(n_2281), .D(n_2278), 
		.Z(n_2283));
	notech_reg regs_reg_3_31(.CP(n_63684), .D(n_24965), .CD(n_62374), .Q(regs_3
		[31]));
	notech_mux2 i_7520(.S(n_56008), .A(n_12830), .B(regs_3[31]), .Z(n_24965)
		);
	notech_reg_set cr0_reg_0(.CP(n_63684), .D(n_24971), .SD(n_62374), .Q(\nbus_14546[0] 
		));
	notech_mux2 i_7528(.S(n_97990346), .A(opa[0]), .B(n_61279), .Z(n_24971)
		);
	notech_ao4 i_141648371(.A(n_61094), .B(n_30779), .C(n_338161009), .D(n_26603
		), .Z(n_2281));
	notech_reg cr0_reg_1(.CP(n_63684), .D(n_24977), .CD(n_62374), .Q(\nbus_14542[1] 
		));
	notech_mux2 i_7536(.S(n_97990346), .A(opa[1]), .B(\nbus_14542[1] ), .Z(n_24977
		));
	notech_reg cr0_reg_2(.CP(n_63684), .D(n_24983), .CD(n_62374), .Q(cr0[2])
		);
	notech_mux2 i_7544(.S(n_97990346), .A(opa[2]), .B(cr0[2]), .Z(n_24983)
		);
	notech_ao4 i_141748370(.A(n_332160949), .B(n_74622849), .C(n_74822851), 
		.D(n_26278), .Z(n_2279));
	notech_reg cr0_reg_3(.CP(n_63684), .D(n_24989), .CD(n_62373), .Q(\nbus_14542[3] 
		));
	notech_mux2 i_7552(.S(n_97990346), .A(n_60971), .B(\nbus_14542[3] ), .Z(n_24989
		));
	notech_and3 i_142348364(.A(n_2275), .B(n_227795867), .C(n_2057), .Z(n_2278
		));
	notech_reg cr0_reg_4(.CP(n_63684), .D(n_24995), .CD(n_62373), .Q(\nbus_14542[4] 
		));
	notech_mux2 i_7560(.S(n_97990346), .A(opa[4]), .B(\nbus_14542[4] ), .Z(n_24995
		));
	notech_ao4 i_142048367(.A(n_75522858), .B(n_26277), .C(n_75622859), .D(n_26276
		), .Z(n_227795867));
	notech_reg cr0_reg_5(.CP(n_63684), .D(n_25001), .CD(n_62373), .Q(\nbus_14542[5] 
		));
	notech_mux2 i_7568(.S(n_97990346), .A(n_60980), .B(\nbus_14542[5] ), .Z(n_25001
		));
	notech_reg cr0_reg_6(.CP(n_63684), .D(n_25007), .CD(n_62370), .Q(\nbus_14542[6] 
		));
	notech_mux2 i_7576(.S(n_97990346), .A(opa[6]), .B(\nbus_14542[6] ), .Z(n_25007
		));
	notech_ao4 i_142148366(.A(n_75222855), .B(n_26272), .C(n_74922852), .D(n_26268
		), .Z(n_2275));
	notech_reg cr0_reg_7(.CP(n_63640), .D(n_25013), .CD(n_62370), .Q(\nbus_14542[7] 
		));
	notech_mux2 i_7584(.S(n_97990346), .A(opa[7]), .B(\nbus_14542[7] ), .Z(n_25013
		));
	notech_reg cr0_reg_8(.CP(n_63640), .D(n_25019), .CD(n_62373), .Q(\nbus_14542[8] 
		));
	notech_mux2 i_7592(.S(n_97990346), .A(opa[8]), .B(\nbus_14542[8] ), .Z(n_25019
		));
	notech_reg cr0_reg_9(.CP(n_63642), .D(n_25025), .CD(n_62373), .Q(\nbus_14542[9] 
		));
	notech_mux2 i_7600(.S(n_97990346), .A(opa[9]), .B(\nbus_14542[9] ), .Z(n_25025
		));
	notech_ao4 i_194247851(.A(n_57117), .B(n_31774), .C(n_57609), .D(n_33120
		), .Z(n_2272));
	notech_reg cr0_reg_10(.CP(n_63642), .D(n_25031), .CD(n_62373), .Q(\nbus_14542[10] 
		));
	notech_mux2 i_7608(.S(n_97990346), .A(opa[10]), .B(\nbus_14542[10] ), .Z
		(n_25031));
	notech_ao4 i_194347850(.A(n_57136), .B(n_31742), .C(n_57152), .D(n_33119
		), .Z(n_2271));
	notech_reg cr0_reg_11(.CP(n_63642), .D(n_25037), .CD(n_62373), .Q(\nbus_14542[11] 
		));
	notech_mux2 i_7616(.S(n_97990346), .A(opa[11]), .B(\nbus_14542[11] ), .Z
		(n_25037));
	notech_and2 i_194747846(.A(n_2269), .B(n_2268), .Z(n_2270));
	notech_reg cr0_reg_12(.CP(n_63642), .D(n_25043), .CD(n_62373), .Q(\nbus_14542[12] 
		));
	notech_mux2 i_7624(.S(n_97990346), .A(opa[12]), .B(\nbus_14542[12] ), .Z
		(n_25043));
	notech_ao4 i_194547848(.A(n_57163), .B(n_31838), .C(n_57178), .D(n_31999
		), .Z(n_2269));
	notech_reg cr0_reg_13(.CP(n_63642), .D(n_25049), .CD(n_62375), .Q(\nbus_14542[13] 
		));
	notech_mux2 i_7632(.S(n_97990346), .A(opa[13]), .B(\nbus_14542[13] ), .Z
		(n_25049));
	notech_ao4 i_194647847(.A(n_57189), .B(n_31710), .C(n_57199), .D(n_31934
		), .Z(n_2268));
	notech_reg cr0_reg_14(.CP(n_63642), .D(n_25055), .CD(n_62375), .Q(\nbus_14542[14] 
		));
	notech_mux2 i_7640(.S(n_97990346), .A(opa[14]), .B(\nbus_14542[14] ), .Z
		(n_25055));
	notech_and4 i_195547838(.A(n_2265), .B(n_2264), .C(n_2262), .D(n_2261), 
		.Z(n_2267));
	notech_reg cr0_reg_15(.CP(n_63642), .D(n_25061), .CD(n_62375), .Q(\nbus_14542[15] 
		));
	notech_mux2 i_7648(.S(n_97990346), .A(opa[15]), .B(\nbus_14542[15] ), .Z
		(n_25061));
	notech_reg cr0_reg_16(.CP(n_63642), .D(n_25067), .CD(n_62375), .Q(cr0[16
		]));
	notech_mux2 i_7656(.S(n_61596), .A(opa[16]), .B(cr0[16]), .Z(n_25067));
	notech_ao4 i_194947844(.A(n_57059), .B(n_31678), .C(n_57072), .D(n_31806
		), .Z(n_2265));
	notech_reg cr0_reg_17(.CP(n_63642), .D(n_25073), .CD(n_62375), .Q(\nbus_14542[17] 
		));
	notech_mux2 i_7664(.S(n_61596), .A(opa[17]), .B(\nbus_14542[17] ), .Z(n_25073
		));
	notech_ao4 i_195047843(.A(n_57086), .B(n_31870), .C(n_57097), .D(n_31575
		), .Z(n_2264));
	notech_reg cr0_reg_18(.CP(n_63642), .D(n_25079), .CD(n_62375), .Q(\nbus_14542[18] 
		));
	notech_mux2 i_7672(.S(n_61596), .A(opa[18]), .B(\nbus_14542[18] ), .Z(n_25079
		));
	notech_reg cr0_reg_19(.CP(n_63642), .D(n_25085), .CD(n_62375), .Q(\nbus_14542[19] 
		));
	notech_mux2 i_7680(.S(n_61596), .A(opa[19]), .B(\nbus_14542[19] ), .Z(n_25085
		));
	notech_ao4 i_195247841(.A(n_58696), .B(n_31967), .C(n_59095), .D(n_31902
		), .Z(n_2262));
	notech_reg cr0_reg_20(.CP(n_63642), .D(n_25092), .CD(n_62375), .Q(\nbus_14542[20] 
		));
	notech_mux2 i_7688(.S(n_61596), .A(opa[20]), .B(\nbus_14542[20] ), .Z(n_25092
		));
	notech_ao4 i_195347840(.A(n_57211), .B(n_31411), .C(n_57225), .D(n_31646
		), .Z(n_2261));
	notech_reg cr0_reg_21(.CP(n_63642), .D(n_25100), .CD(n_62375), .Q(\nbus_14542[21] 
		));
	notech_mux2 i_7696(.S(n_61596), .A(opa[21]), .B(\nbus_14542[21] ), .Z(n_25100
		));
	notech_nand2 i_10049744(.A(n_63772), .B(opc_10[3]), .Z(n_74522848));
	notech_reg cr0_reg_22(.CP(n_63642), .D(n_25106), .CD(n_62375), .Q(\nbus_14542[22] 
		));
	notech_mux2 i_7704(.S(n_61596), .A(opa[22]), .B(\nbus_14542[22] ), .Z(n_25106
		));
	notech_nao3 i_33649743(.A(n_61928), .B(opa[3]), .C(n_63712), .Z(n_74622849
		));
	notech_reg cr0_reg_23(.CP(n_63642), .D(n_25113), .CD(n_62374), .Q(\nbus_14542[23] 
		));
	notech_mux2 i_7712(.S(n_61596), .A(opa[23]), .B(\nbus_14542[23] ), .Z(n_25113
		));
	notech_nao3 i_34149742(.A(n_63772), .B(opa[3]), .C(n_63702), .Z(n_74822851
		));
	notech_reg cr0_reg_24(.CP(n_63642), .D(n_25119), .CD(n_62374), .Q(\nbus_14542[24] 
		));
	notech_mux2 i_7720(.S(n_61596), .A(opa[24]), .B(\nbus_14542[24] ), .Z(n_25119
		));
	notech_nand2 i_36149737(.A(n_63744), .B(opc[3]), .Z(n_74922852));
	notech_reg cr0_reg_25(.CP(n_63642), .D(n_25126), .CD(n_62374), .Q(\nbus_14542[25] 
		));
	notech_mux2 i_7728(.S(n_61596), .A(opa[25]), .B(\nbus_14542[25] ), .Z(n_25126
		));
	notech_nand3 i_35749738(.A(n_63698), .B(n_63764), .C(opa[3]), .Z(n_75222855
		));
	notech_reg cr0_reg_26(.CP(n_63642), .D(n_25132), .CD(n_62374), .Q(\nbus_14542[26] 
		));
	notech_mux2 i_7736(.S(n_61596), .A(opa[26]), .B(\nbus_14542[26] ), .Z(n_25132
		));
	notech_nand3 i_35649739(.A(n_63698), .B(n_61928), .C(opa[3]), .Z(n_75322856
		));
	notech_reg cr0_reg_27(.CP(n_63642), .D(n_25138), .CD(n_62374), .Q(\nbus_14542[27] 
		));
	notech_mux2 i_7744(.S(n_61596), .A(opa[27]), .B(\nbus_14542[27] ), .Z(n_25138
		));
	notech_nand3 i_35249741(.A(n_63720), .B(n_63764), .C(opb[3]), .Z(n_75522858
		));
	notech_reg cr0_reg_28(.CP(n_63568), .D(n_25144), .CD(n_62375), .Q(\nbus_14542[28] 
		));
	notech_mux2 i_7752(.S(n_61596), .A(opa[28]), .B(\nbus_14542[28] ), .Z(n_25144
		));
	notech_nand3 i_35349740(.A(n_63720), .B(n_61928), .C(opb[3]), .Z(n_75622859
		));
	notech_reg cr0_reg_29(.CP(n_63568), .D(n_25150), .CD(n_62375), .Q(\nbus_14542[29] 
		));
	notech_mux2 i_7760(.S(n_61596), .A(opa[29]), .B(\nbus_14542[29] ), .Z(n_25150
		));
	notech_reg cr0_reg_30(.CP(n_63568), .D(n_25156), .CD(n_62374), .Q(\nbus_14542[30] 
		));
	notech_mux2 i_7768(.S(n_61596), .A(opa[30]), .B(\nbus_14542[30] ), .Z(n_25156
		));
	notech_reg cr0_reg_31(.CP(n_63568), .D(n_25162), .CD(n_62374), .Q(\nbus_14542[31] 
		));
	notech_mux2 i_7776(.S(n_61596), .A(opa[31]), .B(\nbus_14542[31] ), .Z(n_25162
		));
	notech_ao4 i_214047653(.A(n_57117), .B(n_31778), .C(n_57609), .D(n_33122
		), .Z(n_2258));
	notech_reg mask8b_reg_0(.CP(n_63568), .D(n_25168), .CD(n_62368), .Q(mask8b
		[0]));
	notech_mux2 i_7784(.S(n_31070), .A(mask8b[0]), .B(n_31064), .Z(n_25168)
		);
	notech_ao4 i_214147652(.A(n_57136), .B(n_31746), .C(n_57152), .D(n_33121
		), .Z(n_225795868));
	notech_reg mask8b_reg_1(.CP(n_63568), .D(n_25174), .CD(n_62368), .Q(mask8b
		[1]));
	notech_mux2 i_7792(.S(n_31070), .A(mask8b[1]), .B(n_31065), .Z(n_25174)
		);
	notech_and2 i_214547648(.A(n_2255), .B(n_2254), .Z(n_225695869));
	notech_reg mask8b_reg_2(.CP(n_63568), .D(n_25180), .CD(n_62368), .Q(mask8b
		[2]));
	notech_mux2 i_7800(.S(n_31070), .A(mask8b[2]), .B(n_11287), .Z(n_25180)
		);
	notech_ao4 i_214347650(.A(n_57163), .B(n_31842), .C(n_57178), .D(n_32003
		), .Z(n_2255));
	notech_reg opb_reg_0(.CP(n_63568), .D(n_25186), .CD(n_62368), .Q(opb[0])
		);
	notech_mux2 i_7808(.S(n_208880594), .A(n_31073), .B(opb[0]), .Z(n_25186)
		);
	notech_ao4 i_214447649(.A(n_57189), .B(n_31714), .C(n_57199), .D(n_31938
		), .Z(n_2254));
	notech_reg opb_reg_1(.CP(n_63568), .D(n_25192), .CD(n_62368), .Q(opb[1])
		);
	notech_mux2 i_7816(.S(n_208880594), .A(n_31076), .B(opb[1]), .Z(n_25192)
		);
	notech_and4 i_215347640(.A(n_2251), .B(n_2250), .C(n_2248), .D(n_2247), 
		.Z(n_2253));
	notech_reg opb_reg_2(.CP(n_63568), .D(n_25198), .CD(n_62369), .Q(opb[2])
		);
	notech_mux2 i_7824(.S(n_208880594), .A(n_31077), .B(opb[2]), .Z(n_25198)
		);
	notech_reg opb_reg_3(.CP(n_63568), .D(n_25204), .CD(n_62369), .Q(opb[3])
		);
	notech_mux2 i_7832(.S(n_208880594), .A(n_4431), .B(opb[3]), .Z(n_25204)
		);
	notech_ao4 i_214747646(.A(n_57059), .B(n_31682), .C(n_57072), .D(n_31810
		), .Z(n_2251));
	notech_reg opb_reg_4(.CP(n_63568), .D(n_25210), .CD(n_62368), .Q(opb[4])
		);
	notech_mux2 i_7840(.S(n_208880594), .A(n_13641), .B(opb[4]), .Z(n_25210)
		);
	notech_ao4 i_214847645(.A(n_57086), .B(n_31874), .C(n_57097), .D(n_31579
		), .Z(n_2250));
	notech_reg opb_reg_5(.CP(n_63650), .D(n_25216), .CD(n_62369), .Q(opb[5])
		);
	notech_mux2 i_7848(.S(n_208880594), .A(n_13647), .B(opb[5]), .Z(n_25216)
		);
	notech_reg opb_reg_6(.CP(n_63500), .D(n_25222), .CD(n_62368), .Q(opb[6])
		);
	notech_mux2 i_7856(.S(n_208880594), .A(n_13653), .B(opb[6]), .Z(n_25222)
		);
	notech_ao4 i_215047643(.A(n_58696), .B(n_31971), .C(n_59099), .D(n_31906
		), .Z(n_2248));
	notech_reg opb_reg_7(.CP(n_63500), .D(n_25228), .CD(n_62367), .Q(opb[7])
		);
	notech_mux2 i_7865(.S(n_208880594), .A(n_13659), .B(opb[7]), .Z(n_25228)
		);
	notech_ao4 i_215147642(.A(n_57211), .B(n_31415), .C(n_57225), .D(n_31650
		), .Z(n_2247));
	notech_reg opb_reg_8(.CP(n_63500), .D(n_25234), .CD(n_62367), .Q(opb[8])
		);
	notech_mux2 i_7873(.S(n_208880594), .A(n_31078), .B(opb[8]), .Z(n_25234)
		);
	notech_reg opb_reg_9(.CP(n_63500), .D(n_25240), .CD(n_62367), .Q(opb[9])
		);
	notech_mux2 i_7881(.S(n_208880594), .A(n_31079), .B(opb[9]), .Z(n_25240)
		);
	notech_reg opb_reg_10(.CP(n_63500), .D(n_25246), .CD(n_62367), .Q(opb[10
		]));
	notech_mux2 i_7889(.S(n_208880594), .A(n_30637), .B(opb[10]), .Z(n_25246
		));
	notech_ao4 i_215447639(.A(n_57117), .B(n_31777), .C(n_57604), .D(n_33124
		), .Z(n_2244));
	notech_reg opb_reg_11(.CP(n_63500), .D(n_25252), .CD(n_62368), .Q(opb[11
		]));
	notech_mux2 i_7897(.S(n_208880594), .A(n_30419), .B(opb[11]), .Z(n_25252
		));
	notech_ao4 i_215547638(.A(n_57130), .B(n_31745), .C(n_57152), .D(n_33123
		), .Z(n_2243));
	notech_reg opb_reg_12(.CP(n_63500), .D(n_25258), .CD(n_62368), .Q(opb[12
		]));
	notech_mux2 i_7905(.S(n_208880594), .A(n_30423), .B(opb[12]), .Z(n_25258
		));
	notech_and2 i_215947634(.A(n_2241), .B(n_2240), .Z(n_2242));
	notech_reg opb_reg_13(.CP(n_63500), .D(n_25264), .CD(n_62368), .Q(opb[13
		]));
	notech_mux2 i_7913(.S(n_208880594), .A(n_30413), .B(opb[13]), .Z(n_25264
		));
	notech_ao4 i_215747636(.A(n_57163), .B(n_31841), .C(n_57178), .D(n_32002
		), .Z(n_2241));
	notech_reg opb_reg_14(.CP(n_63500), .D(n_25270), .CD(n_62368), .Q(opb[14
		]));
	notech_mux2 i_7921(.S(n_208880594), .A(n_31080), .B(opb[14]), .Z(n_25270
		));
	notech_ao4 i_215847635(.A(n_57189), .B(n_31713), .C(n_57199), .D(n_31937
		), .Z(n_2240));
	notech_reg opb_reg_15(.CP(n_63500), .D(n_25276), .CD(n_62368), .Q(opb[15
		]));
	notech_mux2 i_7929(.S(n_208880594), .A(n_446668050), .B(opb[15]), .Z(n_25276
		));
	notech_and4 i_216747626(.A(n_223795870), .B(n_223695871), .C(n_223495873
		), .D(n_223395874), .Z(n_2239));
	notech_reg opb_reg_16(.CP(n_63580), .D(n_25282), .CD(n_62370), .Q(opb[16
		]));
	notech_mux2 i_7937(.S(n_331981796), .A(n_13713), .B(opb[16]), .Z(n_25282
		));
	notech_reg opb_reg_17(.CP(n_63580), .D(n_25288), .CD(n_62370), .Q(opb[17
		]));
	notech_mux2 i_7945(.S(n_331981796), .A(n_31081), .B(opb[17]), .Z(n_25288
		));
	notech_ao4 i_216147632(.A(n_57059), .B(n_31681), .C(n_57072), .D(n_31809
		), .Z(n_223795870));
	notech_reg opb_reg_18(.CP(n_63580), .D(n_25294), .CD(n_62370), .Q(opb[18
		]));
	notech_mux2 i_7953(.S(n_331981796), .A(n_31082), .B(opb[18]), .Z(n_25294
		));
	notech_ao4 i_216247631(.A(n_57086), .B(n_31873), .C(n_57103), .D(n_31578
		), .Z(n_223695871));
	notech_reg opb_reg_19(.CP(n_63580), .D(n_25300), .CD(n_62370), .Q(opb[19
		]));
	notech_mux2 i_7961(.S(n_331981796), .A(n_13731), .B(opb[19]), .Z(n_25300
		));
	notech_reg opb_reg_20(.CP(n_63580), .D(n_25306), .CD(n_62370), .Q(opb[20
		]));
	notech_mux2 i_7969(.S(n_331981796), .A(n_13737), .B(opb[20]), .Z(n_25306
		));
	notech_ao4 i_216447629(.A(n_58696), .B(n_31970), .C(n_59099), .D(n_31905
		), .Z(n_223495873));
	notech_reg opb_reg_21(.CP(n_63580), .D(n_25312), .CD(n_62370), .Q(opb[21
		]));
	notech_mux2 i_7977(.S(n_331981796), .A(n_13743), .B(opb[21]), .Z(n_25312
		));
	notech_ao4 i_216547628(.A(n_57211), .B(n_31414), .C(n_57225), .D(n_31649
		), .Z(n_223395874));
	notech_reg opb_reg_22(.CP(n_63580), .D(n_25318), .CD(n_62370), .Q(opb[22
		]));
	notech_mux2 i_7985(.S(n_331981796), .A(n_13749), .B(opb[22]), .Z(n_25318
		));
	notech_reg opb_reg_23(.CP(n_63580), .D(n_25324), .CD(n_62370), .Q(opb[23
		]));
	notech_mux2 i_7993(.S(n_331981796), .A(n_13755), .B(opb[23]), .Z(n_25324
		));
	notech_reg opb_reg_24(.CP(n_63580), .D(n_25330), .CD(n_62370), .Q(opb[24
		]));
	notech_mux2 i_8001(.S(n_331981796), .A(n_13761), .B(opb[24]), .Z(n_25330
		));
	notech_ao4 i_216847625(.A(n_57117), .B(n_31776), .C(n_57604), .D(n_33126
		), .Z(n_2230));
	notech_reg opb_reg_25(.CP(n_63580), .D(n_25336), .CD(n_62370), .Q(opb[25
		]));
	notech_mux2 i_8009(.S(n_331981796), .A(n_13767), .B(opb[25]), .Z(n_25336
		));
	notech_ao4 i_216947624(.A(n_57130), .B(n_31744), .C(n_57152), .D(n_33125
		), .Z(n_2229));
	notech_reg opb_reg_26(.CP(n_63580), .D(n_25342), .CD(n_62369), .Q(opb[26
		]));
	notech_mux2 i_8017(.S(n_331981796), .A(n_13773), .B(opb[26]), .Z(n_25342
		));
	notech_and2 i_217347620(.A(n_2227), .B(n_2226), .Z(n_2228));
	notech_reg opb_reg_27(.CP(n_63580), .D(n_25348), .CD(n_62369), .Q(opb[27
		]));
	notech_mux2 i_8025(.S(n_331981796), .A(n_13779), .B(opb[27]), .Z(n_25348
		));
	notech_ao4 i_217147622(.A(n_57163), .B(n_31840), .C(n_57174), .D(n_32001
		), .Z(n_2227));
	notech_reg opb_reg_28(.CP(n_63580), .D(n_25354), .CD(n_62369), .Q(opb[28
		]));
	notech_mux2 i_8033(.S(n_331981796), .A(n_13785), .B(opb[28]), .Z(n_25354
		));
	notech_ao4 i_217247621(.A(n_57189), .B(n_31712), .C(n_57199), .D(n_31936
		), .Z(n_2226));
	notech_reg opb_reg_29(.CP(n_63580), .D(n_25360), .CD(n_62369), .Q(opb[29
		]));
	notech_mux2 i_8041(.S(n_331981796), .A(n_4429), .B(opb[29]), .Z(n_25360)
		);
	notech_and4 i_218147612(.A(n_2223), .B(n_2222), .C(n_2220), .D(n_2219), 
		.Z(n_2225));
	notech_reg opb_reg_30(.CP(n_63580), .D(n_25366), .CD(n_62369), .Q(opb[30
		]));
	notech_mux2 i_8049(.S(n_331981796), .A(n_13797), .B(opb[30]), .Z(n_25366
		));
	notech_reg opb_reg_31(.CP(n_63580), .D(n_25372), .CD(n_62369), .Q(opb[31
		]));
	notech_mux2 i_8057(.S(n_331981796), .A(n_13803), .B(n_60629), .Z(n_25372
		));
	notech_ao4 i_217547618(.A(n_57059), .B(n_31680), .C(n_57068), .D(n_31808
		), .Z(n_2223));
	notech_reg regs_reg_2_0(.CP(n_63580), .D(n_25378), .CD(n_62369), .Q(regs_2
		[0]));
	notech_mux2 i_8065(.S(\nbus_11305[0] ), .A(regs_2[0]), .B(n_12292), .Z(n_25378
		));
	notech_ao4 i_217647617(.A(n_57086), .B(n_31872), .C(n_57097), .D(n_31577
		), .Z(n_2222));
	notech_reg regs_reg_2_1(.CP(n_63580), .D(n_25384), .CD(n_62369), .Q(regs_2
		[1]));
	notech_mux2 i_8073(.S(\nbus_11305[0] ), .A(regs_2[1]), .B(n_12298), .Z(n_25384
		));
	notech_reg regs_reg_2_2(.CP(n_63580), .D(n_25390), .CD(n_62369), .Q(regs_2
		[2]));
	notech_mux2 i_8081(.S(\nbus_11305[0] ), .A(regs_2[2]), .B(n_441067994), 
		.Z(n_25390));
	notech_ao4 i_217847615(.A(n_58696), .B(n_31969), .C(n_59099), .D(n_31904
		), .Z(n_2220));
	notech_reg regs_reg_2_3(.CP(n_63578), .D(n_25396), .CD(n_62381), .Q(regs_2
		[3]));
	notech_mux2 i_8089(.S(\nbus_11305[0] ), .A(regs_2[3]), .B(n_31083), .Z(n_25396
		));
	notech_ao4 i_217947614(.A(n_57211), .B(n_31413), .C(n_57225), .D(n_31648
		), .Z(n_2219));
	notech_reg regs_reg_2_4(.CP(n_63578), .D(n_25402), .CD(n_62381), .Q(regs_2
		[4]));
	notech_mux2 i_8097(.S(\nbus_11305[0] ), .A(regs_2[4]), .B(n_31084), .Z(n_25402
		));
	notech_reg regs_reg_2_5(.CP(n_63654), .D(n_25408), .CD(n_62381), .Q(regs_2
		[5]));
	notech_mux2 i_8105(.S(\nbus_11305[0] ), .A(regs_2[5]), .B(n_30398), .Z(n_25408
		));
	notech_reg regs_reg_2_6(.CP(n_63654), .D(n_25414), .CD(n_62381), .Q(regs_2
		[6]));
	notech_mux2 i_8113(.S(\nbus_11305[0] ), .A(regs_2[6]), .B(n_31085), .Z(n_25414
		));
	notech_ao4 i_218247611(.A(n_57117), .B(n_31775), .C(n_57604), .D(n_33128
		), .Z(n_2216));
	notech_reg regs_reg_2_7(.CP(n_63654), .D(n_25420), .CD(n_62381), .Q(regs_2
		[7]));
	notech_mux2 i_8121(.S(\nbus_11305[0] ), .A(regs_2[7]), .B(n_4381), .Z(n_25420
		));
	notech_ao4 i_218347610(.A(n_57130), .B(n_31743), .C(n_57152), .D(n_33127
		), .Z(n_2215));
	notech_reg regs_reg_2_8(.CP(n_63654), .D(n_25426), .CD(n_62381), .Q(regs_2
		[8]));
	notech_mux2 i_8129(.S(\nbus_11305[0] ), .A(regs_2[8]), .B(n_12340), .Z(n_25426
		));
	notech_and2 i_218747606(.A(n_2213), .B(n_2212), .Z(n_2214));
	notech_reg regs_reg_2_9(.CP(n_63654), .D(n_25434), .CD(n_62381), .Q(regs_2
		[9]));
	notech_mux2 i_8137(.S(\nbus_11305[0] ), .A(regs_2[9]), .B(n_30397), .Z(n_25434
		));
	notech_ao4 i_218547608(.A(n_57163), .B(n_31839), .C(n_57174), .D(n_32000
		), .Z(n_2213));
	notech_reg regs_reg_2_10(.CP(n_63654), .D(n_25440), .CD(n_62381), .Q(regs_2
		[10]));
	notech_mux2 i_8145(.S(\nbus_11305[0] ), .A(regs_2[10]), .B(n_30644), .Z(n_25440
		));
	notech_ao4 i_218647607(.A(n_57189), .B(n_31711), .C(n_57199), .D(n_31935
		), .Z(n_2212));
	notech_reg regs_reg_2_11(.CP(n_63654), .D(n_25446), .CD(n_62381), .Q(regs_2
		[11]));
	notech_mux2 i_8153(.S(\nbus_11305[0] ), .A(regs_2[11]), .B(n_30437), .Z(n_25446
		));
	notech_and4 i_219547598(.A(n_2209), .B(n_2208), .C(n_2206), .D(n_2205), 
		.Z(n_2211));
	notech_reg regs_reg_2_12(.CP(n_63654), .D(n_25452), .CD(n_62380), .Q(regs_2
		[12]));
	notech_mux2 i_8161(.S(\nbus_11305[0] ), .A(regs_2[12]), .B(n_440867992),
		 .Z(n_25452));
	notech_reg regs_reg_2_13(.CP(n_63654), .D(n_25458), .CD(n_62380), .Q(regs_2
		[13]));
	notech_mux2 i_8169(.S(\nbus_11305[0] ), .A(regs_2[13]), .B(n_30645), .Z(n_25458
		));
	notech_ao4 i_218947604(.A(n_57059), .B(n_31679), .C(n_57068), .D(n_31807
		), .Z(n_2209));
	notech_reg regs_reg_2_14(.CP(n_63654), .D(n_25464), .CD(n_62380), .Q(regs_2
		[14]));
	notech_mux2 i_8177(.S(\nbus_11305[0] ), .A(regs_2[14]), .B(n_31086), .Z(n_25464
		));
	notech_ao4 i_219047603(.A(n_57081), .B(n_31871), .C(n_57097), .D(n_31576
		), .Z(n_2208));
	notech_reg regs_reg_2_15(.CP(n_63654), .D(n_25472), .CD(n_62380), .Q(regs_2
		[15]));
	notech_mux2 i_8185(.S(\nbus_11305[0] ), .A(regs_2[15]), .B(n_30438), .Z(n_25472
		));
	notech_reg regs_reg_2_16(.CP(n_63654), .D(n_25478), .CD(n_62380), .Q(regs_2
		[16]));
	notech_mux2 i_8193(.S(n_56019), .A(regs_2[16]), .B(n_12388), .Z(n_25478)
		);
	notech_ao4 i_219247601(.A(n_58696), .B(n_31968), .C(n_59099), .D(n_31903
		), .Z(n_2206));
	notech_reg regs_reg_2_17(.CP(n_63654), .D(n_25486), .CD(n_62380), .Q(regs_2
		[17]));
	notech_mux2 i_8201(.S(n_56019), .A(regs_2[17]), .B(n_31087), .Z(n_25486)
		);
	notech_ao4 i_219347600(.A(n_57211), .B(n_31412), .C(n_57225), .D(n_31647
		), .Z(n_2205));
	notech_reg regs_reg_2_18(.CP(n_63654), .D(n_25492), .CD(n_62380), .Q(regs_2
		[18]));
	notech_mux2 i_8209(.S(n_56019), .A(regs_2[18]), .B(n_12400), .Z(n_25492)
		);
	notech_nand2 i_112766178(.A(n_83739557), .B(n_83839558), .Z(n_220495876)
		);
	notech_reg regs_reg_2_19(.CP(n_63654), .D(n_25498), .CD(n_62380), .Q(regs_2
		[19]));
	notech_mux2 i_8217(.S(n_56019), .A(regs_2[19]), .B(n_31088), .Z(n_25498)
		);
	notech_reg regs_reg_2_20(.CP(n_63654), .D(n_25504), .CD(n_62380), .Q(regs_2
		[20]));
	notech_mux2 i_8225(.S(n_56019), .A(regs_2[20]), .B(n_3032), .Z(n_25504)
		);
	notech_reg regs_reg_2_21(.CP(n_63654), .D(n_25510), .CD(n_62380), .Q(regs_2
		[21]));
	notech_mux2 i_8233(.S(n_56019), .A(regs_2[21]), .B(n_12418), .Z(n_25510)
		);
	notech_reg regs_reg_2_22(.CP(n_63654), .D(n_25516), .CD(n_62384), .Q(regs_2
		[22]));
	notech_mux2 i_8241(.S(n_56019), .A(regs_2[22]), .B(n_338681853), .Z(n_25516
		));
	notech_reg regs_reg_2_23(.CP(n_63578), .D(n_25522), .CD(n_62384), .Q(regs_2
		[23]));
	notech_mux2 i_8249(.S(n_56019), .A(regs_2[23]), .B(n_12430), .Z(n_25522)
		);
	notech_reg regs_reg_2_24(.CP(n_63578), .D(n_25528), .CD(n_62384), .Q(regs_2
		[24]));
	notech_mux2 i_8257(.S(n_56019), .A(regs_2[24]), .B(n_337681843), .Z(n_25528
		));
	notech_reg regs_reg_2_25(.CP(n_63578), .D(n_25534), .CD(n_62384), .Q(regs_2
		[25]));
	notech_mux2 i_8265(.S(n_56019), .A(regs_2[25]), .B(n_336681833), .Z(n_25534
		));
	notech_reg regs_reg_2_26(.CP(n_63578), .D(n_25540), .CD(n_62384), .Q(regs_2
		[26]));
	notech_mux2 i_8273(.S(n_56019), .A(regs_2[26]), .B(n_31089), .Z(n_25540)
		);
	notech_reg regs_reg_2_27(.CP(n_63578), .D(n_25546), .CD(n_62385), .Q(regs_2
		[27]));
	notech_mux2 i_8281(.S(n_56019), .A(regs_2[27]), .B(n_12454), .Z(n_25546)
		);
	notech_reg regs_reg_2_28(.CP(n_63578), .D(n_25552), .CD(n_62385), .Q(regs_2
		[28]));
	notech_mux2 i_8289(.S(n_56019), .A(regs_2[28]), .B(n_31090), .Z(n_25552)
		);
	notech_reg regs_reg_2_29(.CP(n_63578), .D(n_25558), .CD(n_62385), .Q(regs_2
		[29]));
	notech_mux2 i_8297(.S(n_56019), .A(regs_2[29]), .B(n_30406), .Z(n_25558)
		);
	notech_reg regs_reg_2_30(.CP(n_63578), .D(n_25564), .CD(n_62385), .Q(regs_2
		[30]));
	notech_mux2 i_8305(.S(n_56019), .A(regs_2[30]), .B(n_12472), .Z(n_25564)
		);
	notech_reg regs_reg_2_31(.CP(n_63578), .D(n_25570), .CD(n_62384), .Q(regs_2
		[31]));
	notech_mux2 i_8313(.S(n_56019), .A(regs_2[31]), .B(n_31091), .Z(n_25570)
		);
	notech_ao4 i_225747536(.A(n_57112), .B(n_31773), .C(n_57609), .D(n_33130
		), .Z(n_2191));
	notech_reg regs_reg_1_0(.CP(n_63578), .D(n_25576), .CD(n_62381), .Q(ecx[
		0]));
	notech_mux2 i_8321(.S(\nbus_11304[0] ), .A(ecx[0]), .B(n_11935), .Z(n_25576
		));
	notech_ao4 i_225847535(.A(n_57130), .B(n_31741), .C(n_57152), .D(n_33129
		), .Z(n_2190));
	notech_reg regs_reg_1_1(.CP(n_63654), .D(n_25582), .CD(n_62384), .Q(ecx[
		1]));
	notech_mux2 i_8329(.S(\nbus_11304[0] ), .A(ecx[1]), .B(n_31092), .Z(n_25582
		));
	notech_and2 i_226247531(.A(n_2188), .B(n_2187), .Z(n_2189));
	notech_reg regs_reg_1_2(.CP(n_63500), .D(n_25588), .CD(n_62381), .Q(ecx[
		2]));
	notech_mux2 i_8337(.S(\nbus_11304[0] ), .A(ecx[2]), .B(n_30439), .Z(n_25588
		));
	notech_ao4 i_226047533(.A(n_57163), .B(n_31837), .C(n_57174), .D(n_31998
		), .Z(n_2188));
	notech_reg regs_reg_1_3(.CP(n_63576), .D(n_25594), .CD(n_62381), .Q(ecx[
		3]));
	notech_mux2 i_8345(.S(\nbus_11304[0] ), .A(ecx[3]), .B(n_31093), .Z(n_25594
		));
	notech_ao4 i_226147532(.A(n_57189), .B(n_31709), .C(n_57199), .D(n_31933
		), .Z(n_2187));
	notech_reg regs_reg_1_4(.CP(n_63650), .D(n_25600), .CD(n_62384), .Q(ecx[
		4]));
	notech_mux2 i_8353(.S(\nbus_11304[0] ), .A(ecx[4]), .B(n_30908), .Z(n_25600
		));
	notech_and4 i_227047523(.A(n_2184), .B(n_2183), .C(n_2179), .D(n_217860435
		), .Z(n_2186));
	notech_reg regs_reg_1_5(.CP(n_63650), .D(n_25606), .CD(n_62384), .Q(ecx[
		5]));
	notech_mux2 i_8361(.S(\nbus_11304[0] ), .A(ecx[5]), .B(n_30909), .Z(n_25606
		));
	notech_reg regs_reg_1_6(.CP(n_63650), .D(n_25612), .CD(n_62384), .Q(ecx[
		6]));
	notech_mux2 i_8369(.S(\nbus_11304[0] ), .A(ecx[6]), .B(n_31094), .Z(n_25612
		));
	notech_ao4 i_226447529(.A(n_57059), .B(n_31677), .C(n_57068), .D(n_31805
		), .Z(n_2184));
	notech_reg regs_reg_1_7(.CP(n_63650), .D(n_25618), .CD(n_62384), .Q(ecx[
		7]));
	notech_mux2 i_8377(.S(\nbus_11304[0] ), .A(ecx[7]), .B(n_30656), .Z(n_25618
		));
	notech_ao4 i_226547528(.A(n_57081), .B(n_31869), .C(n_57097), .D(n_31574
		), .Z(n_2183));
	notech_reg regs_reg_1_8(.CP(n_63650), .D(n_25624), .CD(n_62384), .Q(ecx[
		8]));
	notech_mux2 i_8385(.S(\nbus_11304[0] ), .A(ecx[8]), .B(n_11983), .Z(n_25624
		));
	notech_reg regs_reg_1_9(.CP(n_63650), .D(n_25630), .CD(n_62378), .Q(ecx[
		9]));
	notech_mux2 i_8393(.S(\nbus_11304[0] ), .A(ecx[9]), .B(n_4374), .Z(n_25630
		));
	notech_ao4 i_226747526(.A(n_58696), .B(n_31966), .C(n_59099), .D(n_31901
		), .Z(n_2179));
	notech_reg regs_reg_1_10(.CP(n_63650), .D(n_25636), .CD(n_62378), .Q(ecx
		[10]));
	notech_mux2 i_8401(.S(\nbus_11304[0] ), .A(ecx[10]), .B(n_380564336), .Z
		(n_25636));
	notech_ao4 i_226847525(.A(n_57211), .B(n_31410), .C(n_57225), .D(n_31645
		), .Z(n_217860435));
	notech_reg regs_reg_1_11(.CP(n_63650), .D(n_25642), .CD(n_62376), .Q(ecx
		[11]));
	notech_mux2 i_8409(.S(\nbus_11304[0] ), .A(ecx[11]), .B(n_440367987), .Z
		(n_25642));
	notech_reg regs_reg_1_12(.CP(n_63650), .D(n_25648), .CD(n_62376), .Q(ecx
		[12]));
	notech_mux2 i_8417(.S(\nbus_11304[0] ), .A(ecx[12]), .B(n_440267986), .Z
		(n_25648));
	notech_reg regs_reg_1_13(.CP(n_63650), .D(n_25655), .CD(n_62378), .Q(ecx
		[13]));
	notech_mux2 i_8425(.S(\nbus_11304[0] ), .A(ecx[13]), .B(n_380464335), .Z
		(n_25655));
	notech_reg regs_reg_1_14(.CP(n_63650), .D(n_25662), .CD(n_62378), .Q(ecx
		[14]));
	notech_mux2 i_8434(.S(\nbus_11304[0] ), .A(ecx[14]), .B(n_31095), .Z(n_25662
		));
	notech_reg regs_reg_1_15(.CP(n_63688), .D(n_25669), .CD(n_62378), .Q(ecx
		[15]));
	notech_mux2 i_8443(.S(\nbus_11304[0] ), .A(ecx[15]), .B(n_441167995), .Z
		(n_25669));
	notech_reg regs_reg_1_16(.CP(n_63688), .D(n_25677), .CD(n_62378), .Q(ecx
		[16]));
	notech_mux2 i_8452(.S(\nbus_11304[16] ), .A(ecx[16]), .B(n_12031), .Z(n_25677
		));
	notech_reg regs_reg_1_17(.CP(n_63688), .D(n_25686), .CD(n_62378), .Q(ecx
		[17]));
	notech_mux2 i_8460(.S(\nbus_11304[16] ), .A(ecx[17]), .B(n_31096), .Z(n_25686
		));
	notech_reg regs_reg_1_18(.CP(n_63688), .D(n_25693), .CD(n_62376), .Q(ecx
		[18]));
	notech_mux2 i_8468(.S(\nbus_11304[16] ), .A(ecx[18]), .B(n_12043), .Z(n_25693
		));
	notech_reg regs_reg_1_19(.CP(n_63688), .D(n_25700), .CD(n_62376), .Q(ecx
		[19]));
	notech_mux2 i_8476(.S(\nbus_11304[16] ), .A(ecx[19]), .B(n_31097), .Z(n_25700
		));
	notech_reg regs_reg_1_20(.CP(n_63688), .D(n_25707), .CD(n_62376), .Q(ecx
		[20]));
	notech_mux2 i_8484(.S(\nbus_11304[16] ), .A(ecx[20]), .B(n_12055), .Z(n_25707
		));
	notech_reg regs_reg_1_21(.CP(n_63688), .D(n_25714), .CD(n_62376), .Q(ecx
		[21]));
	notech_mux2 i_8492(.S(\nbus_11304[16] ), .A(ecx[21]), .B(n_12061), .Z(n_25714
		));
	notech_reg regs_reg_1_22(.CP(n_63688), .D(n_25720), .CD(n_62376), .Q(ecx
		[22]));
	notech_mux2 i_8500(.S(\nbus_11304[16] ), .A(ecx[22]), .B(n_12067), .Z(n_25720
		));
	notech_reg regs_reg_1_23(.CP(n_63688), .D(n_25726), .CD(n_62376), .Q(ecx
		[23]));
	notech_mux2 i_8508(.S(\nbus_11304[16] ), .A(ecx[23]), .B(n_12073), .Z(n_25726
		));
	notech_reg regs_reg_1_24(.CP(n_63688), .D(n_25732), .CD(n_62376), .Q(ecx
		[24]));
	notech_mux2 i_8516(.S(\nbus_11304[16] ), .A(ecx[24]), .B(n_12079), .Z(n_25732
		));
	notech_reg regs_reg_1_25(.CP(n_63688), .D(n_25738), .CD(n_62376), .Q(ecx
		[25]));
	notech_mux2 i_8525(.S(\nbus_11304[16] ), .A(ecx[25]), .B(n_12085), .Z(n_25738
		));
	notech_reg regs_reg_1_26(.CP(n_63688), .D(n_25744), .CD(n_62376), .Q(ecx
		[26]));
	notech_mux2 i_8533(.S(\nbus_11304[16] ), .A(ecx[26]), .B(n_12091), .Z(n_25744
		));
	notech_reg regs_reg_1_27(.CP(n_63688), .D(n_25751), .CD(n_62376), .Q(ecx
		[27]));
	notech_mux2 i_8541(.S(\nbus_11304[16] ), .A(ecx[27]), .B(n_12097), .Z(n_25751
		));
	notech_reg regs_reg_1_28(.CP(n_63688), .D(n_25757), .CD(n_62379), .Q(ecx
		[28]));
	notech_mux2 i_8549(.S(\nbus_11304[16] ), .A(ecx[28]), .B(n_31100), .Z(n_25757
		));
	notech_nand2 i_32027(.A(n_63748), .B(n_27378), .Z(n_27371));
	notech_reg regs_reg_1_29(.CP(n_63688), .D(n_25763), .CD(n_62379), .Q(ecx
		[29]));
	notech_mux2 i_8557(.S(\nbus_11304[16] ), .A(ecx[29]), .B(n_12109), .Z(n_25763
		));
	notech_reg regs_reg_1_30(.CP(n_63688), .D(n_25769), .CD(n_62379), .Q(ecx
		[30]));
	notech_mux2 i_8565(.S(\nbus_11304[16] ), .A(ecx[30]), .B(n_12115), .Z(n_25769
		));
	notech_reg regs_reg_1_31(.CP(n_63688), .D(n_25775), .CD(n_62379), .Q(ecx
		[31]));
	notech_mux2 i_8573(.S(\nbus_11304[16] ), .A(ecx[31]), .B(n_31101), .Z(n_25775
		));
	notech_reg_set divq_reg_0(.CP(n_63688), .D(n_25781), .SD(1'b1), .Q(divq[
		0]));
	notech_mux2 i_8581(.S(n_56397), .A(divq[0]), .B(n_7784), .Z(n_25781));
	notech_reg_set divq_reg_1(.CP(n_63650), .D(n_25787), .SD(1'b1), .Q(divq[
		1]));
	notech_mux2 i_8589(.S(n_56397), .A(divq[1]), .B(n_7789), .Z(n_25787));
	notech_reg_set divq_reg_2(.CP(n_63688), .D(n_25793), .SD(1'b1), .Q(divq[
		2]));
	notech_mux2 i_8597(.S(n_56397), .A(divq[2]), .B(n_7794), .Z(n_25793));
	notech_reg_set divq_reg_3(.CP(n_63652), .D(n_25799), .SD(1'b1), .Q(divq[
		3]));
	notech_mux2 i_8605(.S(n_56397), .A(divq[3]), .B(n_7799), .Z(n_25799));
	notech_reg_set divq_reg_4(.CP(n_63652), .D(n_25805), .SD(1'b1), .Q(divq[
		4]));
	notech_mux2 i_8613(.S(n_56397), .A(divq[4]), .B(n_7804), .Z(n_25805));
	notech_reg_set divq_reg_5(.CP(n_63652), .D(n_25811), .SD(1'b1), .Q(divq[
		5]));
	notech_mux2 i_8621(.S(n_56397), .A(divq[5]), .B(n_7809), .Z(n_25811));
	notech_reg_set divq_reg_6(.CP(n_63652), .D(n_25817), .SD(1'b1), .Q(divq[
		6]));
	notech_mux2 i_8629(.S(n_56397), .A(divq[6]), .B(n_7814), .Z(n_25817));
	notech_reg_set divq_reg_7(.CP(n_63652), .D(n_25823), .SD(1'b1), .Q(divq[
		7]));
	notech_mux2 i_8637(.S(n_56397), .A(divq[7]), .B(n_7819), .Z(n_25823));
	notech_reg_set divq_reg_8(.CP(n_63652), .D(n_25831), .SD(1'b1), .Q(divq[
		8]));
	notech_mux2 i_8645(.S(n_56397), .A(divq[8]), .B(n_7824), .Z(n_25831));
	notech_reg_set divq_reg_9(.CP(n_63652), .D(n_25842), .SD(1'b1), .Q(divq[
		9]));
	notech_mux2 i_8653(.S(n_56397), .A(divq[9]), .B(n_7829), .Z(n_25842));
	notech_reg_set divq_reg_10(.CP(n_63652), .D(n_25848), .SD(1'b1), .Q(divq
		[10]));
	notech_mux2 i_8661(.S(n_56397), .A(divq[10]), .B(n_7834), .Z(n_25848));
	notech_reg_set divq_reg_11(.CP(n_63652), .D(n_25854), .SD(1'b1), .Q(divq
		[11]));
	notech_mux2 i_8669(.S(n_56397), .A(divq[11]), .B(n_7839), .Z(n_25854));
	notech_reg_set divq_reg_12(.CP(n_63652), .D(n_25860), .SD(1'b1), .Q(divq
		[12]));
	notech_mux2 i_8677(.S(n_56397), .A(divq[12]), .B(n_215266559), .Z(n_25860
		));
	notech_reg_set divq_reg_13(.CP(n_63652), .D(n_25866), .SD(1'b1), .Q(divq
		[13]));
	notech_mux2 i_8685(.S(n_56397), .A(divq[13]), .B(n_187762904), .Z(n_25866
		));
	notech_reg_set divq_reg_14(.CP(n_63652), .D(n_25872), .SD(1'b1), .Q(divq
		[14]));
	notech_mux2 i_8693(.S(n_56397), .A(divq[14]), .B(n_7854), .Z(n_25872));
	notech_reg_set divq_reg_15(.CP(n_63652), .D(n_25878), .SD(1'b1), .Q(divq
		[15]));
	notech_mux2 i_8701(.S(n_56397), .A(divq[15]), .B(n_214466554), .Z(n_25878
		));
	notech_reg_set divq_reg_16(.CP(n_63652), .D(n_25884), .SD(1'b1), .Q(divq
		[16]));
	notech_mux2 i_8709(.S(n_56399), .A(divq[16]), .B(n_7864), .Z(n_25884));
	notech_reg_set divq_reg_17(.CP(n_63652), .D(n_25890), .SD(1'b1), .Q(divq
		[17]));
	notech_mux2 i_8717(.S(n_56399), .A(divq[17]), .B(n_7869), .Z(n_25890));
	notech_reg_set divq_reg_18(.CP(n_63652), .D(n_25897), .SD(1'b1), .Q(divq
		[18]));
	notech_mux2 i_8725(.S(n_56399), .A(divq[18]), .B(n_7874), .Z(n_25897));
	notech_reg_set divq_reg_19(.CP(n_63652), .D(n_25903), .SD(1'b1), .Q(divq
		[19]));
	notech_mux2 i_8733(.S(n_56399), .A(divq[19]), .B(n_7879), .Z(n_25903));
	notech_reg_set divq_reg_20(.CP(n_63652), .D(n_25909), .SD(1'b1), .Q(divq
		[20]));
	notech_mux2 i_8741(.S(n_56399), .A(divq[20]), .B(n_7884), .Z(n_25909));
	notech_reg_set divq_reg_21(.CP(n_63652), .D(n_25919), .SD(1'b1), .Q(divq
		[21]));
	notech_mux2 i_8749(.S(n_56399), .A(divq[21]), .B(n_7889), .Z(n_25919));
	notech_reg_set divq_reg_22(.CP(n_63576), .D(n_25925), .SD(1'b1), .Q(divq
		[22]));
	notech_mux2 i_8757(.S(n_56399), .A(divq[22]), .B(n_7894), .Z(n_25925));
	notech_reg_set divq_reg_23(.CP(n_63576), .D(n_25931), .SD(1'b1), .Q(divq
		[23]));
	notech_mux2 i_8765(.S(n_56399), .A(divq[23]), .B(n_7899), .Z(n_25931));
	notech_reg_set divq_reg_24(.CP(n_63576), .D(n_25937), .SD(1'b1), .Q(divq
		[24]));
	notech_mux2 i_8773(.S(n_56399), .A(divq[24]), .B(n_7904), .Z(n_25937));
	notech_reg_set divq_reg_25(.CP(n_63576), .D(n_25943), .SD(1'b1), .Q(divq
		[25]));
	notech_mux2 i_8781(.S(n_56399), .A(divq[25]), .B(n_7909), .Z(n_25943));
	notech_reg_set divq_reg_26(.CP(n_63576), .D(n_25949), .SD(1'b1), .Q(divq
		[26]));
	notech_mux2 i_8789(.S(n_56399), .A(divq[26]), .B(n_7914), .Z(n_25949));
	notech_reg_set divq_reg_27(.CP(n_63576), .D(n_25955), .SD(1'b1), .Q(divq
		[27]));
	notech_mux2 i_8797(.S(n_56399), .A(divq[27]), .B(n_7919), .Z(n_25955));
	notech_reg_set divq_reg_28(.CP(n_63576), .D(n_25961), .SD(1'b1), .Q(divq
		[28]));
	notech_mux2 i_8805(.S(n_56399), .A(divq[28]), .B(n_7924), .Z(n_25961));
	notech_reg_set divq_reg_29(.CP(n_63576), .D(n_25967), .SD(1'b1), .Q(divq
		[29]));
	notech_mux2 i_8813(.S(n_56399), .A(divq[29]), .B(n_7929), .Z(n_25967));
	notech_reg_set divq_reg_30(.CP(n_63576), .D(n_25973), .SD(1'b1), .Q(divq
		[30]));
	notech_mux2 i_8821(.S(n_56399), .A(divq[30]), .B(n_7934), .Z(n_25973));
	notech_reg_set divq_reg_31(.CP(n_63576), .D(n_25979), .SD(1'b1), .Q(divq
		[31]));
	notech_mux2 i_8829(.S(n_56399), .A(divq[31]), .B(n_7939), .Z(n_25979));
	notech_reg_set divq_reg_32(.CP(n_63500), .D(n_25985), .SD(1'b1), .Q(divq
		[32]));
	notech_mux2 i_8837(.S(n_56392), .A(divq[32]), .B(n_7944), .Z(n_25985));
	notech_reg_set divq_reg_33(.CP(n_63576), .D(n_25991), .SD(1'b1), .Q(divq
		[33]));
	notech_mux2 i_8845(.S(n_56392), .A(divq[33]), .B(n_31102), .Z(n_25991)
		);
	notech_reg_set divq_reg_34(.CP(n_63582), .D(n_25997), .SD(1'b1), .Q(divq
		[34]));
	notech_mux2 i_8853(.S(n_56392), .A(divq[34]), .B(n_31103), .Z(n_25997)
		);
	notech_reg_set divq_reg_35(.CP(n_63502), .D(n_26003), .SD(1'b1), .Q(divq
		[35]));
	notech_mux2 i_8861(.S(n_56392), .A(divq[35]), .B(n_31104), .Z(n_26003)
		);
	notech_reg_set divq_reg_36(.CP(n_63502), .D(n_26009), .SD(1'b1), .Q(divq
		[36]));
	notech_mux2 i_8870(.S(n_56392), .A(divq[36]), .B(n_31105), .Z(n_26009)
		);
	notech_reg_set divq_reg_37(.CP(n_63502), .D(n_26015), .SD(1'b1), .Q(divq
		[37]));
	notech_mux2 i_8878(.S(n_56392), .A(divq[37]), .B(n_31106), .Z(n_26015)
		);
	notech_reg_set divq_reg_38(.CP(n_63502), .D(n_26021), .SD(1'b1), .Q(divq
		[38]));
	notech_mux2 i_8886(.S(n_56392), .A(divq[38]), .B(n_31107), .Z(n_26021)
		);
	notech_reg_set divq_reg_39(.CP(n_63502), .D(n_26027), .SD(1'b1), .Q(divq
		[39]));
	notech_mux2 i_8894(.S(n_56392), .A(divq[39]), .B(n_31108), .Z(n_26027)
		);
	notech_reg_set divq_reg_40(.CP(n_63502), .D(n_26034), .SD(1'b1), .Q(divq
		[40]));
	notech_mux2 i_8902(.S(n_56392), .A(divq[40]), .B(n_31109), .Z(n_26034)
		);
	notech_reg_set divq_reg_41(.CP(n_63502), .D(n_26040), .SD(1'b1), .Q(divq
		[41]));
	notech_mux2 i_8910(.S(n_56392), .A(divq[41]), .B(n_31110), .Z(n_26040)
		);
	notech_reg_set divq_reg_42(.CP(n_63502), .D(n_26050), .SD(1'b1), .Q(divq
		[42]));
	notech_mux2 i_8918(.S(n_56392), .A(divq[42]), .B(n_31111), .Z(n_26050)
		);
	notech_reg_set divq_reg_43(.CP(n_63502), .D(n_26056), .SD(1'b1), .Q(divq
		[43]));
	notech_mux2 i_8926(.S(n_56392), .A(divq[43]), .B(n_31112), .Z(n_26056)
		);
	notech_reg_set divq_reg_44(.CP(n_63502), .D(n_26065), .SD(1'b1), .Q(divq
		[44]));
	notech_mux2 i_8934(.S(n_56392), .A(divq[44]), .B(n_31113), .Z(n_26065)
		);
	notech_reg_set divq_reg_45(.CP(n_63584), .D(n_26071), .SD(1'b1), .Q(divq
		[45]));
	notech_mux2 i_8942(.S(n_56392), .A(divq[45]), .B(n_31114), .Z(n_26071)
		);
	notech_reg_set divq_reg_46(.CP(n_63584), .D(n_26077), .SD(1'b1), .Q(divq
		[46]));
	notech_mux2 i_8951(.S(n_56392), .A(divq[46]), .B(n_31115), .Z(n_26077)
		);
	notech_reg_set divq_reg_47(.CP(n_63584), .D(n_26083), .SD(1'b1), .Q(divq
		[47]));
	notech_mux2 i_8959(.S(n_56392), .A(divq[47]), .B(n_31116), .Z(n_26083)
		);
	notech_reg_set divq_reg_48(.CP(n_63584), .D(n_26090), .SD(1'b1), .Q(divq
		[48]));
	notech_mux2 i_8967(.S(n_56394), .A(divq[48]), .B(n_31117), .Z(n_26090)
		);
	notech_reg_set divq_reg_49(.CP(n_63584), .D(n_26096), .SD(1'b1), .Q(divq
		[49]));
	notech_mux2 i_8975(.S(n_56394), .A(divq[49]), .B(n_31120), .Z(n_26096)
		);
	notech_reg_set divq_reg_50(.CP(n_63584), .D(n_26102), .SD(1'b1), .Q(divq
		[50]));
	notech_mux2 i_8983(.S(n_56394), .A(divq[50]), .B(n_31121), .Z(n_26102)
		);
	notech_reg_set divq_reg_51(.CP(n_63584), .D(n_26108), .SD(1'b1), .Q(divq
		[51]));
	notech_mux2 i_8991(.S(n_56394), .A(divq[51]), .B(n_31124), .Z(n_26108)
		);
	notech_reg_set divq_reg_52(.CP(n_63584), .D(n_26114), .SD(1'b1), .Q(divq
		[52]));
	notech_mux2 i_8999(.S(n_56394), .A(divq[52]), .B(n_31127), .Z(n_26114)
		);
	notech_reg_set divq_reg_53(.CP(n_63584), .D(n_26120), .SD(1'b1), .Q(divq
		[53]));
	notech_mux2 i_9007(.S(n_56394), .A(divq[53]), .B(n_31128), .Z(n_26120)
		);
	notech_reg_set divq_reg_54(.CP(n_63584), .D(n_26126), .SD(1'b1), .Q(divq
		[54]));
	notech_mux2 i_9015(.S(n_56394), .A(divq[54]), .B(n_31129), .Z(n_26126)
		);
	notech_reg_set divq_reg_55(.CP(n_63584), .D(n_26132), .SD(1'b1), .Q(divq
		[55]));
	notech_mux2 i_9023(.S(n_56394), .A(divq[55]), .B(n_31130), .Z(n_26132)
		);
	notech_reg_set divq_reg_56(.CP(n_63584), .D(n_26139), .SD(1'b1), .Q(divq
		[56]));
	notech_mux2 i_9031(.S(n_56394), .A(divq[56]), .B(n_31131), .Z(n_26139)
		);
	notech_reg_set divq_reg_57(.CP(n_63584), .D(n_26145), .SD(1'b1), .Q(divq
		[57]));
	notech_mux2 i_9039(.S(n_56394), .A(divq[57]), .B(n_31132), .Z(n_26145)
		);
	notech_reg_set divq_reg_58(.CP(n_63584), .D(n_26151), .SD(1'b1), .Q(divq
		[58]));
	notech_mux2 i_9047(.S(n_56394), .A(divq[58]), .B(n_31133), .Z(n_26151)
		);
	notech_reg_set divq_reg_59(.CP(n_63584), .D(n_26157), .SD(1'b1), .Q(divq
		[59]));
	notech_mux2 i_9055(.S(n_56394), .A(divq[59]), .B(n_31134), .Z(n_26157)
		);
	notech_reg_set divq_reg_60(.CP(n_63584), .D(n_26163), .SD(1'b1), .Q(divq
		[60]));
	notech_mux2 i_9063(.S(n_56394), .A(divq[60]), .B(n_31135), .Z(n_26163)
		);
	notech_reg_set divq_reg_61(.CP(n_63584), .D(n_26169), .SD(1'b1), .Q(divq
		[61]));
	notech_mux2 i_9071(.S(n_56394), .A(divq[61]), .B(n_31136), .Z(n_26169)
		);
	notech_reg_set divq_reg_62(.CP(n_63584), .D(n_26175), .SD(1'b1), .Q(divq
		[62]));
	notech_mux2 i_9079(.S(n_56394), .A(divq[62]), .B(n_31137), .Z(n_26175)
		);
	notech_nand3 i_28272(.A(n_63720), .B(n_63764), .C(opa[5]), .Z(n_31126)
		);
	notech_reg_set divq_reg_63(.CP(n_63584), .D(n_26181), .SD(1'b1), .Q(divq
		[63]));
	notech_mux2 i_9087(.S(n_56394), .A(divq[63]), .B(n_176994252), .Z(n_26181
		));
	notech_nand3 i_28273(.A(n_63720), .B(n_63764), .C(opb[5]), .Z(n_31125)
		);
	notech_reg_set divr_reg_0(.CP(n_63656), .D(n_26187), .SD(1'b1), .Q(divr[
		0]));
	notech_mux2 i_9095(.S(n_56440), .A(divr[0]), .B(n_16502), .Z(n_26187));
	notech_nand3 i_28275(.A(n_63720), .B(n_61928), .C(opb[5]), .Z(n_31123)
		);
	notech_reg_set divr_reg_1(.CP(n_63582), .D(n_26193), .SD(1'b1), .Q(divr[
		1]));
	notech_mux2 i_9103(.S(n_56440), .A(divr[1]), .B(n_16507), .Z(n_26193));
	notech_nand3 i_28276(.A(n_63698), .B(n_61928), .C(opa[5]), .Z(n_31122)
		);
	notech_reg_set divr_reg_2(.CP(n_63656), .D(n_26199), .SD(1'b1), .Q(divr[
		2]));
	notech_mux2 i_9111(.S(n_56440), .A(divr[2]), .B(n_16512), .Z(n_26199));
	notech_nand2 i_28279(.A(n_63776), .B(opc_10[5]), .Z(n_31119));
	notech_reg_set divr_reg_3(.CP(n_63656), .D(n_26205), .SD(1'b1), .Q(divr[
		3]));
	notech_mux2 i_9119(.S(n_56440), .A(divr[3]), .B(n_16517), .Z(n_26205));
	notech_nand2 i_28280(.A(n_63776), .B(opc[5]), .Z(n_31118));
	notech_reg_set divr_reg_4(.CP(n_63656), .D(n_26211), .SD(1'b1), .Q(divr[
		4]));
	notech_mux2 i_9127(.S(n_56440), .A(divr[4]), .B(n_16522), .Z(n_26211));
	notech_nao3 i_28299(.A(n_63776), .B(opa[5]), .C(\opcode[1] ), .Z(n_31099
		));
	notech_reg_set divr_reg_5(.CP(n_63656), .D(n_26217), .SD(1'b1), .Q(divr[
		5]));
	notech_mux2 i_9135(.S(n_56440), .A(divr[5]), .B(n_16527), .Z(n_26217));
	notech_nao3 i_28300(.A(n_61928), .B(opa[5]), .C(\opcode[1] ), .Z(n_31098
		));
	notech_reg_set divr_reg_6(.CP(n_63656), .D(n_26223), .SD(1'b1), .Q(divr[
		6]));
	notech_mux2 i_9143(.S(n_56440), .A(divr[6]), .B(n_16532), .Z(n_26223));
	notech_nand3 i_28323(.A(n_63698), .B(n_63734), .C(opa[4]), .Z(n_31075)
		);
	notech_reg_set divr_reg_7(.CP(n_63656), .D(n_26229), .SD(1'b1), .Q(divr[
		7]));
	notech_mux2 i_9151(.S(n_56440), .A(divr[7]), .B(n_16537), .Z(n_26229));
	notech_nand3 i_28324(.A(n_63698), .B(n_63734), .C(opb[4]), .Z(n_31074)
		);
	notech_reg_set divr_reg_8(.CP(n_63656), .D(n_26235), .SD(1'b1), .Q(divr[
		8]));
	notech_mux2 i_9159(.S(n_56440), .A(divr[8]), .B(n_16542), .Z(n_26235));
	notech_nand3 i_28326(.A(n_63698), .B(n_61930), .C(opb[4]), .Z(n_31072)
		);
	notech_reg_set divr_reg_9(.CP(n_63656), .D(n_26241), .SD(1'b1), .Q(divr[
		9]));
	notech_mux2 i_9167(.S(n_56440), .A(divr[9]), .B(n_16547), .Z(n_26241));
	notech_nand3 i_28327(.A(n_63698), .B(n_61928), .C(opa[4]), .Z(n_31071)
		);
	notech_reg_set divr_reg_10(.CP(n_63656), .D(n_26247), .SD(1'b1), .Q(divr
		[10]));
	notech_mux2 i_9175(.S(n_56440), .A(divr[10]), .B(n_188562912), .Z(n_26247
		));
	notech_nand2 i_28330(.A(n_63776), .B(opc_10[4]), .Z(n_31068));
	notech_reg_set divr_reg_11(.CP(n_63656), .D(n_26253), .SD(1'b1), .Q(divr
		[11]));
	notech_mux2 i_9183(.S(n_56440), .A(divr[11]), .B(n_216866571), .Z(n_26253
		));
	notech_nand2 i_28331(.A(n_63776), .B(opc[4]), .Z(n_31067));
	notech_reg_set divr_reg_12(.CP(n_63656), .D(n_26259), .SD(1'b1), .Q(divr
		[12]));
	notech_mux2 i_9191(.S(n_56440), .A(divr[12]), .B(n_216466567), .Z(n_26259
		));
	notech_nao3 i_28350(.A(n_63776), .B(opa[4]), .C(\opcode[1] ), .Z(n_31048
		));
	notech_reg_set divr_reg_13(.CP(n_63656), .D(n_26265), .SD(1'b1), .Q(divr
		[13]));
	notech_mux2 i_9199(.S(n_56440), .A(divr[13]), .B(n_188162908), .Z(n_26265
		));
	notech_nao3 i_28351(.A(n_61928), .B(opa[4]), .C(\opcode[1] ), .Z(n_31047
		));
	notech_reg_set divr_reg_14(.CP(n_63656), .D(n_26274), .SD(1'b1), .Q(divr
		[14]));
	notech_mux2 i_9207(.S(n_56440), .A(divr[14]), .B(n_16572), .Z(n_26274)
		);
	notech_reg_set divr_reg_15(.CP(n_63656), .D(n_26284), .SD(1'b1), .Q(divr
		[15]));
	notech_mux2 i_9216(.S(n_56440), .A(divr[15]), .B(n_215766563), .Z(n_26284
		));
	notech_reg_set divr_reg_16(.CP(n_63656), .D(n_26290), .SD(1'b1), .Q(divr
		[16]));
	notech_mux2 i_9225(.S(n_56442), .A(divr[16]), .B(n_16582), .Z(n_26290)
		);
	notech_reg_set divr_reg_17(.CP(n_63656), .D(n_26296), .SD(1'b1), .Q(divr
		[17]));
	notech_mux2 i_9233(.S(n_56442), .A(divr[17]), .B(n_16587), .Z(n_26296)
		);
	notech_reg_set divr_reg_18(.CP(n_63656), .D(n_26302), .SD(1'b1), .Q(divr
		[18]));
	notech_mux2 i_9241(.S(n_56442), .A(divr[18]), .B(n_16592), .Z(n_26302)
		);
	notech_reg_set divr_reg_19(.CP(n_63656), .D(n_26308), .SD(1'b1), .Q(divr
		[19]));
	notech_mux2 i_9249(.S(n_56442), .A(divr[19]), .B(n_16597), .Z(n_26308)
		);
	notech_reg_set divr_reg_20(.CP(n_63582), .D(n_26314), .SD(1'b1), .Q(divr
		[20]));
	notech_mux2 i_9257(.S(n_56442), .A(divr[20]), .B(n_16602), .Z(n_26314)
		);
	notech_reg_set divr_reg_21(.CP(n_63582), .D(n_26320), .SD(1'b1), .Q(divr
		[21]));
	notech_mux2 i_9265(.S(n_56442), .A(divr[21]), .B(n_16607), .Z(n_26320)
		);
	notech_reg_set divr_reg_22(.CP(n_63582), .D(n_26326), .SD(1'b1), .Q(divr
		[22]));
	notech_mux2 i_9273(.S(n_56442), .A(divr[22]), .B(n_16612), .Z(n_26326)
		);
	notech_reg_set divr_reg_23(.CP(n_63582), .D(n_26332), .SD(1'b1), .Q(divr
		[23]));
	notech_mux2 i_9281(.S(n_56442), .A(divr[23]), .B(n_16617), .Z(n_26332)
		);
	notech_reg_set divr_reg_24(.CP(n_63582), .D(n_26338), .SD(1'b1), .Q(divr
		[24]));
	notech_mux2 i_9289(.S(n_56442), .A(divr[24]), .B(n_16622), .Z(n_26338)
		);
	notech_reg_set divr_reg_25(.CP(n_63582), .D(n_26344), .SD(1'b1), .Q(divr
		[25]));
	notech_mux2 i_9297(.S(n_56442), .A(divr[25]), .B(n_16627), .Z(n_26344)
		);
	notech_reg_set divr_reg_26(.CP(n_63582), .D(n_26350), .SD(1'b1), .Q(divr
		[26]));
	notech_mux2 i_9305(.S(n_56442), .A(divr[26]), .B(n_16632), .Z(n_26350)
		);
	notech_reg_set divr_reg_27(.CP(n_63582), .D(n_26356), .SD(1'b1), .Q(divr
		[27]));
	notech_mux2 i_9313(.S(n_56442), .A(divr[27]), .B(n_16637), .Z(n_26356)
		);
	notech_reg_set divr_reg_28(.CP(n_63582), .D(n_26362), .SD(1'b1), .Q(divr
		[28]));
	notech_mux2 i_9321(.S(n_56442), .A(divr[28]), .B(n_16642), .Z(n_26362)
		);
	notech_reg_set divr_reg_29(.CP(n_63582), .D(n_26368), .SD(1'b1), .Q(divr
		[29]));
	notech_mux2 i_9329(.S(n_56442), .A(divr[29]), .B(n_16647), .Z(n_26368)
		);
	notech_reg_set divr_reg_30(.CP(n_63502), .D(n_26374), .SD(1'b1), .Q(divr
		[30]));
	notech_mux2 i_9337(.S(n_56442), .A(divr[30]), .B(n_16652), .Z(n_26374)
		);
	notech_or2 i_24749487(.A(n_75322856), .B(n_26275), .Z(n_2057));
	notech_reg_set divr_reg_31(.CP(n_63502), .D(n_26380), .SD(1'b1), .Q(divr
		[31]));
	notech_mux2 i_9345(.S(n_56442), .A(divr[31]), .B(n_16657), .Z(n_26380)
		);
	notech_reg_set divr_reg_32(.CP(n_63586), .D(n_26387), .SD(1'b1), .Q(divr
		[32]));
	notech_mux2 i_9353(.S(n_56435), .A(divr[32]), .B(n_16662), .Z(n_26387)
		);
	notech_reg_set divr_reg_33(.CP(n_63504), .D(n_26395), .SD(1'b1), .Q(divr
		[33]));
	notech_mux2 i_9361(.S(n_56435), .A(divr[33]), .B(n_16667), .Z(n_26395)
		);
	notech_reg_set divr_reg_34(.CP(n_63504), .D(n_26404), .SD(1'b1), .Q(divr
		[34]));
	notech_mux2 i_9369(.S(n_56435), .A(divr[34]), .B(n_16672), .Z(n_26404)
		);
	notech_reg_set divr_reg_35(.CP(n_63504), .D(n_26410), .SD(1'b1), .Q(divr
		[35]));
	notech_mux2 i_9377(.S(n_56435), .A(divr[35]), .B(n_16677), .Z(n_26410)
		);
	notech_nao3 i_25249482(.A(n_63776), .B(opc_10[3]), .C(n_26271), .Z(n_2052
		));
	notech_reg_set divr_reg_36(.CP(n_63504), .D(n_26416), .SD(1'b1), .Q(divr
		[36]));
	notech_mux2 i_9385(.S(n_56435), .A(divr[36]), .B(n_16682), .Z(n_26416)
		);
	notech_reg_set divr_reg_37(.CP(n_63504), .D(n_26422), .SD(1'b1), .Q(divr
		[37]));
	notech_mux2 i_9393(.S(n_56435), .A(divr[37]), .B(n_16687), .Z(n_26422)
		);
	notech_reg_set divr_reg_38(.CP(n_63504), .D(n_26428), .SD(1'b1), .Q(divr
		[38]));
	notech_mux2 i_9402(.S(n_56435), .A(divr[38]), .B(n_16692), .Z(n_26428)
		);
	notech_reg_set divr_reg_39(.CP(n_63504), .D(n_26434), .SD(1'b1), .Q(divr
		[39]));
	notech_mux2 i_9410(.S(n_56435), .A(divr[39]), .B(n_16697), .Z(n_26434)
		);
	notech_reg_set divr_reg_40(.CP(n_63504), .D(n_26440), .SD(1'b1), .Q(divr
		[40]));
	notech_mux2 i_9420(.S(n_56435), .A(divr[40]), .B(n_16702), .Z(n_26440)
		);
	notech_or2 i_25749477(.A(n_338361011), .B(n_332460952), .Z(n_2045));
	notech_reg_set divr_reg_41(.CP(n_63504), .D(n_26446), .SD(1'b1), .Q(divr
		[41]));
	notech_mux2 i_9430(.S(n_56435), .A(divr[41]), .B(n_16707), .Z(n_26446)
		);
	notech_reg_set divr_reg_42(.CP(n_63504), .D(n_26452), .SD(1'b1), .Q(divr
		[42]));
	notech_mux2 i_9438(.S(n_56435), .A(divr[42]), .B(n_16712), .Z(n_26452)
		);
	notech_reg_set divr_reg_43(.CP(n_63586), .D(n_26458), .SD(1'b1), .Q(divr
		[43]));
	notech_mux2 i_9446(.S(n_56435), .A(divr[43]), .B(n_16717), .Z(n_26458)
		);
	notech_reg_set divr_reg_44(.CP(n_63586), .D(n_26464), .SD(1'b1), .Q(divr
		[44]));
	notech_mux2 i_9454(.S(n_56435), .A(divr[44]), .B(n_16722), .Z(n_26464)
		);
	notech_reg_set divr_reg_45(.CP(n_63586), .D(n_26470), .SD(1'b1), .Q(divr
		[45]));
	notech_mux2 i_9462(.S(n_56435), .A(divr[45]), .B(n_16727), .Z(n_26470)
		);
	notech_reg_set divr_reg_46(.CP(n_63586), .D(n_26476), .SD(1'b1), .Q(divr
		[46]));
	notech_mux2 i_9470(.S(n_56435), .A(divr[46]), .B(n_16732), .Z(n_26476)
		);
	notech_reg_set divr_reg_47(.CP(n_63586), .D(n_26482), .SD(1'b1), .Q(divr
		[47]));
	notech_mux2 i_9478(.S(n_56435), .A(divr[47]), .B(n_16737), .Z(n_26482)
		);
	notech_reg_set divr_reg_48(.CP(n_63586), .D(n_26488), .SD(1'b1), .Q(divr
		[48]));
	notech_mux2 i_9486(.S(n_56437), .A(divr[48]), .B(n_16742), .Z(n_26488)
		);
	notech_reg_set divr_reg_49(.CP(n_63586), .D(n_26494), .SD(1'b1), .Q(divr
		[49]));
	notech_mux2 i_9494(.S(n_56437), .A(divr[49]), .B(n_16747), .Z(n_26494)
		);
	notech_and2 i_118648595(.A(n_338061008), .B(n_1634), .Z(n_2034));
	notech_reg_set divr_reg_50(.CP(n_63586), .D(n_26500), .SD(1'b1), .Q(divr
		[50]));
	notech_mux2 i_9502(.S(n_56437), .A(divr[50]), .B(n_16752), .Z(n_26500)
		);
	notech_nand3 i_118048597(.A(n_28551), .B(n_28558), .C(n_28552), .Z(n_203360404
		));
	notech_reg_set divr_reg_51(.CP(n_63586), .D(n_26506), .SD(1'b1), .Q(divr
		[51]));
	notech_mux2 i_9510(.S(n_56437), .A(divr[51]), .B(n_16757), .Z(n_26506)
		);
	notech_nand3 i_149724(.A(n_83739557), .B(n_27379), .C(n_83839558), .Z(n_203260403
		));
	notech_reg_set divr_reg_52(.CP(n_63586), .D(n_26512), .SD(1'b1), .Q(divr
		[52]));
	notech_mux2 i_9518(.S(n_56437), .A(divr[52]), .B(n_16762), .Z(n_26512)
		);
	notech_nao3 i_21158216(.A(n_57656), .B(n_336260990), .C(n_336460992), .Z
		(n_30694));
	notech_reg_set divr_reg_53(.CP(n_63586), .D(n_26518), .SD(1'b1), .Q(divr
		[53]));
	notech_mux2 i_9526(.S(n_56437), .A(divr[53]), .B(n_16767), .Z(n_26518)
		);
	notech_reg_set divr_reg_54(.CP(n_63586), .D(n_26524), .SD(1'b1), .Q(divr
		[54]));
	notech_mux2 i_9534(.S(n_56437), .A(divr[54]), .B(n_16772), .Z(n_26524)
		);
	notech_and3 i_159151499(.A(n_2021), .B(n_2020), .C(n_2028), .Z(n_2029)
		);
	notech_reg_set divr_reg_55(.CP(n_63586), .D(n_26530), .SD(1'b1), .Q(divr
		[55]));
	notech_mux2 i_9542(.S(n_56437), .A(divr[55]), .B(n_16777), .Z(n_26530)
		);
	notech_and4 i_159051500(.A(n_202660402), .B(n_202560401), .C(n_2023), .D
		(n_1948), .Z(n_2028));
	notech_reg_set divr_reg_56(.CP(n_63586), .D(n_26536), .SD(1'b1), .Q(divr
		[56]));
	notech_mux2 i_9550(.S(n_56437), .A(divr[56]), .B(n_16782), .Z(n_26536)
		);
	notech_reg_set divr_reg_57(.CP(n_63586), .D(n_26542), .SD(1'b1), .Q(divr
		[57]));
	notech_mux2 i_9558(.S(n_56437), .A(divr[57]), .B(n_16787), .Z(n_26542)
		);
	notech_ao4 i_158451506(.A(n_126826595), .B(n_58920), .C(n_126726594), .D
		(n_58438), .Z(n_202660402));
	notech_reg_set divr_reg_58(.CP(n_63586), .D(n_26548), .SD(1'b1), .Q(divr
		[58]));
	notech_mux2 i_9566(.S(n_56437), .A(divr[58]), .B(n_16792), .Z(n_26548)
		);
	notech_ao4 i_158351507(.A(n_337761005), .B(n_60510), .C(n_55966), .D(n_33110
		), .Z(n_202560401));
	notech_reg_set divr_reg_59(.CP(n_63586), .D(n_26554), .SD(1'b1), .Q(divr
		[59]));
	notech_mux2 i_9574(.S(n_56437), .A(divr[59]), .B(n_16797), .Z(n_26554)
		);
	notech_reg_set divr_reg_60(.CP(n_63586), .D(n_26560), .SD(1'b1), .Q(divr
		[60]));
	notech_mux2 i_9582(.S(n_56437), .A(divr[60]), .B(n_16802), .Z(n_26560)
		);
	notech_ao4 i_158251508(.A(n_55975), .B(n_32084), .C(n_55955), .D(n_31018
		), .Z(n_2023));
	notech_reg_set divr_reg_61(.CP(n_63504), .D(n_26566), .SD(1'b1), .Q(divr
		[61]));
	notech_mux2 i_9590(.S(n_56437), .A(divr[61]), .B(n_16807), .Z(n_26566)
		);
	notech_reg_set divr_reg_62(.CP(n_63504), .D(n_26572), .SD(1'b1), .Q(divr
		[62]));
	notech_mux2 i_9598(.S(n_56437), .A(divr[62]), .B(n_16812), .Z(n_26572)
		);
	notech_ao4 i_158651504(.A(n_337861006), .B(n_31501), .C(n_55946), .D(n_31533
		), .Z(n_2021));
	notech_reg_set divr_reg_63(.CP(n_63506), .D(n_26578), .SD(1'b1), .Q(divr
		[63]));
	notech_mux2 i_9606(.S(n_56437), .A(divr[63]), .B(n_16817), .Z(n_26578)
		);
	notech_ao4 i_158551505(.A(n_126926596), .B(n_33172), .C(n_101026337), .D
		(n_127026597), .Z(n_2020));
	notech_reg sign_div_reg(.CP(n_63506), .D(n_26584), .CD(n_62379), .Q(sign_div
		));
	notech_mux2 i_9614(.S(n_339389278), .A(n_30736), .B(sign_div), .Z(n_26584
		));
	notech_reg_set opc_reg_0(.CP(n_63506), .D(n_26591), .SD(1'b1), .Q(opc[0]
		));
	notech_mux2 i_9622(.S(\nbus_11289[0] ), .A(opc[0]), .B(n_9816), .Z(n_26591
		));
	notech_reg_set opc_reg_1(.CP(n_63506), .D(n_26597), .SD(1'b1), .Q(opc[1]
		));
	notech_mux2 i_9630(.S(\nbus_11289[0] ), .A(opc[1]), .B(n_31140), .Z(n_26597
		));
	notech_nand3 i_137751713(.A(n_2015), .B(n_2014), .C(n_201360398), .Z(n_2017
		));
	notech_reg_set opc_reg_2(.CP(n_63506), .D(n_26605), .SD(1'b1), .Q(opc[2]
		));
	notech_mux2 i_9638(.S(\nbus_11289[0] ), .A(opc[2]), .B(n_9826), .Z(n_26605
		));
	notech_reg_set opc_reg_3(.CP(n_63506), .D(n_26611), .SD(1'b1), .Q(opc[3]
		));
	notech_mux2 i_9646(.S(\nbus_11289[0] ), .A(opc[3]), .B(n_31141), .Z(n_26611
		));
	notech_ao4 i_137151719(.A(n_124626573), .B(n_58429), .C(n_337561003), .D
		(n_60519), .Z(n_2015));
	notech_reg_set opc_reg_4(.CP(n_63506), .D(n_26617), .SD(1'b1), .Q(opc[4]
		));
	notech_mux2 i_9654(.S(\nbus_11289[0] ), .A(opc[4]), .B(n_30427), .Z(n_26617
		));
	notech_ao4 i_137051720(.A(n_55913), .B(n_33109), .C(n_55793), .D(n_33107
		), .Z(n_2014));
	notech_reg_set opc_reg_5(.CP(n_63506), .D(n_26625), .SD(1'b1), .Q(opc[5]
		));
	notech_mux2 i_9662(.S(n_31142), .A(opc[5]), .B(n_9841), .Z(n_26625));
	notech_ao4 i_137451716(.A(n_61092), .B(n_30830), .C(n_57006), .D(n_31532
		), .Z(n_201360398));
	notech_reg_set opc_reg_6(.CP(n_63506), .D(n_26633), .SD(1'b1), .Q(opc[6]
		));
	notech_mux2 i_9670(.S(n_31142), .A(opc[6]), .B(n_9846), .Z(n_26633));
	notech_nand2 i_137651714(.A(n_201160396), .B(n_2010), .Z(n_201260397));
	notech_reg_set opc_reg_7(.CP(n_63506), .D(n_26640), .SD(1'b1), .Q(opc[7]
		));
	notech_mux2 i_9678(.S(n_31142), .A(opc[7]), .B(n_9851), .Z(n_26640));
	notech_ao4 i_137351717(.A(n_31500), .B(n_328660914), .C(n_124726574), .D
		(n_33171), .Z(n_201160396));
	notech_reg_set opc_reg_8(.CP(n_63506), .D(n_26646), .SD(1'b1), .Q(opc[8]
		));
	notech_mux2 i_9686(.S(\nbus_11289[8] ), .A(opc[8]), .B(n_9856), .Z(n_26646
		));
	notech_ao4 i_137251718(.A(n_106826395), .B(n_124826575), .C(n_124526572)
		, .D(n_58893), .Z(n_2010));
	notech_reg_set opc_reg_9(.CP(n_63506), .D(n_26652), .SD(1'b1), .Q(opc[9]
		));
	notech_mux2 i_9694(.S(\nbus_11289[8] ), .A(opc[9]), .B(n_9861), .Z(n_26652
		));
	notech_reg_set opc_reg_10(.CP(n_63506), .D(n_26658), .SD(1'b1), .Q(opc[
		10]));
	notech_mux2 i_9702(.S(\nbus_11289[8] ), .A(opc[10]), .B(n_9866), .Z(n_26658
		));
	notech_reg_set opc_reg_11(.CP(n_63506), .D(n_26666), .SD(1'b1), .Q(opc[
		11]));
	notech_mux2 i_9710(.S(\nbus_11289[8] ), .A(opc[11]), .B(n_9871), .Z(n_26666
		));
	notech_nand3 i_115851930(.A(n_200460393), .B(n_200360392), .C(n_2002), .Z
		(n_200660395));
	notech_reg_set opc_reg_12(.CP(n_63506), .D(n_26672), .SD(1'b1), .Q(opc[
		12]));
	notech_mux2 i_9718(.S(\nbus_11289[8] ), .A(opc[12]), .B(n_9876), .Z(n_26672
		));
	notech_reg_set opc_reg_13(.CP(n_63506), .D(n_26678), .SD(1'b1), .Q(opc[
		13]));
	notech_mux2 i_9726(.S(\nbus_11289[8] ), .A(opc[13]), .B(n_9881), .Z(n_26678
		));
	notech_ao4 i_115251936(.A(n_122726554), .B(n_58420), .C(n_337361001), .D
		(n_60528), .Z(n_200460393));
	notech_reg_set opc_reg_14(.CP(n_63506), .D(n_26684), .SD(1'b1), .Q(opc[
		14]));
	notech_mux2 i_9734(.S(\nbus_11289[8] ), .A(opc[14]), .B(n_9886), .Z(n_26684
		));
	notech_ao4 i_115151937(.A(n_55884), .B(n_33106), .C(n_333260960), .D(n_33105
		), .Z(n_200360392));
	notech_reg_set opc_reg_15(.CP(n_63506), .D(n_26690), .SD(1'b1), .Q(opc[
		15]));
	notech_mux2 i_9742(.S(\nbus_11289[8] ), .A(opc[15]), .B(n_9891), .Z(n_26690
		));
	notech_ao4 i_115551933(.A(n_61094), .B(n_30854), .C(n_57006), .D(n_31531
		), .Z(n_2002));
	notech_reg_set opc_reg_16(.CP(n_63506), .D(n_26696), .SD(1'b1), .Q(opc[
		16]));
	notech_mux2 i_9750(.S(n_31159), .A(opc[16]), .B(n_31143), .Z(n_26696));
	notech_nand2 i_115751931(.A(n_2000), .B(n_199960390), .Z(n_200160391));
	notech_reg_set opc_reg_17(.CP(n_63456), .D(n_26702), .SD(1'b1), .Q(opc[
		17]));
	notech_mux2 i_9758(.S(n_31159), .A(opc[17]), .B(n_31144), .Z(n_26702));
	notech_ao4 i_115451934(.A(n_331060938), .B(n_31499), .C(n_122826555), .D
		(n_33170), .Z(n_2000));
	notech_reg_set opc_reg_18(.CP(n_63456), .D(n_26708), .SD(1'b1), .Q(opc[
		18]));
	notech_mux2 i_9768(.S(n_31159), .A(opc[18]), .B(n_31145), .Z(n_26708));
	notech_ao4 i_115351935(.A(n_109226419), .B(n_122926556), .C(n_122626553)
		, .D(n_58902), .Z(n_199960390));
	notech_reg_set opc_reg_19(.CP(n_63456), .D(n_26714), .SD(1'b1), .Q(opc[
		19]));
	notech_mux2 i_9776(.S(n_31159), .A(opc[19]), .B(n_31146), .Z(n_26714));
	notech_reg_set opc_reg_20(.CP(n_63456), .D(n_26720), .SD(1'b1), .Q(opc[
		20]));
	notech_mux2 i_9784(.S(n_31159), .A(opc[20]), .B(n_31147), .Z(n_26720));
	notech_reg_set opc_reg_21(.CP(n_63456), .D(n_26726), .SD(1'b1), .Q(opc[
		21]));
	notech_mux2 i_9792(.S(n_31159), .A(opc[21]), .B(n_31148), .Z(n_26726));
	notech_reg_set opc_reg_22(.CP(n_63456), .D(n_26732), .SD(1'b1), .Q(opc[
		22]));
	notech_mux2 i_9800(.S(n_31159), .A(opc[22]), .B(n_31149), .Z(n_26732));
	notech_ao4 i_29652779(.A(n_57225), .B(n_31666), .C(n_57211), .D(n_31431)
		, .Z(n_1994));
	notech_reg_set opc_reg_23(.CP(n_63456), .D(n_26738), .SD(1'b1), .Q(opc[
		23]));
	notech_mux2 i_9809(.S(n_31159), .A(opc[23]), .B(n_31150), .Z(n_26738));
	notech_ao4 i_29552780(.A(n_59095), .B(n_31922), .C(n_58696), .D(n_31987)
		, .Z(n_1993));
	notech_reg_set opc_reg_24(.CP(n_63456), .D(n_26744), .SD(1'b1), .Q(opc[
		24]));
	notech_mux2 i_9817(.S(n_31159), .A(opc[24]), .B(n_31151), .Z(n_26744));
	notech_and2 i_29952776(.A(n_1990), .B(n_1989), .Z(n_1991));
	notech_reg_set opc_reg_25(.CP(n_63456), .D(n_26750), .SD(1'b1), .Q(opc[
		25]));
	notech_mux2 i_9825(.S(n_31159), .A(opc[25]), .B(n_31152), .Z(n_26750));
	notech_ao4 i_29452781(.A(n_31595), .B(n_57097), .C(n_57081), .D(n_31890)
		, .Z(n_1990));
	notech_reg_set opc_reg_26(.CP(n_63456), .D(n_26756), .SD(1'b1), .Q(opc[
		26]));
	notech_mux2 i_9833(.S(n_31159), .A(opc[26]), .B(n_31153), .Z(n_26756));
	notech_ao4 i_29352782(.A(n_57072), .B(n_31826), .C(n_57059), .D(n_31698)
		, .Z(n_1989));
	notech_reg_set opc_reg_27(.CP(n_63456), .D(n_26762), .SD(1'b1), .Q(opc[
		27]));
	notech_mux2 i_9841(.S(n_31159), .A(opc[27]), .B(n_31154), .Z(n_26762));
	notech_and4 i_30152774(.A(n_198695889), .B(n_198595890), .C(n_198395892)
		, .D(n_1982), .Z(n_198860388));
	notech_reg_set opc_reg_28(.CP(n_63456), .D(n_26768), .SD(1'b1), .Q(opc[
		28]));
	notech_mux2 i_9849(.S(n_31159), .A(opc[28]), .B(n_31155), .Z(n_26768));
	notech_reg_set opc_reg_29(.CP(n_63672), .D(n_26774), .SD(1'b1), .Q(opc[
		29]));
	notech_mux2 i_9857(.S(n_31159), .A(opc[29]), .B(n_31156), .Z(n_26774));
	notech_ao4 i_29252783(.A(n_57199), .B(n_31955), .C(n_57189), .D(n_31730)
		, .Z(n_198695889));
	notech_reg_set opc_reg_30(.CP(n_63378), .D(n_26780), .SD(1'b1), .Q(opc[
		30]));
	notech_mux2 i_9865(.S(n_31159), .A(opc[30]), .B(n_31157), .Z(n_26780));
	notech_ao4 i_29152784(.A(n_57178), .B(n_32019), .C(n_57163), .D(n_31858)
		, .Z(n_198595890));
	notech_reg_set opc_reg_31(.CP(n_63378), .D(n_26786), .SD(1'b1), .Q(opc[
		31]));
	notech_mux2 i_9873(.S(n_31159), .A(n_60602), .B(n_31158), .Z(n_26786));
	notech_reg nZF_reg(.CP(n_63378), .D(n_26792), .CD(n_62380), .Q(nZF));
	notech_mux2 i_9881(.S(n_16830), .A(nZF), .B(n_16833), .Z(n_26792));
	notech_ao4 i_29052785(.A(n_57152), .B(n_33112), .C(n_57136), .D(n_31762)
		, .Z(n_198395892));
	notech_reg regs_reg_0_0(.CP(n_63378), .D(n_26798), .CD(n_62380), .Q(regs_0
		[0]));
	notech_mux2 i_9889(.S(n_4456), .A(n_11566), .B(regs_0[0]), .Z(n_26798)
		);
	notech_ao4 i_28952786(.A(n_57609), .B(n_33111), .C(n_57112), .D(n_31794)
		, .Z(n_1982));
	notech_reg regs_reg_0_1(.CP(n_63378), .D(n_26804), .CD(n_62379), .Q(regs_0
		[1]));
	notech_mux2 i_9897(.S(n_4456), .A(n_30907), .B(regs_0[1]), .Z(n_26804)
		);
	notech_reg regs_reg_0_2(.CP(n_63378), .D(n_26810), .CD(n_62379), .Q(regs_0
		[2]));
	notech_mux2 i_9905(.S(n_4456), .A(n_30400), .B(regs_0[2]), .Z(n_26810)
		);
	notech_reg regs_reg_0_3(.CP(n_63378), .D(n_26816), .CD(n_62379), .Q(regs_0
		[3]));
	notech_mux2 i_9913(.S(n_4456), .A(n_4416), .B(regs_0[3]), .Z(n_26816));
	notech_reg regs_reg_0_4(.CP(n_63378), .D(n_26825), .CD(n_62378), .Q(regs_0
		[4]));
	notech_mux2 i_9921(.S(n_4456), .A(n_30399), .B(regs_0[4]), .Z(n_26825)
		);
	notech_ao4 i_22052855(.A(n_57097), .B(n_31597), .C(n_57225), .D(n_31668)
		, .Z(n_197895895));
	notech_reg regs_reg_0_5(.CP(n_63378), .D(n_26831), .CD(n_62378), .Q(regs_0
		[5]));
	notech_mux2 i_9929(.S(n_4456), .A(n_4377), .B(regs_0[5]), .Z(n_26831));
	notech_ao4 i_21952856(.A(n_57211), .B(n_31433), .C(n_59095), .D(n_31924)
		, .Z(n_197795896));
	notech_reg regs_reg_0_6(.CP(n_63476), .D(n_26837), .CD(n_62378), .Q(regs_0
		[6]));
	notech_mux2 i_9937(.S(n_4456), .A(n_11602), .B(regs_0[6]), .Z(n_26837)
		);
	notech_and2 i_22352852(.A(n_197595898), .B(n_197495899), .Z(n_197695897)
		);
	notech_reg regs_reg_0_7(.CP(n_63476), .D(n_26843), .CD(n_62378), .Q(regs_0
		[7]));
	notech_mux2 i_9945(.S(n_4456), .A(n_4376), .B(regs_0[7]), .Z(n_26843));
	notech_ao4 i_21852857(.A(n_58696), .B(n_31989), .C(n_57081), .D(n_31892)
		, .Z(n_197595898));
	notech_reg regs_reg_0_8(.CP(n_63476), .D(n_26849), .CD(n_62378), .Q(regs_0
		[8]));
	notech_mux2 i_9953(.S(n_4456), .A(n_11614), .B(regs_0[8]), .Z(n_26849)
		);
	notech_ao4 i_21752858(.A(n_57072), .B(n_31828), .C(n_57059), .D(n_31700)
		, .Z(n_197495899));
	notech_reg regs_reg_0_9(.CP(n_63476), .D(n_26855), .CD(n_62379), .Q(regs_0
		[9]));
	notech_mux2 i_9961(.S(n_4456), .A(n_30392), .B(regs_0[9]), .Z(n_26855)
		);
	notech_and4 i_22552850(.A(n_197195902), .B(n_197095903), .C(n_196895905)
		, .D(n_1967), .Z(n_197395900));
	notech_reg regs_reg_0_10(.CP(n_63476), .D(n_26861), .CD(n_62379), .Q(regs_0
		[10]));
	notech_mux2 i_9969(.S(n_4456), .A(n_30643), .B(regs_0[10]), .Z(n_26861)
		);
	notech_reg regs_reg_0_11(.CP(n_63476), .D(n_26867), .CD(n_62379), .Q(regs_0
		[11]));
	notech_mux2 i_9977(.S(n_4456), .A(n_441467998), .B(regs_0[11]), .Z(n_26867
		));
	notech_ao4 i_21652859(.A(n_57199), .B(n_31957), .C(n_57189), .D(n_31732)
		, .Z(n_197195902));
	notech_reg regs_reg_0_12(.CP(n_63476), .D(n_26873), .CD(n_62379), .Q(regs_0
		[12]));
	notech_mux2 i_9985(.S(n_4456), .A(n_441367997), .B(regs_0[12]), .Z(n_26873
		));
	notech_ao4 i_21552860(.A(n_57178), .B(n_32021), .C(n_57163), .D(n_31860)
		, .Z(n_197095903));
	notech_reg regs_reg_0_13(.CP(n_63476), .D(n_26879), .CD(n_62356), .Q(regs_0
		[13]));
	notech_mux2 i_9993(.S(n_4456), .A(n_11644), .B(regs_0[13]), .Z(n_26879)
		);
	notech_reg regs_reg_0_14(.CP(n_63476), .D(n_26885), .CD(n_62356), .Q(regs_0
		[14]));
	notech_mux2 i_10001(.S(n_4456), .A(n_11650), .B(regs_0[14]), .Z(n_26885)
		);
	notech_ao4 i_21452861(.A(n_57152), .B(n_33116), .C(n_57136), .D(n_31764)
		, .Z(n_196895905));
	notech_reg regs_reg_0_15(.CP(n_63476), .D(n_26891), .CD(n_62356), .Q(regs_0
		[15]));
	notech_mux2 i_10009(.S(n_4456), .A(n_441267996), .B(regs_0[15]), .Z(n_26891
		));
	notech_ao4 i_21352862(.A(n_57609), .B(n_33115), .C(n_57112), .D(n_31796)
		, .Z(n_1967));
	notech_reg regs_reg_0_16(.CP(n_63476), .D(n_26897), .CD(n_62356), .Q(regs_0
		[16]));
	notech_mux2 i_10017(.S(n_56041), .A(n_31161), .B(regs_0[16]), .Z(n_26897
		));
	notech_reg regs_reg_0_17(.CP(n_63476), .D(n_26903), .CD(n_62356), .Q(regs_0
		[17]));
	notech_mux2 i_10025(.S(n_56041), .A(n_11668), .B(regs_0[17]), .Z(n_26903
		));
	notech_reg regs_reg_0_18(.CP(n_63476), .D(n_26909), .CD(n_62356), .Q(regs_0
		[18]));
	notech_mux2 i_10033(.S(n_56041), .A(n_31162), .B(regs_0[18]), .Z(n_26909
		));
	notech_ao4 i_17152904(.A(n_57225), .B(n_31667), .C(n_57211), .D(n_31432)
		, .Z(n_196395907));
	notech_reg regs_reg_0_19(.CP(n_63476), .D(n_26915), .CD(n_62356), .Q(regs_0
		[19]));
	notech_mux2 i_10041(.S(n_56041), .A(n_31163), .B(regs_0[19]), .Z(n_26915
		));
	notech_ao4 i_17052905(.A(n_59095), .B(n_31923), .C(n_58696), .D(n_31988)
		, .Z(n_196295908));
	notech_reg regs_reg_0_20(.CP(n_63476), .D(n_26921), .CD(n_62356), .Q(regs_0
		[20]));
	notech_mux2 i_10049(.S(n_56041), .A(n_31164), .B(regs_0[20]), .Z(n_26921
		));
	notech_and2 i_17452901(.A(n_196095910), .B(n_1958), .Z(n_196195909));
	notech_reg regs_reg_0_21(.CP(n_63476), .D(n_26927), .CD(n_62356), .Q(regs_0
		[21]));
	notech_mux2 i_10057(.S(n_56041), .A(n_3042), .B(regs_0[21]), .Z(n_26927)
		);
	notech_ao4 i_16952906(.A(n_57097), .B(n_31596), .C(n_57086), .D(n_31891)
		, .Z(n_196095910));
	notech_reg regs_reg_0_22(.CP(n_63476), .D(n_26933), .CD(n_62354), .Q(regs_0
		[22]));
	notech_mux2 i_10065(.S(n_56041), .A(n_31165), .B(regs_0[22]), .Z(n_26933
		));
	notech_ao4 i_16852907(.A(n_57068), .B(n_31827), .C(n_57059), .D(n_31699)
		, .Z(n_1958));
	notech_reg regs_reg_0_23(.CP(n_63476), .D(n_26941), .CD(n_62354), .Q(regs_0
		[23]));
	notech_mux2 i_10074(.S(n_56041), .A(n_11704), .B(regs_0[23]), .Z(n_26941
		));
	notech_and4 i_17652899(.A(n_195595912), .B(n_195495913), .C(n_195295915)
		, .D(n_1951), .Z(n_1957));
	notech_reg regs_reg_0_24(.CP(n_63476), .D(n_26948), .CD(n_62354), .Q(regs_0
		[24]));
	notech_mux2 i_10082(.S(n_56041), .A(n_31166), .B(regs_0[24]), .Z(n_26948
		));
	notech_reg regs_reg_0_25(.CP(n_63474), .D(n_26956), .CD(n_62354), .Q(regs_0
		[25]));
	notech_mux2 i_10090(.S(n_56041), .A(n_11716), .B(regs_0[25]), .Z(n_26956
		));
	notech_ao4 i_16752908(.A(n_57199), .B(n_31956), .C(n_57189), .D(n_31731)
		, .Z(n_195595912));
	notech_reg regs_reg_0_26(.CP(n_63474), .D(n_26963), .CD(n_62354), .Q(regs_0
		[26]));
	notech_mux2 i_10098(.S(n_56041), .A(n_31167), .B(regs_0[26]), .Z(n_26963
		));
	notech_ao4 i_16652909(.A(n_57178), .B(n_32020), .C(n_57163), .D(n_31859)
		, .Z(n_195495913));
	notech_reg regs_reg_0_27(.CP(n_63546), .D(n_26969), .CD(n_62354), .Q(regs_0
		[27]));
	notech_mux2 i_10106(.S(n_56041), .A(n_31168), .B(regs_0[27]), .Z(n_26969
		));
	notech_reg regs_reg_0_28(.CP(n_63546), .D(n_26975), .CD(n_62354), .Q(regs_0
		[28]));
	notech_mux2 i_10114(.S(n_56041), .A(n_31169), .B(regs_0[28]), .Z(n_26975
		));
	notech_ao4 i_16552910(.A(n_57152), .B(n_33114), .C(n_57136), .D(n_31763)
		, .Z(n_195295915));
	notech_reg regs_reg_0_29(.CP(n_63546), .D(n_26982), .CD(n_62354), .Q(regs_0
		[29]));
	notech_mux2 i_10122(.S(n_56041), .A(n_30407), .B(regs_0[29]), .Z(n_26982
		));
	notech_ao4 i_16452911(.A(n_57609), .B(n_33113), .C(n_57112), .D(n_31795)
		, .Z(n_1951));
	notech_reg regs_reg_0_30(.CP(n_63546), .D(n_26989), .CD(n_62354), .Q(regs_0
		[30]));
	notech_mux2 i_10130(.S(n_56041), .A(n_31170), .B(regs_0[30]), .Z(n_26989
		));
	notech_nand3 i_2621784(.A(n_194995916), .B(n_2029), .C(n_193795917), .Z(n_1950
		));
	notech_reg regs_reg_0_31(.CP(n_63546), .D(n_26995), .CD(n_62354), .Q(regs_0
		[31]));
	notech_mux2 i_10138(.S(n_56041), .A(n_31171), .B(regs_0[31]), .Z(n_26995
		));
	notech_nao3 i_158151509(.A(n_63776), .B(opc_10[25]), .C(n_337961007), .Z
		(n_194995916));
	notech_reg cr1_reg_0(.CP(n_63546), .D(n_27001), .CD(n_62357), .Q(nbus_14541
		[0]));
	notech_mux2 i_10146(.S(n_98090347), .A(opa[0]), .B(nbus_14541[0]), .Z(n_27001
		));
	notech_nand2 i_157951511(.A(sav_esp[25]), .B(n_61864), .Z(n_1948));
	notech_reg cr1_reg_1(.CP(n_63546), .D(n_27007), .CD(n_62357), .Q(nbus_14541
		[1]));
	notech_mux2 i_10154(.S(n_98090347), .A(opa[1]), .B(nbus_14541[1]), .Z(n_27007
		));
	notech_reg cr1_reg_2(.CP(n_63546), .D(n_27013), .CD(n_62357), .Q(nbus_14541
		[2]));
	notech_mux2 i_10162(.S(n_98090347), .A(opa[2]), .B(nbus_14541[2]), .Z(n_27013
		));
	notech_reg cr1_reg_3(.CP(n_63546), .D(n_27019), .CD(n_62357), .Q(nbus_14541
		[3]));
	notech_mux2 i_10170(.S(n_98090347), .A(opa[3]), .B(nbus_14541[3]), .Z(n_27019
		));
	notech_reg cr1_reg_4(.CP(n_63546), .D(n_27025), .CD(n_62357), .Q(nbus_14541
		[4]));
	notech_mux2 i_10178(.S(n_98090347), .A(opa[4]), .B(nbus_14541[4]), .Z(n_27025
		));
	notech_reg cr1_reg_5(.CP(n_63546), .D(n_27031), .CD(n_62358), .Q(nbus_14541
		[5]));
	notech_mux2 i_10186(.S(n_98090347), .A(opa[5]), .B(nbus_14541[5]), .Z(n_27031
		));
	notech_reg cr1_reg_6(.CP(n_63546), .D(n_27037), .CD(n_62358), .Q(nbus_14541
		[6]));
	notech_mux2 i_10194(.S(n_98090347), .A(opa[6]), .B(nbus_14541[6]), .Z(n_27037
		));
	notech_reg cr1_reg_7(.CP(n_63546), .D(n_27043), .CD(n_62358), .Q(nbus_14541
		[7]));
	notech_mux2 i_10202(.S(n_98090347), .A(opa[7]), .B(nbus_14541[7]), .Z(n_27043
		));
	notech_reg cr1_reg_8(.CP(n_63546), .D(n_27049), .CD(n_62358), .Q(nbus_14541
		[8]));
	notech_mux2 i_10210(.S(n_98090347), .A(opa[8]), .B(nbus_14541[8]), .Z(n_27049
		));
	notech_reg cr1_reg_9(.CP(n_63546), .D(n_27055), .CD(n_62357), .Q(nbus_14541
		[9]));
	notech_mux2 i_10218(.S(n_98090347), .A(opa[9]), .B(nbus_14541[9]), .Z(n_27055
		));
	notech_reg cr1_reg_10(.CP(n_63546), .D(n_27061), .CD(n_62356), .Q(nbus_14541
		[10]));
	notech_mux2 i_10226(.S(n_98090347), .A(opa[10]), .B(nbus_14541[10]), .Z(n_27061
		));
	notech_reg cr1_reg_11(.CP(n_63546), .D(n_27067), .CD(n_62357), .Q(nbus_14541
		[11]));
	notech_mux2 i_10234(.S(n_98090347), .A(opa[11]), .B(nbus_14541[11]), .Z(n_27067
		));
	notech_or2 i_158051510(.A(n_126226589), .B(n_363350926), .Z(n_193795917)
		);
	notech_reg cr1_reg_12(.CP(n_63546), .D(n_27073), .CD(n_62356), .Q(nbus_14541
		[12]));
	notech_mux2 i_10242(.S(n_98090347), .A(opa[12]), .B(nbus_14541[12]), .Z(n_27073
		));
	notech_or4 i_2521527(.A(n_2017), .B(n_201260397), .C(n_1935), .D(n_1924)
		, .Z(n_1936));
	notech_reg cr1_reg_13(.CP(n_63474), .D(n_27079), .CD(n_62356), .Q(nbus_14541
		[13]));
	notech_mux2 i_10250(.S(n_98090347), .A(opa[13]), .B(nbus_14541[13]), .Z(n_27079
		));
	notech_ao3 i_136951721(.A(n_63776), .B(opc_10[24]), .C(n_337661004), .Z(n_1935
		));
	notech_reg cr1_reg_14(.CP(n_63474), .D(n_27087), .CD(n_62357), .Q(nbus_14541
		[14]));
	notech_mux2 i_10258(.S(n_98090347), .A(opa[14]), .B(nbus_14541[14]), .Z(n_27087
		));
	notech_reg cr1_reg_15(.CP(n_63474), .D(n_27098), .CD(n_62357), .Q(nbus_14541
		[15]));
	notech_mux2 i_10266(.S(n_98090347), .A(opa[15]), .B(nbus_14541[15]), .Z(n_27098
		));
	notech_reg cr1_reg_16(.CP(n_63474), .D(n_27104), .CD(n_62357), .Q(nbus_14541
		[16]));
	notech_mux2 i_10274(.S(n_56063), .A(opa[16]), .B(nbus_14541[16]), .Z(n_27104
		));
	notech_reg cr1_reg_17(.CP(n_63474), .D(n_27110), .CD(n_62357), .Q(nbus_14541
		[17]));
	notech_mux2 i_10286(.S(n_56063), .A(opa[17]), .B(nbus_14541[17]), .Z(n_27110
		));
	notech_reg cr1_reg_18(.CP(n_63474), .D(n_27116), .CD(n_62357), .Q(nbus_14541
		[18]));
	notech_mux2 i_10295(.S(n_56063), .A(opa[18]), .B(nbus_14541[18]), .Z(n_27116
		));
	notech_reg cr1_reg_19(.CP(n_63474), .D(n_27122), .CD(n_62352), .Q(nbus_14541
		[19]));
	notech_mux2 i_10303(.S(n_56063), .A(opa[19]), .B(nbus_14541[19]), .Z(n_27122
		));
	notech_reg cr1_reg_20(.CP(n_63474), .D(n_27128), .CD(n_62352), .Q(nbus_14541
		[20]));
	notech_mux2 i_10311(.S(n_56063), .A(opa[20]), .B(nbus_14541[20]), .Z(n_27128
		));
	notech_reg cr1_reg_21(.CP(n_63474), .D(n_27134), .CD(n_62351), .Q(nbus_14541
		[21]));
	notech_mux2 i_10320(.S(n_56063), .A(opa[21]), .B(nbus_14541[21]), .Z(n_27134
		));
	notech_reg cr1_reg_22(.CP(n_63546), .D(n_27140), .CD(n_62351), .Q(nbus_14541
		[22]));
	notech_mux2 i_10328(.S(n_56063), .A(opa[22]), .B(nbus_14541[22]), .Z(n_27140
		));
	notech_reg cr1_reg_23(.CP(n_63472), .D(n_27146), .CD(n_62352), .Q(nbus_14541
		[23]));
	notech_mux2 i_10336(.S(n_56063), .A(opa[23]), .B(nbus_14541[23]), .Z(n_27146
		));
	notech_reg cr1_reg_24(.CP(n_63472), .D(n_27152), .CD(n_62352), .Q(nbus_14541
		[24]));
	notech_mux2 i_10344(.S(n_56063), .A(opa[24]), .B(nbus_14541[24]), .Z(n_27152
		));
	notech_nor2 i_136851722(.A(n_124126568), .B(n_364628688), .Z(n_1924));
	notech_reg cr1_reg_25(.CP(n_63542), .D(n_27158), .CD(n_62352), .Q(nbus_14541
		[25]));
	notech_mux2 i_10352(.S(n_56063), .A(opa[25]), .B(nbus_14541[25]), .Z(n_27158
		));
	notech_or4 i_2421334(.A(n_200660395), .B(n_200160391), .C(n_1922), .D(n_1911
		), .Z(n_1923));
	notech_reg cr1_reg_26(.CP(n_63542), .D(n_27164), .CD(n_62352), .Q(nbus_14541
		[26]));
	notech_mux2 i_10360(.S(n_56063), .A(opa[26]), .B(nbus_14541[26]), .Z(n_27164
		));
	notech_ao3 i_115051938(.A(n_63776), .B(opc_10[23]), .C(n_337461002), .Z(n_1922
		));
	notech_reg cr1_reg_27(.CP(n_63542), .D(n_27170), .CD(n_62352), .Q(nbus_14541
		[27]));
	notech_mux2 i_10368(.S(n_56063), .A(opa[27]), .B(nbus_14541[27]), .Z(n_27170
		));
	notech_reg cr1_reg_28(.CP(n_63542), .D(n_27176), .CD(n_62351), .Q(nbus_14541
		[28]));
	notech_mux2 i_10376(.S(n_56063), .A(opa[28]), .B(nbus_14541[28]), .Z(n_27176
		));
	notech_reg cr1_reg_29(.CP(n_63542), .D(n_27182), .CD(n_62351), .Q(nbus_14541
		[29]));
	notech_mux2 i_10384(.S(n_56063), .A(opa[29]), .B(nbus_14541[29]), .Z(n_27182
		));
	notech_reg cr1_reg_30(.CP(n_63542), .D(n_27188), .CD(n_62351), .Q(nbus_14541
		[30]));
	notech_mux2 i_10393(.S(n_56063), .A(opa[30]), .B(nbus_14541[30]), .Z(n_27188
		));
	notech_reg cr1_reg_31(.CP(n_63542), .D(n_27194), .CD(n_62351), .Q(nbus_14541
		[31]));
	notech_mux2 i_10401(.S(n_56063), .A(opa[31]), .B(nbus_14541[31]), .Z(n_27194
		));
	notech_reg cr2_reg_reg_0(.CP(n_63542), .D(n_27203), .CD(n_62351), .Q(cr2_reg
		[0]));
	notech_mux2 i_10409(.S(\nbus_11278[0] ), .A(cr2_reg[0]), .B(n_8107), .Z(n_27203
		));
	notech_reg cr2_reg_reg_1(.CP(n_63542), .D(n_27209), .CD(n_62351), .Q(cr2_reg
		[1]));
	notech_mux2 i_10417(.S(\nbus_11278[0] ), .A(cr2_reg[1]), .B(n_8113), .Z(n_27209
		));
	notech_reg cr2_reg_reg_2(.CP(n_63626), .D(n_27215), .CD(n_62351), .Q(cr2_reg
		[2]));
	notech_mux2 i_10425(.S(\nbus_11278[0] ), .A(cr2_reg[2]), .B(n_8119), .Z(n_27215
		));
	notech_reg cr2_reg_reg_3(.CP(n_63626), .D(n_27221), .CD(n_62351), .Q(cr2_reg
		[3]));
	notech_mux2 i_10433(.S(\nbus_11278[0] ), .A(cr2_reg[3]), .B(n_8125), .Z(n_27221
		));
	notech_reg cr2_reg_reg_4(.CP(n_63626), .D(n_27227), .CD(n_62351), .Q(cr2_reg
		[4]));
	notech_mux2 i_10441(.S(\nbus_11278[0] ), .A(cr2_reg[4]), .B(n_8131), .Z(n_27227
		));
	notech_reg cr2_reg_reg_5(.CP(n_63626), .D(n_27233), .CD(n_62351), .Q(cr2_reg
		[5]));
	notech_mux2 i_10449(.S(\nbus_11278[0] ), .A(cr2_reg[5]), .B(n_8137), .Z(n_27233
		));
	notech_nor2 i_114951939(.A(n_122226549), .B(n_363450925), .Z(n_1911));
	notech_reg cr2_reg_reg_6(.CP(n_63626), .D(n_27239), .CD(n_62353), .Q(cr2_reg
		[6]));
	notech_mux2 i_10457(.S(\nbus_11278[0] ), .A(cr2_reg[6]), .B(n_8143), .Z(n_27239
		));
	notech_reg cr2_reg_reg_7(.CP(n_63626), .D(n_27245), .CD(n_62353), .Q(cr2_reg
		[7]));
	notech_mux2 i_10465(.S(\nbus_11278[0] ), .A(cr2_reg[7]), .B(n_8149), .Z(n_27245
		));
	notech_reg cr2_reg_reg_8(.CP(n_63626), .D(n_27251), .CD(n_62353), .Q(cr2_reg
		[8]));
	notech_mux2 i_10473(.S(\nbus_11278[0] ), .A(cr2_reg[8]), .B(n_8155), .Z(n_27251
		));
	notech_reg cr2_reg_reg_9(.CP(n_63626), .D(n_27257), .CD(n_62353), .Q(cr2_reg
		[9]));
	notech_mux2 i_10481(.S(\nbus_11278[0] ), .A(cr2_reg[9]), .B(n_8161), .Z(n_27257
		));
	notech_reg cr2_reg_reg_10(.CP(n_63626), .D(n_27263), .CD(n_62353), .Q(cr2_reg
		[10]));
	notech_mux2 i_10489(.S(\nbus_11278[0] ), .A(cr2_reg[10]), .B(n_8167), .Z
		(n_27263));
	notech_reg cr2_reg_reg_11(.CP(n_63626), .D(n_27269), .CD(n_62354), .Q(cr2_reg
		[11]));
	notech_mux2 i_10497(.S(\nbus_11278[0] ), .A(cr2_reg[11]), .B(n_8173), .Z
		(n_27269));
	notech_reg cr2_reg_reg_12(.CP(n_63626), .D(n_27275), .CD(n_62354), .Q(cr2_reg
		[12]));
	notech_mux2 i_10505(.S(\nbus_11278[0] ), .A(cr2_reg[12]), .B(n_8179), .Z
		(n_27275));
	notech_reg cr2_reg_reg_13(.CP(n_63626), .D(n_27281), .CD(n_62353), .Q(cr2_reg
		[13]));
	notech_mux2 i_10513(.S(\nbus_11278[0] ), .A(cr2_reg[13]), .B(n_8185), .Z
		(n_27281));
	notech_reg cr2_reg_reg_14(.CP(n_63626), .D(n_27287), .CD(n_62353), .Q(cr2_reg
		[14]));
	notech_mux2 i_10521(.S(\nbus_11278[0] ), .A(cr2_reg[14]), .B(n_8191), .Z
		(n_27287));
	notech_reg cr2_reg_reg_15(.CP(n_63626), .D(n_27293), .CD(n_62353), .Q(cr2_reg
		[15]));
	notech_mux2 i_10529(.S(\nbus_11278[0] ), .A(cr2_reg[15]), .B(n_8197), .Z
		(n_27293));
	notech_reg cr2_reg_reg_16(.CP(n_63626), .D(n_27299), .CD(n_62352), .Q(cr2_reg
		[16]));
	notech_mux2 i_10537(.S(\nbus_11278[0] ), .A(cr2_reg[16]), .B(n_8203), .Z
		(n_27299));
	notech_reg cr2_reg_reg_17(.CP(n_63626), .D(n_27305), .CD(n_62352), .Q(cr2_reg
		[17]));
	notech_mux2 i_10545(.S(\nbus_11278[0] ), .A(cr2_reg[17]), .B(n_8209), .Z
		(n_27305));
	notech_reg cr2_reg_reg_18(.CP(n_63626), .D(n_27311), .CD(n_62352), .Q(cr2_reg
		[18]));
	notech_mux2 i_10553(.S(n_55811), .A(cr2_reg[18]), .B(n_8215), .Z(n_27311
		));
	notech_reg cr2_reg_reg_19(.CP(n_63626), .D(n_27317), .CD(n_62352), .Q(cr2_reg
		[19]));
	notech_mux2 i_10561(.S(n_55811), .A(cr2_reg[19]), .B(n_8221), .Z(n_27317
		));
	notech_reg cr2_reg_reg_20(.CP(n_63542), .D(n_27323), .CD(n_62352), .Q(cr2_reg
		[20]));
	notech_mux2 i_10569(.S(n_55811), .A(cr2_reg[20]), .B(n_8227), .Z(n_27323
		));
	notech_reg cr2_reg_reg_21(.CP(n_63626), .D(n_27329), .CD(n_62353), .Q(cr2_reg
		[21]));
	notech_mux2 i_10577(.S(n_55811), .A(cr2_reg[21]), .B(n_8233), .Z(n_27329
		));
	notech_reg cr2_reg_reg_22(.CP(n_63544), .D(n_27335), .CD(n_62353), .Q(cr2_reg
		[22]));
	notech_mux2 i_10585(.S(n_55811), .A(cr2_reg[22]), .B(n_8239), .Z(n_27335
		));
	notech_reg cr2_reg_reg_23(.CP(n_63544), .D(n_27341), .CD(n_62353), .Q(cr2_reg
		[23]));
	notech_mux2 i_10593(.S(n_55811), .A(cr2_reg[23]), .B(n_8245), .Z(n_27341
		));
	notech_reg cr2_reg_reg_24(.CP(n_63544), .D(n_27347), .CD(n_62353), .Q(cr2_reg
		[24]));
	notech_mux2 i_10601(.S(n_55811), .A(cr2_reg[24]), .B(n_8251), .Z(n_27347
		));
	notech_reg cr2_reg_reg_25(.CP(n_63544), .D(n_27353), .CD(n_62364), .Q(cr2_reg
		[25]));
	notech_mux2 i_10609(.S(n_55811), .A(cr2_reg[25]), .B(n_8257), .Z(n_27353
		));
	notech_reg cr2_reg_reg_26(.CP(n_63544), .D(n_27359), .CD(n_62364), .Q(cr2_reg
		[26]));
	notech_mux2 i_10617(.S(n_55811), .A(cr2_reg[26]), .B(n_8263), .Z(n_27359
		));
	notech_reg cr2_reg_reg_27(.CP(n_63544), .D(n_27365), .CD(n_62364), .Q(cr2_reg
		[27]));
	notech_mux2 i_10625(.S(n_55811), .A(cr2_reg[27]), .B(n_8269), .Z(n_27365
		));
	notech_reg cr2_reg_reg_28(.CP(n_63544), .D(n_27372), .CD(n_62364), .Q(cr2_reg
		[28]));
	notech_mux2 i_10633(.S(n_55811), .A(cr2_reg[28]), .B(n_8275), .Z(n_27372
		));
	notech_reg cr2_reg_reg_29(.CP(n_63544), .D(n_27381), .CD(n_62364), .Q(cr2_reg
		[29]));
	notech_mux2 i_10641(.S(n_55811), .A(cr2_reg[29]), .B(n_8281), .Z(n_27381
		));
	notech_reg cr2_reg_reg_30(.CP(n_63544), .D(n_27387), .CD(n_62364), .Q(cr2_reg
		[30]));
	notech_mux2 i_10649(.S(n_55811), .A(cr2_reg[30]), .B(n_8287), .Z(n_27387
		));
	notech_reg cr2_reg_reg_31(.CP(n_63544), .D(n_27393), .CD(n_62365), .Q(cr2_reg
		[31]));
	notech_mux2 i_10657(.S(n_55811), .A(cr2_reg[31]), .B(n_8293), .Z(n_27393
		));
	notech_reg cr3_reg_0(.CP(n_63544), .D(n_27399), .CD(n_62364), .Q(\nbus_14540[0] 
		));
	notech_mux2 i_10665(.S(n_98190348), .A(opa[0]), .B(\nbus_14540[0] ), .Z(n_27399
		));
	notech_reg cr3_reg_1(.CP(n_63544), .D(n_27405), .CD(n_62364), .Q(\nbus_14540[1] 
		));
	notech_mux2 i_10673(.S(n_98190348), .A(opa[1]), .B(\nbus_14540[1] ), .Z(n_27405
		));
	notech_reg cr3_reg_2(.CP(n_63544), .D(n_27411), .CD(n_62364), .Q(\nbus_14540[2] 
		));
	notech_mux2 i_10681(.S(n_98190348), .A(opa[2]), .B(\nbus_14540[2] ), .Z(n_27411
		));
	notech_reg cr3_reg_3(.CP(n_63544), .D(n_27417), .CD(n_62363), .Q(\nbus_14540[3] 
		));
	notech_mux2 i_10689(.S(n_98190348), .A(opa[3]), .B(\nbus_14540[3] ), .Z(n_27417
		));
	notech_reg cr3_reg_4(.CP(n_63544), .D(n_27423), .CD(n_62363), .Q(\nbus_14540[4] 
		));
	notech_mux2 i_10697(.S(n_98190348), .A(opa[4]), .B(\nbus_14540[4] ), .Z(n_27423
		));
	notech_reg cr3_reg_5(.CP(n_63544), .D(n_27429), .CD(n_62363), .Q(\nbus_14540[5] 
		));
	notech_mux2 i_10705(.S(n_98190348), .A(opa[5]), .B(\nbus_14540[5] ), .Z(n_27429
		));
	notech_reg cr3_reg_6(.CP(n_63544), .D(n_27435), .CD(n_62363), .Q(\nbus_14540[6] 
		));
	notech_mux2 i_10715(.S(n_98190348), .A(opa[6]), .B(\nbus_14540[6] ), .Z(n_27435
		));
	notech_reg cr3_reg_7(.CP(n_63544), .D(n_27441), .CD(n_62363), .Q(\nbus_14540[7] 
		));
	notech_mux2 i_10723(.S(n_98190348), .A(opa[7]), .B(\nbus_14540[7] ), .Z(n_27441
		));
	notech_reg cr3_reg_8(.CP(n_63544), .D(n_27447), .CD(n_62364), .Q(\nbus_14540[8] 
		));
	notech_mux2 i_10731(.S(n_98190348), .A(opa[8]), .B(\nbus_14540[8] ), .Z(n_27447
		));
	notech_reg cr3_reg_9(.CP(n_63472), .D(n_27453), .CD(n_62364), .Q(\nbus_14540[9] 
		));
	notech_mux2 i_10739(.S(n_98190348), .A(opa[9]), .B(\nbus_14540[9] ), .Z(n_27453
		));
	notech_reg cr3_reg_10(.CP(n_63472), .D(n_27459), .CD(n_62363), .Q(\nbus_14540[10] 
		));
	notech_mux2 i_10747(.S(n_98190348), .A(opa[10]), .B(\nbus_14540[10] ), .Z
		(n_27459));
	notech_reg cr3_reg_11(.CP(n_63472), .D(n_27465), .CD(n_62364), .Q(\nbus_14540[11] 
		));
	notech_mux2 i_10755(.S(n_98190348), .A(opa[11]), .B(\nbus_14540[11] ), .Z
		(n_27465));
	notech_reg cr3_reg_12(.CP(n_63472), .D(n_27471), .CD(n_62367), .Q(cr3[12
		]));
	notech_mux2 i_10763(.S(n_98190348), .A(opa[12]), .B(cr3[12]), .Z(n_27471
		));
	notech_reg cr3_reg_13(.CP(n_63472), .D(n_27477), .CD(n_62367), .Q(cr3[13
		]));
	notech_mux2 i_10771(.S(n_98190348), .A(opa[13]), .B(cr3[13]), .Z(n_27477
		));
	notech_reg cr3_reg_14(.CP(n_63472), .D(n_27483), .CD(n_62365), .Q(cr3[14
		]));
	notech_mux2 i_10779(.S(n_98190348), .A(opa[14]), .B(cr3[14]), .Z(n_27483
		));
	notech_reg cr3_reg_15(.CP(n_63472), .D(n_27489), .CD(n_62367), .Q(cr3[15
		]));
	notech_mux2 i_10787(.S(n_98190348), .A(n_61034), .B(cr3[15]), .Z(n_27489
		));
	notech_reg cr3_reg_16(.CP(n_63472), .D(n_27495), .CD(n_62367), .Q(cr3[16
		]));
	notech_mux2 i_10795(.S(n_56936), .A(opa[16]), .B(cr3[16]), .Z(n_27495)
		);
	notech_reg cr3_reg_17(.CP(n_63472), .D(n_27506), .CD(n_62367), .Q(cr3[17
		]));
	notech_mux2 i_10803(.S(n_56936), .A(opa[17]), .B(cr3[17]), .Z(n_27506)
		);
	notech_reg cr3_reg_18(.CP(n_63542), .D(n_27516), .CD(n_62367), .Q(cr3[18
		]));
	notech_mux2 i_10811(.S(n_56936), .A(opa[18]), .B(cr3[18]), .Z(n_27516)
		);
	notech_reg cr3_reg_19(.CP(n_63536), .D(n_27522), .CD(n_62367), .Q(cr3[19
		]));
	notech_mux2 i_10819(.S(n_56936), .A(opa[19]), .B(cr3[19]), .Z(n_27522)
		);
	notech_reg cr3_reg_20(.CP(n_63470), .D(n_27528), .CD(n_62367), .Q(cr3[20
		]));
	notech_mux2 i_10827(.S(n_56936), .A(opa[20]), .B(cr3[20]), .Z(n_27528)
		);
	notech_reg cr3_reg_21(.CP(n_63536), .D(n_27535), .CD(n_62365), .Q(cr3[21
		]));
	notech_mux2 i_10835(.S(n_56936), .A(opa[21]), .B(cr3[21]), .Z(n_27535)
		);
	notech_reg cr3_reg_22(.CP(n_63536), .D(n_27541), .CD(n_62365), .Q(cr3[22
		]));
	notech_mux2 i_10843(.S(n_56936), .A(opa[22]), .B(cr3[22]), .Z(n_27541)
		);
	notech_ao4 i_185354144(.A(n_184660383), .B(n_32266), .C(n_60188), .D(n_323660864
		), .Z(n_1862));
	notech_reg cr3_reg_23(.CP(n_63536), .D(n_27547), .CD(n_62365), .Q(cr3[23
		]));
	notech_mux2 i_10851(.S(n_56936), .A(opa[23]), .B(cr3[23]), .Z(n_27547)
		);
	notech_reg cr3_reg_24(.CP(n_63536), .D(n_27553), .CD(n_62365), .Q(cr3[24
		]));
	notech_mux2 i_10859(.S(n_56936), .A(opa[24]), .B(cr3[24]), .Z(n_27553)
		);
	notech_reg cr3_reg_25(.CP(n_63536), .D(n_27559), .CD(n_62365), .Q(cr3[25
		]));
	notech_mux2 i_10867(.S(n_56936), .A(opa[25]), .B(cr3[25]), .Z(n_27559)
		);
	notech_reg cr3_reg_26(.CP(n_63536), .D(n_27565), .CD(n_62365), .Q(cr3[26
		]));
	notech_mux2 i_10875(.S(n_56936), .A(opa[26]), .B(cr3[26]), .Z(n_27565)
		);
	notech_reg cr3_reg_27(.CP(n_63536), .D(n_27571), .CD(n_62365), .Q(cr3[27
		]));
	notech_mux2 i_10883(.S(n_56936), .A(opa[27]), .B(cr3[27]), .Z(n_27571)
		);
	notech_ao4 i_98854995(.A(n_63748), .B(n_61958), .C(n_61056), .D(n_55831)
		, .Z(n_184660383));
	notech_reg cr3_reg_28(.CP(n_63536), .D(n_27577), .CD(n_62365), .Q(cr3[28
		]));
	notech_mux2 i_10891(.S(n_56936), .A(opa[28]), .B(cr3[28]), .Z(n_27577)
		);
	notech_reg cr3_reg_29(.CP(n_63536), .D(n_27583), .CD(n_62365), .Q(cr3[29
		]));
	notech_mux2 i_10899(.S(n_56936), .A(opa[29]), .B(cr3[29]), .Z(n_27583)
		);
	notech_or4 i_5455872(.A(n_61819), .B(n_57535), .C(n_57662), .D(n_32220),
		 .Z(n_184360381));
	notech_reg cr3_reg_30(.CP(n_63622), .D(n_27591), .CD(n_62365), .Q(cr3[30
		]));
	notech_mux2 i_10907(.S(n_56936), .A(opa[30]), .B(cr3[30]), .Z(n_27591)
		);
	notech_or4 i_29018(.A(n_32628), .B(n_32394), .C(n_61056), .D(n_57656), .Z
		(n_30380));
	notech_reg cr3_reg_31(.CP(n_63622), .D(n_27597), .CD(n_62359), .Q(cr3[31
		]));
	notech_mux2 i_10915(.S(n_56936), .A(opa[31]), .B(cr3[31]), .Z(n_27597)
		);
	notech_reg opa_reg_0(.CP(n_63622), .D(n_27603), .CD(n_62359), .Q(opa[0])
		);
	notech_mux2 i_10923(.S(n_31239), .A(opa[0]), .B(n_31231), .Z(n_27603));
	notech_nao3 i_28902(.A(n_336560993), .B(n_61730), .C(n_61883), .Z(n_30496
		));
	notech_reg opa_reg_1(.CP(n_63622), .D(n_27609), .CD(n_62359), .Q(opa[1])
		);
	notech_mux2 i_10931(.S(n_31239), .A(opa[1]), .B(n_31233), .Z(n_27609));
	notech_nao3 i_29025(.A(n_184060379), .B(n_316260790), .C(n_61883), .Z(n_30373
		));
	notech_reg opa_reg_2(.CP(n_63622), .D(n_27615), .CD(n_62359), .Q(opa[2])
		);
	notech_mux2 i_10939(.S(n_31239), .A(opa[2]), .B(n_31234), .Z(n_27615));
	notech_or4 i_29019(.A(n_61912), .B(n_61898), .C(n_61883), .D(n_30380), .Z
		(n_30379));
	notech_reg opa_reg_3(.CP(n_63622), .D(n_27621), .CD(n_62359), .Q(opa[3])
		);
	notech_mux2 i_10947(.S(n_31239), .A(opa[3]), .B(n_31235), .Z(n_27621));
	notech_or4 i_28895(.A(n_61883), .B(n_57672), .C(n_61717), .D(n_1850), .Z
		(n_30503));
	notech_reg opa_reg_4(.CP(n_63622), .D(n_27628), .CD(n_62359), .Q(opa[4])
		);
	notech_mux2 i_10955(.S(n_31239), .A(opa[4]), .B(n_31236), .Z(n_27628));
	notech_reg opa_reg_5(.CP(n_63622), .D(n_27639), .CD(n_62359), .Q(opa[5])
		);
	notech_mux2 i_10963(.S(n_31239), .A(opa[5]), .B(n_301460643), .Z(n_27639
		));
	notech_reg opa_reg_6(.CP(n_63622), .D(n_27645), .CD(n_62359), .Q(opa[6])
		);
	notech_mux2 i_10971(.S(n_31239), .A(opa[6]), .B(n_31237), .Z(n_27645));
	notech_and2 i_151858119(.A(n_57714), .B(instrc[116]), .Z(n_30727));
	notech_reg opa_reg_7(.CP(n_63622), .D(n_27651), .CD(n_62359), .Q(opa[7])
		);
	notech_mux2 i_10979(.S(n_31239), .A(opa[7]), .B(n_31238), .Z(n_27651));
	notech_ao4 i_176358173(.A(n_1855), .B(n_30414), .C(n_32317), .D(n_30904)
		, .Z(n_184060379));
	notech_reg opa_reg_8(.CP(n_63622), .D(n_27657), .CD(n_62359), .Q(opa[8])
		);
	notech_mux2 i_10987(.S(n_333181808), .A(n_31240), .B(opa[8]), .Z(n_27657
		));
	notech_ao4 i_154759212(.A(n_100842449), .B(n_30379), .C(n_30373), .D(\nbus_11290[2] 
		), .Z(n_183660378));
	notech_reg opa_reg_9(.CP(n_63622), .D(n_27663), .CD(n_62358), .Q(opa[9])
		);
	notech_mux2 i_10995(.S(n_333181808), .A(n_31241), .B(opa[9]), .Z(n_27663
		));
	notech_reg opa_reg_10(.CP(n_63622), .D(n_27669), .CD(n_62358), .Q(opa[10
		]));
	notech_mux2 i_11003(.S(n_333181808), .A(n_31242), .B(opa[10]), .Z(n_27669
		));
	notech_ao4 i_154859211(.A(n_30376), .B(n_33167), .C(n_30378), .D(n_58247
		), .Z(n_183160376));
	notech_reg opa_reg_11(.CP(n_63622), .D(n_27675), .CD(n_62358), .Q(opa[11
		]));
	notech_mux2 i_11011(.S(n_333181808), .A(n_31243), .B(opa[11]), .Z(n_27675
		));
	notech_ao4 i_155059209(.A(n_100542446), .B(n_30379), .C(n_30373), .D(\nbus_11290[6] 
		), .Z(n_183060375));
	notech_reg opa_reg_12(.CP(n_63622), .D(n_27681), .CD(n_62358), .Q(opa[12
		]));
	notech_mux2 i_11019(.S(n_333181808), .A(n_31244), .B(n_61016), .Z(n_27681
		));
	notech_reg opa_reg_13(.CP(n_63622), .D(n_27687), .CD(n_62358), .Q(opa[13
		]));
	notech_mux2 i_11027(.S(n_333181808), .A(n_31245), .B(n_61025), .Z(n_27687
		));
	notech_ao4 i_155159208(.A(n_30376), .B(n_33166), .C(n_30378), .D(n_58265
		), .Z(n_182560374));
	notech_reg opa_reg_14(.CP(n_63622), .D(n_27693), .CD(n_62358), .Q(opa[14
		]));
	notech_mux2 i_11035(.S(n_333181808), .A(n_31246), .B(opa[14]), .Z(n_27693
		));
	notech_ao4 i_155359206(.A(n_100242443), .B(n_30379), .C(n_30373), .D(\nbus_11290[7] 
		), .Z(n_1821));
	notech_reg opa_reg_15(.CP(n_63622), .D(n_27699), .CD(n_62359), .Q(opa[15
		]));
	notech_mux2 i_11043(.S(n_333181808), .A(n_31247), .B(n_61034), .Z(n_27699
		));
	notech_reg opa_reg_16(.CP(n_63622), .D(n_27705), .CD(n_62358), .Q(opa[16
		]));
	notech_mux2 i_11051(.S(n_31248), .A(opa[16]), .B(n_17144), .Z(n_27705)
		);
	notech_ao4 i_155459205(.A(n_30376), .B(n_33165), .C(n_30378), .D(n_58275
		), .Z(n_1814));
	notech_reg opa_reg_17(.CP(n_63676), .D(n_27711), .CD(n_62358), .Q(opa[17
		]));
	notech_mux2 i_11059(.S(n_31248), .A(opa[17]), .B(n_17150), .Z(n_27711)
		);
	notech_ao4 i_155659203(.A(n_99942440), .B(n_30503), .C(n_30496), .D(n_59032
		), .Z(n_1812));
	notech_reg opa_reg_18(.CP(n_63620), .D(n_27717), .CD(n_62362), .Q(opa[18
		]));
	notech_mux2 i_11067(.S(n_31248), .A(opa[18]), .B(n_17156), .Z(n_27717)
		);
	notech_reg opa_reg_19(.CP(n_63676), .D(n_27723), .CD(n_62363), .Q(opa[19
		]));
	notech_mux2 i_11075(.S(n_31248), .A(opa[19]), .B(n_17162), .Z(n_27723)
		);
	notech_ao4 i_155759202(.A(n_30499), .B(n_58294), .C(n_30501), .D(n_33168
		), .Z(n_1810));
	notech_reg opa_reg_20(.CP(n_63676), .D(n_27729), .CD(n_62362), .Q(opa[20
		]));
	notech_mux2 i_11083(.S(n_31248), .A(opa[20]), .B(n_17168), .Z(n_27729)
		);
	notech_reg opa_reg_21(.CP(n_63676), .D(n_27735), .CD(n_62362), .Q(opa[21
		]));
	notech_mux2 i_11091(.S(n_31248), .A(opa[21]), .B(n_17174), .Z(n_27735)
		);
	notech_ao4 i_157959181(.A(n_101142452), .B(n_30379), .C(n_30373), .D(n_58956
		), .Z(n_179760373));
	notech_reg opa_reg_22(.CP(n_63676), .D(n_27741), .CD(n_62363), .Q(opa[22
		]));
	notech_mux2 i_11099(.S(n_31248), .A(opa[22]), .B(n_17180), .Z(n_27741)
		);
	notech_reg opa_reg_23(.CP(n_63676), .D(n_27747), .CD(n_62363), .Q(opa[23
		]));
	notech_mux2 i_11107(.S(n_31248), .A(opa[23]), .B(n_17186), .Z(n_27747)
		);
	notech_ao4 i_158059180(.A(n_33169), .B(n_30376), .C(n_58238), .D(n_30378
		), .Z(n_179595933));
	notech_reg opa_reg_24(.CP(n_63676), .D(n_27756), .CD(n_62363), .Q(opa[24
		]));
	notech_mux2 i_11115(.S(n_31248), .A(opa[24]), .B(n_17192), .Z(n_27756)
		);
	notech_reg opa_reg_25(.CP(n_63676), .D(n_27762), .CD(n_62363), .Q(opa[25
		]));
	notech_mux2 i_11123(.S(n_31248), .A(opa[25]), .B(n_17198), .Z(n_27762)
		);
	notech_reg opa_reg_26(.CP(n_63676), .D(n_27768), .CD(n_62363), .Q(opa[26
		]));
	notech_mux2 i_11131(.S(n_31248), .A(opa[26]), .B(n_17204), .Z(n_27768)
		);
	notech_reg opa_reg_27(.CP(n_63676), .D(n_27774), .CD(n_62362), .Q(opa[27
		]));
	notech_mux2 i_11139(.S(n_31248), .A(opa[27]), .B(n_17210), .Z(n_27774)
		);
	notech_nand2 i_76559940(.A(n_61616), .B(read_data[0]), .Z(n_179195937)
		);
	notech_reg opa_reg_28(.CP(n_63676), .D(n_27780), .CD(n_62362), .Q(opa[28
		]));
	notech_mux2 i_11148(.S(n_31248), .A(opa[28]), .B(n_17216), .Z(n_27780)
		);
	notech_reg opa_reg_29(.CP(n_63676), .D(n_27786), .CD(n_62362), .Q(opa[29
		]));
	notech_mux2 i_11156(.S(n_31248), .A(opa[29]), .B(n_17222), .Z(n_27786)
		);
	notech_reg opa_reg_30(.CP(n_63676), .D(n_27792), .CD(n_62359), .Q(opa[30
		]));
	notech_mux2 i_11164(.S(n_31248), .A(opa[30]), .B(n_17228), .Z(n_27792)
		);
	notech_reg opa_reg_31(.CP(n_63676), .D(n_27799), .CD(n_62362), .Q(opa[31
		]));
	notech_mux2 i_11172(.S(n_31248), .A(opa[31]), .B(n_17234), .Z(n_27799)
		);
	notech_reg tcmp_reg(.CP(n_63676), .D(n_27805), .CD(n_62362), .Q(tcmp));
	notech_mux2 i_11180(.S(n_7370), .A(tcmp), .B(n_315392472), .Z(n_27805)
		);
	notech_nand2 i_73059975(.A(n_61616), .B(read_data[9]), .Z(n_178695942)
		);
	notech_reg sema_rw_reg(.CP(n_63676), .D(n_27811), .CD(n_62362), .Q(sema_rw
		));
	notech_mux2 i_11188(.S(n_31250), .A(sema_rw), .B(n_30627), .Z(n_27811)
		);
	notech_reg_set fsm_reg_0(.CP(n_63676), .D(n_27818), .SD(n_62362), .Q(fsm
		[0]));
	notech_mux2 i_11196(.S(\nbus_11314[0] ), .A(n_61898), .B(n_30434), .Z(n_27818
		));
	notech_reg_set fsm_reg_1(.CP(n_63676), .D(n_27825), .SD(n_62362), .Q(fsm
		[1]));
	notech_mux2 i_11204(.S(\nbus_11314[0] ), .A(n_61912), .B(n_13943), .Z(n_27825
		));
	notech_reg_set fsm_reg_2(.CP(n_63676), .D(n_27839), .SD(n_62362), .Q(fsm
		[2]));
	notech_mux2 i_11212(.S(\nbus_11314[0] ), .A(fsm[2]), .B(n_13949), .Z(n_27839
		));
	notech_reg_set fsm_reg_3(.CP(n_63620), .D(n_27847), .SD(n_62408), .Q(fsm
		[3]));
	notech_mux2 i_11220(.S(\nbus_11314[0] ), .A(fsm[3]), .B(n_31253), .Z(n_27847
		));
	notech_nand2 i_72559980(.A(n_61616), .B(read_data[7]), .Z(n_178195947)
		);
	notech_reg fsm_reg_4(.CP(n_63620), .D(n_27853), .CD(n_62408), .Q(fsm[4])
		);
	notech_mux2 i_11228(.S(\nbus_11314[0] ), .A(fsm[4]), .B(n_31255), .Z(n_27853
		));
	notech_reg vliw_pc_reg_0(.CP(n_63620), .D(n_27859), .CD(n_62408), .Q(vliw_pc
		[0]));
	notech_mux2 i_11236(.S(\nbus_11286[0] ), .A(vliw_pc[0]), .B(n_339281859)
		, .Z(n_27859));
	notech_reg vliw_pc_reg_1(.CP(n_63620), .D(n_27865), .CD(n_62408), .Q(vliw_pc
		[1]));
	notech_mux2 i_11244(.S(\nbus_11286[0] ), .A(vliw_pc[1]), .B(n_316092479)
		, .Z(n_27865));
	notech_reg vliw_pc_reg_2(.CP(n_63620), .D(n_27871), .CD(n_62408), .Q(vliw_pc
		[2]));
	notech_mux2 i_11252(.S(\nbus_11286[0] ), .A(vliw_pc[2]), .B(n_316192480)
		, .Z(n_27871));
	notech_reg vliw_pc_reg_3(.CP(n_63620), .D(n_27877), .CD(n_62408), .Q(vliw_pc
		[3]));
	notech_mux2 i_11260(.S(\nbus_11286[0] ), .A(vliw_pc[3]), .B(n_316292481)
		, .Z(n_27877));
	notech_nand2 i_72059985(.A(n_61616), .B(read_data[6]), .Z(n_177695950)
		);
	notech_reg vliw_pc_reg_4(.CP(n_63620), .D(n_27883), .CD(n_62408), .Q(vliw_pc
		[4]));
	notech_mux2 i_11268(.S(\nbus_11286[0] ), .A(vliw_pc[4]), .B(n_316392482)
		, .Z(n_27883));
	notech_reg_set opd_reg_0(.CP(n_63620), .D(n_27889), .SD(1'b1), .Q(opd[0]
		));
	notech_mux2 i_11276(.S(n_209580601), .A(n_21307), .B(opd[0]), .Z(n_27889
		));
	notech_reg_set opd_reg_1(.CP(n_63620), .D(n_27895), .SD(1'b1), .Q(opd[1]
		));
	notech_mux2 i_11284(.S(n_209580601), .A(n_31259), .B(opd[1]), .Z(n_27895
		));
	notech_reg_set opd_reg_2(.CP(n_63620), .D(n_27901), .SD(1'b1), .Q(opd[2]
		));
	notech_mux2 i_11292(.S(n_209580601), .A(n_21317), .B(opd[2]), .Z(n_27901
		));
	notech_reg_set opd_reg_3(.CP(n_63536), .D(n_27907), .SD(1'b1), .Q(opd[3]
		));
	notech_mux2 i_11300(.S(n_209580601), .A(n_21322), .B(opd[3]), .Z(n_27907
		));
	notech_nand2 i_71559990(.A(n_61616), .B(read_data[2]), .Z(n_1771));
	notech_reg_set opd_reg_4(.CP(n_63470), .D(n_27915), .SD(1'b1), .Q(opd[4]
		));
	notech_mux2 i_11308(.S(n_209580601), .A(n_21327), .B(opd[4]), .Z(n_27915
		));
	notech_reg_set opd_reg_5(.CP(n_63624), .D(n_27926), .SD(1'b1), .Q(opd[5]
		));
	notech_mux2 i_11316(.S(n_209580601), .A(n_21332), .B(opd[5]), .Z(n_27926
		));
	notech_reg_set opd_reg_6(.CP(n_63538), .D(n_27937), .SD(1'b1), .Q(opd[6]
		));
	notech_mux2 i_11324(.S(\nbus_11356[6] ), .A(opd[6]), .B(n_21337), .Z(n_27937
		));
	notech_reg_set opd_reg_7(.CP(n_63538), .D(n_27943), .SD(1'b1), .Q(opd[7]
		));
	notech_mux2 i_11333(.S(\nbus_11356[6] ), .A(opd[7]), .B(n_21342), .Z(n_27943
		));
	notech_reg_set opd_reg_8(.CP(n_63538), .D(n_27949), .SD(1'b1), .Q(opd[8]
		));
	notech_mux2 i_11341(.S(\nbus_11356[6] ), .A(opd[8]), .B(n_21347), .Z(n_27949
		));
	notech_nor2 i_140160726(.A(n_1854), .B(n_1852), .Z(n_176660368));
	notech_reg_set opd_reg_9(.CP(n_63538), .D(n_27955), .SD(1'b1), .Q(opd[9]
		));
	notech_mux2 i_11349(.S(\nbus_11356[6] ), .A(opd[9]), .B(n_21352), .Z(n_27955
		));
	notech_reg_set opd_reg_10(.CP(n_63538), .D(n_27961), .SD(1'b1), .Q(opd[
		10]));
	notech_mux2 i_11357(.S(\nbus_11356[6] ), .A(opd[10]), .B(n_21357), .Z(n_27961
		));
	notech_reg_set opd_reg_11(.CP(n_63538), .D(n_27970), .SD(1'b1), .Q(opd[
		11]));
	notech_mux2 i_11365(.S(\nbus_11356[6] ), .A(opd[11]), .B(n_21362), .Z(n_27970
		));
	notech_nor2 i_141960652(.A(n_57714), .B(n_57686), .Z(n_28557));
	notech_reg_set opd_reg_12(.CP(n_63538), .D(n_27978), .SD(1'b1), .Q(opd[
		12]));
	notech_mux2 i_11373(.S(\nbus_11356[6] ), .A(opd[12]), .B(n_21367), .Z(n_27978
		));
	notech_or2 i_128260656(.A(n_334560973), .B(n_30340), .Z(n_23519));
	notech_reg_set opd_reg_13(.CP(n_63538), .D(n_27986), .SD(1'b1), .Q(opd[
		13]));
	notech_mux2 i_11382(.S(\nbus_11356[6] ), .A(opd[13]), .B(n_21372), .Z(n_27986
		));
	notech_ao4 i_176660738(.A(n_1854), .B(n_1852), .C(n_32317), .D(n_30904),
		 .Z(n_176360365));
	notech_reg_set opd_reg_14(.CP(n_63538), .D(n_27993), .SD(1'b1), .Q(opd[
		14]));
	notech_mux2 i_11390(.S(\nbus_11356[6] ), .A(opd[14]), .B(n_21377), .Z(n_27993
		));
	notech_nao3 i_31660695(.A(n_176360365), .B(n_61730), .C(n_61883), .Z(n_30378
		));
	notech_reg_set opd_reg_15(.CP(n_63624), .D(n_28000), .SD(1'b1), .Q(opd[
		15]));
	notech_mux2 i_11398(.S(\nbus_11356[6] ), .A(opd[15]), .B(n_21382), .Z(n_28000
		));
	notech_or4 i_31560696(.A(n_61912), .B(n_61898), .C(n_61880), .D(n_2805),
		 .Z(n_30376));
	notech_reg_set opd_reg_16(.CP(n_63624), .D(n_28010), .SD(1'b1), .Q(opd[
		16]));
	notech_mux2 i_11406(.S(n_4457), .A(n_21387), .B(opd[16]), .Z(n_28010));
	notech_or4 i_31460697(.A(n_61883), .B(n_57672), .C(n_335660984), .D(n_61717
		), .Z(n_30501));
	notech_reg_set opd_reg_17(.CP(n_63624), .D(n_28016), .SD(1'b1), .Q(opd[
		17]));
	notech_mux2 i_11414(.S(n_4457), .A(n_21392), .B(opd[17]), .Z(n_28016));
	notech_nao3 i_31360698(.A(n_335960987), .B(n_61730), .C(n_61883), .Z(n_30499
		));
	notech_reg_set opd_reg_18(.CP(n_63624), .D(n_28022), .SD(1'b1), .Q(opd[
		18]));
	notech_mux2 i_11422(.S(n_4457), .A(n_21397), .B(opd[18]), .Z(n_28022));
	notech_reg_set opd_reg_19(.CP(n_63624), .D(n_28028), .SD(1'b1), .Q(opd[
		19]));
	notech_mux2 i_11430(.S(n_4457), .A(n_21402), .B(opd[19]), .Z(n_28028));
	notech_ao3 i_95262440(.A(n_30274), .B(n_1661), .C(n_335060978), .Z(n_176160363
		));
	notech_reg_set opd_reg_20(.CP(n_63624), .D(n_28034), .SD(1'b1), .Q(opd[
		20]));
	notech_mux2 i_11439(.S(n_4457), .A(n_21407), .B(opd[20]), .Z(n_28034));
	notech_reg_set opd_reg_21(.CP(n_63624), .D(n_28040), .SD(1'b1), .Q(opd[
		21]));
	notech_mux2 i_11447(.S(n_4457), .A(n_21412), .B(opd[21]), .Z(n_28040));
	notech_reg_set opd_reg_22(.CP(n_63624), .D(n_28046), .SD(1'b1), .Q(opd[
		22]));
	notech_mux2 i_11455(.S(n_4457), .A(n_21417), .B(opd[22]), .Z(n_28046));
	notech_ao4 i_95362439(.A(n_58664), .B(nbus_11271[1]), .C(n_334560973), .D
		(n_30891), .Z(n_175860360));
	notech_reg_set opd_reg_23(.CP(n_63624), .D(n_28052), .SD(1'b1), .Q(opd[
		23]));
	notech_mux2 i_11463(.S(n_4457), .A(n_21422), .B(opd[23]), .Z(n_28052));
	notech_ao4 i_95462438(.A(n_30916), .B(n_23511), .C(n_334460972), .D(n_56956
		), .Z(n_175760359));
	notech_reg_set opd_reg_24(.CP(n_63624), .D(n_28058), .SD(1'b1), .Q(opd[
		24]));
	notech_mux2 i_11471(.S(n_4457), .A(n_21427), .B(opd[24]), .Z(n_28058));
	notech_and4 i_96362429(.A(n_175260356), .B(n_175160355), .C(n_174960353)
		, .D(n_174860352), .Z(n_175660358));
	notech_reg_set opd_reg_25(.CP(n_63624), .D(n_28064), .SD(1'b1), .Q(opd[
		25]));
	notech_mux2 i_11479(.S(n_4457), .A(n_21432), .B(opd[25]), .Z(n_28064));
	notech_reg_set opd_reg_26(.CP(n_63624), .D(n_28070), .SD(1'b1), .Q(opd[
		26]));
	notech_mux2 i_11487(.S(n_4457), .A(n_21437), .B(opd[26]), .Z(n_28070));
	notech_ao4 i_95762435(.A(n_30896), .B(n_23519), .C(n_30914), .D(n_23510)
		, .Z(n_175260356));
	notech_reg_set opd_reg_27(.CP(n_63624), .D(n_28076), .SD(1'b1), .Q(opd[
		27]));
	notech_mux2 i_11495(.S(n_4457), .A(n_21442), .B(opd[27]), .Z(n_28076));
	notech_ao4 i_95862434(.A(n_391264443), .B(n_33103), .C(n_391164442), .D(n_334360971
		), .Z(n_175160355));
	notech_reg_set opd_reg_28(.CP(n_63624), .D(n_28083), .SD(1'b1), .Q(opd[
		28]));
	notech_mux2 i_11503(.S(n_4457), .A(n_21447), .B(opd[28]), .Z(n_28083));
	notech_reg_set opd_reg_29(.CP(n_63624), .D(n_28091), .SD(1'b1), .Q(opd[
		29]));
	notech_mux2 i_11511(.S(n_4457), .A(n_21452), .B(opd[29]), .Z(n_28091));
	notech_ao4 i_96062432(.A(n_335260980), .B(n_59005), .C(n_335160979), .D(n_58229
		), .Z(n_174960353));
	notech_reg_set opd_reg_30(.CP(n_63624), .D(n_28100), .SD(1'b1), .Q(opd[
		30]));
	notech_mux2 i_11519(.S(n_4457), .A(n_21457), .B(opd[30]), .Z(n_28100));
	notech_ao4 i_96162431(.A(n_58696), .B(n_30280), .C(n_164896005), .D(n_23760
		), .Z(n_174860352));
	notech_reg_set opd_reg_31(.CP(n_63624), .D(n_28107), .SD(1'b1), .Q(opd[
		31]));
	notech_mux2 i_11527(.S(n_4457), .A(n_218780688), .B(n_58018), .Z(n_28107
		));
	notech_reg io_add_reg_0(.CP(n_63624), .D(n_28113), .CD(n_62408), .Q(io_add
		[0]));
	notech_mux2 i_11535(.S(n_31260), .A(io_add[0]), .B(n_326895684), .Z(n_28113
		));
	notech_and3 i_107662325(.A(n_28190), .B(n_174460348), .C(n_167495980), .Z
		(n_174660350));
	notech_reg io_add_reg_1(.CP(n_63538), .D(n_28120), .CD(n_62408), .Q(io_add
		[1]));
	notech_mux2 i_11543(.S(n_31260), .A(io_add[1]), .B(n_326995685), .Z(n_28120
		));
	notech_reg io_add_reg_2(.CP(n_63538), .D(n_28126), .CD(n_62408), .Q(io_add
		[2]));
	notech_mux2 i_11551(.S(n_31260), .A(io_add[2]), .B(n_327095686), .Z(n_28126
		));
	notech_ao4 i_107562326(.A(n_24527), .B(n_33102), .C(n_60453), .D(n_31512
		), .Z(n_174460348));
	notech_reg io_add_reg_3(.CP(n_63540), .D(n_28132), .CD(n_62407), .Q(io_add
		[3]));
	notech_mux2 i_11559(.S(n_31260), .A(io_add[3]), .B(n_327195687), .Z(n_28132
		));
	notech_reg io_add_reg_4(.CP(n_63540), .D(n_28138), .CD(n_62407), .Q(io_add
		[4]));
	notech_mux2 i_11567(.S(n_31260), .A(io_add[4]), .B(n_327295688), .Z(n_28138
		));
	notech_ao4 i_107762324(.A(n_334760975), .B(n_24717), .C(n_61094), .D(n_30763
		), .Z(n_174260346));
	notech_reg io_add_reg_5(.CP(n_63540), .D(n_28145), .CD(n_62407), .Q(io_add
		[5]));
	notech_mux2 i_11575(.S(n_31260), .A(io_add[5]), .B(n_327395689), .Z(n_28145
		));
	notech_ao4 i_107862323(.A(n_381164342), .B(n_56974), .C(n_380764338), .D
		(n_31047), .Z(n_174160345));
	notech_reg io_add_reg_6(.CP(n_63540), .D(n_28151), .CD(n_62407), .Q(io_add
		[6]));
	notech_mux2 i_11583(.S(n_31260), .A(io_add[6]), .B(n_327495690), .Z(n_28151
		));
	notech_and3 i_108862313(.A(n_173860342), .B(n_173760341), .C(n_173660340
		), .Z(n_174060344));
	notech_reg io_add_reg_7(.CP(n_63540), .D(n_28157), .CD(n_62407), .Q(io_add
		[7]));
	notech_mux2 i_11591(.S(n_31260), .A(io_add[7]), .B(n_21074), .Z(n_28157)
		);
	notech_reg io_add_reg_8(.CP(n_63540), .D(n_28164), .CD(n_62408), .Q(io_add
		[8]));
	notech_mux2 i_11599(.S(n_31260), .A(io_add[8]), .B(n_327595691), .Z(n_28164
		));
	notech_ao4 i_108162320(.A(n_381064341), .B(n_33104), .C(n_334660974), .D
		(n_380964340), .Z(n_173860342));
	notech_reg io_add_reg_9(.CP(n_63540), .D(n_28170), .CD(n_62408), .Q(io_add
		[9]));
	notech_mux2 i_11607(.S(n_31260), .A(io_add[9]), .B(n_327695692), .Z(n_28170
		));
	notech_ao4 i_108262319(.A(n_24430), .B(n_31048), .C(n_24424), .D(n_31067
		), .Z(n_173760341));
	notech_reg io_add_reg_10(.CP(n_63540), .D(n_28176), .CD(n_62407), .Q(io_add
		[10]));
	notech_mux2 i_11615(.S(n_31260), .A(io_add[10]), .B(n_327795693), .Z(n_28176
		));
	notech_and3 i_108762314(.A(n_168995966), .B(n_173360337), .C(n_173560339
		), .Z(n_173660340));
	notech_reg io_add_reg_11(.CP(n_63540), .D(n_28182), .CD(n_62407), .Q(io_add
		[11]));
	notech_mux2 i_11623(.S(n_31260), .A(io_add[11]), .B(n_327895694), .Z(n_28182
		));
	notech_ao4 i_108462317(.A(n_24421), .B(n_31068), .C(n_24431), .D(n_31071
		), .Z(n_173560339));
	notech_reg io_add_reg_12(.CP(n_63540), .D(n_28188), .CD(n_62409), .Q(io_add
		[12]));
	notech_mux2 i_11631(.S(n_31260), .A(io_add[12]), .B(n_327995695), .Z(n_28188
		));
	notech_reg io_add_reg_13(.CP(n_63540), .D(n_28195), .CD(n_62409), .Q(io_add
		[13]));
	notech_mux2 i_11639(.S(n_31260), .A(io_add[13]), .B(n_328095696), .Z(n_28195
		));
	notech_ao4 i_108562316(.A(n_24429), .B(n_31075), .C(n_24425), .D(n_31072
		), .Z(n_173360337));
	notech_reg io_add_reg_14(.CP(n_63540), .D(n_28201), .CD(n_62409), .Q(io_add
		[14]));
	notech_mux2 i_11647(.S(n_31260), .A(io_add[14]), .B(n_328195697), .Z(n_28201
		));
	notech_and4 i_109662305(.A(n_28206), .B(n_58055), .C(n_172960333), .D(n_172860332
		), .Z(n_173260336));
	notech_reg io_add_reg_15(.CP(n_63540), .D(n_28208), .CD(n_62409), .Q(io_add
		[15]));
	notech_mux2 i_11655(.S(n_31260), .A(io_add[15]), .B(n_328295698), .Z(n_28208
		));
	notech_reg_set temp_ss_reg_0(.CP(n_63540), .D(n_28214), .SD(1'b1), .Q(temp_ss
		[0]));
	notech_mux2 i_11663(.S(n_31293), .A(temp_ss[0]), .B(n_311492440), .Z(n_28214
		));
	notech_reg_set temp_ss_reg_1(.CP(n_63540), .D(n_28220), .SD(1'b1), .Q(temp_ss
		[1]));
	notech_mux2 i_11671(.S(n_31293), .A(temp_ss[1]), .B(n_311592441), .Z(n_28220
		));
	notech_ao4 i_109062311(.A(n_24528), .B(n_33101), .C(n_24527), .D(n_33100
		), .Z(n_172960333));
	notech_reg_set temp_ss_reg_2(.CP(n_63540), .D(n_28226), .SD(1'b1), .Q(temp_ss
		[2]));
	notech_mux2 i_11679(.S(n_31293), .A(temp_ss[2]), .B(n_311692442), .Z(n_28226
		));
	notech_and3 i_109562306(.A(n_172560329), .B(n_172760331), .C(n_1696), .Z
		(n_172860332));
	notech_reg_set temp_ss_reg_3(.CP(n_63540), .D(n_28232), .SD(1'b1), .Q(temp_ss
		[3]));
	notech_mux2 i_11687(.S(n_31293), .A(temp_ss[3]), .B(n_311792443), .Z(n_28232
		));
	notech_ao4 i_109262309(.A(n_60453), .B(n_31513), .C(n_24717), .D(n_334960977
		), .Z(n_172760331));
	notech_reg_set temp_ss_reg_4(.CP(n_63540), .D(n_28239), .SD(1'b1), .Q(temp_ss
		[4]));
	notech_mux2 i_11695(.S(n_31293), .A(temp_ss[4]), .B(n_311892444), .Z(n_28239
		));
	notech_reg_set temp_ss_reg_5(.CP(n_63540), .D(n_28246), .SD(1'b1), .Q(temp_ss
		[5]));
	notech_mux2 i_11703(.S(n_31293), .A(temp_ss[5]), .B(n_311992445), .Z(n_28246
		));
	notech_ao4 i_109362308(.A(n_381164342), .B(n_56983), .C(n_31098), .D(n_380764338
		), .Z(n_172560329));
	notech_reg_set temp_ss_reg_6(.CP(n_63470), .D(n_28254), .SD(1'b1), .Q(temp_ss
		[6]));
	notech_mux2 i_11712(.S(n_31293), .A(temp_ss[6]), .B(n_312092446), .Z(n_28254
		));
	notech_reg_set temp_ss_reg_7(.CP(n_63470), .D(n_28265), .SD(1'b1), .Q(temp_ss
		[7]));
	notech_mux2 i_11720(.S(n_31293), .A(temp_ss[7]), .B(n_312192447), .Z(n_28265
		));
	notech_reg_set temp_ss_reg_8(.CP(n_63470), .D(n_28271), .SD(1'b1), .Q(temp_ss
		[8]));
	notech_mux2 i_11728(.S(n_31293), .A(temp_ss[8]), .B(n_312292448), .Z(n_28271
		));
	notech_ao4 i_109762304(.A(n_381064341), .B(n_33135), .C(n_334860976), .D
		(n_380964340), .Z(n_172260326));
	notech_reg_set temp_ss_reg_9(.CP(n_63470), .D(n_28277), .SD(1'b1), .Q(temp_ss
		[9]));
	notech_mux2 i_11736(.S(n_31293), .A(temp_ss[9]), .B(n_312392449), .Z(n_28277
		));
	notech_ao4 i_109862303(.A(n_31099), .B(n_24430), .C(n_31118), .D(n_24424
		), .Z(n_172160325));
	notech_reg_set temp_ss_reg_10(.CP(n_63470), .D(n_28283), .SD(1'b1), .Q(temp_ss
		[10]));
	notech_mux2 i_11744(.S(n_31293), .A(temp_ss[10]), .B(n_312492450), .Z(n_28283
		));
	notech_and3 i_110362298(.A(n_170595953), .B(n_171760321), .C(n_171960323
		), .Z(n_172060324));
	notech_reg_set temp_ss_reg_11(.CP(n_63470), .D(n_28289), .SD(1'b1), .Q(temp_ss
		[11]));
	notech_mux2 i_11752(.S(n_31293), .A(temp_ss[11]), .B(n_312592451), .Z(n_28289
		));
	notech_ao4 i_110062301(.A(n_31119), .B(n_24421), .C(n_31122), .D(n_24431
		), .Z(n_171960323));
	notech_reg_set temp_ss_reg_12(.CP(n_63470), .D(n_28295), .SD(1'b1), .Q(temp_ss
		[12]));
	notech_mux2 i_11760(.S(n_31293), .A(temp_ss[12]), .B(n_312792452), .Z(n_28295
		));
	notech_reg_set temp_ss_reg_13(.CP(n_63470), .D(n_28301), .SD(1'b1), .Q(temp_ss
		[13]));
	notech_mux2 i_11768(.S(n_31293), .A(temp_ss[13]), .B(n_312892453), .Z(n_28301
		));
	notech_ao4 i_110162300(.A(n_31126), .B(n_24429), .C(n_31123), .D(n_24425
		), .Z(n_171760321));
	notech_reg_set temp_ss_reg_14(.CP(n_63470), .D(n_28307), .SD(1'b1), .Q(temp_ss
		[14]));
	notech_mux2 i_11776(.S(n_31293), .A(temp_ss[14]), .B(n_312992454), .Z(n_28307
		));
	notech_ao4 i_170061715(.A(n_30378), .B(n_58229), .C(n_30376), .D(n_33103
		), .Z(n_171660320));
	notech_reg_set temp_ss_reg_15(.CP(n_63620), .D(n_28313), .SD(1'b1), .Q(temp_ss
		[15]));
	notech_mux2 i_11785(.S(n_31293), .A(temp_ss[15]), .B(n_313192455), .Z(n_28313
		));
	notech_reg_set temp_ss_reg_16(.CP(n_63528), .D(n_28319), .SD(1'b1), .Q(temp_ss
		[16]));
	notech_mux2 i_11793(.S(n_54423), .A(temp_ss[16]), .B(n_313392456), .Z(n_28319
		));
	notech_ao4 i_170161714(.A(n_30373), .B(n_59005), .C(n_61660), .D(n_31509
		), .Z(n_171460318));
	notech_reg_set temp_ss_reg_17(.CP(n_63468), .D(n_28325), .SD(1'b1), .Q(temp_ss
		[17]));
	notech_mux2 i_11801(.S(n_54423), .A(temp_ss[17]), .B(n_313592457), .Z(n_28325
		));
	notech_ao4 i_172761688(.A(n_32544), .B(n_165695997), .C(n_60188), .D(n_28555
		), .Z(n_171360317));
	notech_reg_set temp_ss_reg_18(.CP(n_63528), .D(n_28331), .SD(1'b1), .Q(temp_ss
		[18]));
	notech_mux2 i_11809(.S(n_54423), .A(temp_ss[18]), .B(n_313792458), .Z(n_28331
		));
	notech_reg_set temp_ss_reg_19(.CP(n_63528), .D(n_28338), .SD(1'b1), .Q(temp_ss
		[19]));
	notech_mux2 i_11818(.S(n_54423), .A(temp_ss[19]), .B(n_313892459), .Z(n_28338
		));
	notech_or4 i_33122(.A(n_58583), .B(n_332160949), .C(n_61786), .D(n_61766
		), .Z(n_26276));
	notech_reg_set temp_ss_reg_20(.CP(n_63528), .D(n_28344), .SD(1'b1), .Q(temp_ss
		[20]));
	notech_mux2 i_11826(.S(n_54423), .A(temp_ss[20]), .B(n_313992460), .Z(n_28344
		));
	notech_or2 i_33123(.A(n_332160949), .B(n_32273), .Z(n_26275));
	notech_reg_set temp_ss_reg_21(.CP(n_63528), .D(n_28350), .SD(1'b1), .Q(temp_ss
		[21]));
	notech_mux2 i_11835(.S(n_54423), .A(temp_ss[21]), .B(n_314092461), .Z(n_28350
		));
	notech_or2 i_9063267(.A(n_332160949), .B(n_30788), .Z(n_26278));
	notech_reg_set temp_ss_reg_22(.CP(n_63528), .D(n_28356), .SD(1'b1), .Q(temp_ss
		[22]));
	notech_mux2 i_11843(.S(n_54423), .A(temp_ss[22]), .B(n_314192462), .Z(n_28356
		));
	notech_or4 i_33121(.A(n_58583), .B(n_26278), .C(n_61786), .D(n_61766), .Z
		(n_26277));
	notech_reg_set temp_ss_reg_23(.CP(n_63528), .D(n_28362), .SD(1'b1), .Q(temp_ss
		[23]));
	notech_mux2 i_11851(.S(n_54423), .A(temp_ss[23]), .B(n_314492463), .Z(n_28362
		));
	notech_nao3 i_33126(.A(n_56002), .B(n_57429), .C(n_332160949), .Z(n_26272
		));
	notech_reg_set temp_ss_reg_24(.CP(n_63528), .D(n_28371), .SD(1'b1), .Q(temp_ss
		[24]));
	notech_mux2 i_11860(.S(n_54423), .A(temp_ss[24]), .B(n_314592464), .Z(n_28371
		));
	notech_or2 i_33127(.A(n_26624), .B(n_56002), .Z(n_26271));
	notech_reg_set temp_ss_reg_25(.CP(n_63528), .D(n_28377), .SD(1'b1), .Q(temp_ss
		[25]));
	notech_mux2 i_11868(.S(n_54423), .A(temp_ss[25]), .B(n_314692465), .Z(n_28377
		));
	notech_or2 i_33130(.A(n_332160949), .B(n_56002), .Z(n_26268));
	notech_reg_set temp_ss_reg_26(.CP(n_63528), .D(n_28383), .SD(1'b1), .Q(temp_ss
		[26]));
	notech_mux2 i_11876(.S(n_54423), .A(temp_ss[26]), .B(n_314792466), .Z(n_28383
		));
	notech_nor2 i_12963230(.A(n_332760955), .B(n_28533), .Z(n_171160315));
	notech_reg_set temp_ss_reg_27(.CP(n_63612), .D(n_28389), .SD(1'b1), .Q(temp_ss
		[27]));
	notech_mux2 i_11884(.S(n_54423), .A(temp_ss[27]), .B(n_314892467), .Z(n_28389
		));
	notech_nao3 i_5263305(.A(n_32323), .B(n_32310), .C(n_334060968), .Z(n_30280
		));
	notech_reg_set temp_ss_reg_28(.CP(n_63612), .D(n_28395), .SD(1'b1), .Q(temp_ss
		[28]));
	notech_mux2 i_11892(.S(n_54423), .A(temp_ss[28]), .B(n_314992468), .Z(n_28395
		));
	notech_or2 i_92762465(.A(n_334360971), .B(n_30379), .Z(n_171060314));
	notech_reg_set temp_ss_reg_29(.CP(n_63612), .D(n_28401), .SD(1'b1), .Q(temp_ss
		[29]));
	notech_mux2 i_11900(.S(n_54423), .A(temp_ss[29]), .B(n_315092469), .Z(n_28401
		));
	notech_reg_set temp_ss_reg_30(.CP(n_63612), .D(n_28407), .SD(1'b1), .Q(temp_ss
		[30]));
	notech_mux2 i_11908(.S(n_54423), .A(temp_ss[30]), .B(n_315192470), .Z(n_28407
		));
	notech_reg_set temp_ss_reg_31(.CP(n_63612), .D(n_28413), .SD(1'b1), .Q(temp_ss
		[31]));
	notech_mux2 i_11916(.S(n_54423), .A(temp_ss[31]), .B(n_315292471), .Z(n_28413
		));
	notech_reg errco_reg_0(.CP(n_63612), .D(n_28419), .CD(n_62410), .Q(errco
		[0]));
	notech_mux2 i_11924(.S(n_55811), .A(errco[0]), .B(n_16495863), .Z(n_28419
		));
	notech_reg errco_reg_1(.CP(n_63612), .D(n_28425), .CD(n_62410), .Q(errco
		[1]));
	notech_mux2 i_11932(.S(n_55811), .A(errco[1]), .B(wr_fault), .Z(n_28425)
		);
	notech_ao4 i_31192(.A(n_28240), .B(nbus_11273[5]), .C(\nbus_11290[5] ), 
		.D(n_331360941), .Z(n_28206));
	notech_reg errco_reg_2(.CP(n_63612), .D(n_28431), .CD(n_62410), .Q(errco
		[2]));
	notech_mux2 i_11940(.S(n_55811), .A(errco[2]), .B(cs[1]), .Z(n_28431));
	notech_ao4 i_31208(.A(n_28240), .B(nbus_11273[4]), .C(n_331360941), .D(\nbus_11290[4] 
		), .Z(n_28190));
	notech_reg errco_reg_3(.CP(n_63612), .D(n_28440), .CD(n_62410), .Q(errco
		[3]));
	notech_ao3 i_11950(.A(n_61094), .B(errco[3]), .C(n_61447), .Z(n_28440)
		);
	notech_or4 i_31363054(.A(n_24430), .B(n_61056), .C(\nbus_11290[5] ), .D(n_58574
		), .Z(n_170595953));
	notech_reg errco_reg_4(.CP(n_63612), .D(n_28443), .CD(n_62410), .Q(errco
		[4]));
	notech_mux2 i_11956(.S(n_55811), .A(errco[4]), .B(n_61447), .Z(n_28443)
		);
	notech_reg errco_reg_5(.CP(n_63612), .D(n_28452), .CD(n_62409), .Q(errco
		[5]));
	notech_ao3 i_11966(.A(n_61094), .B(errco[5]), .C(n_61447), .Z(n_28452)
		);
	notech_reg errco_reg_6(.CP(n_63612), .D(n_28458), .CD(n_62409), .Q(errco
		[6]));
	notech_ao3 i_11974(.A(n_61094), .B(errco[6]), .C(n_61455), .Z(n_28458)
		);
	notech_reg errco_reg_7(.CP(n_63612), .D(n_28464), .CD(n_62409), .Q(errco
		[7]));
	notech_ao3 i_11982(.A(n_61094), .B(errco[7]), .C(n_61447), .Z(n_28464)
		);
	notech_reg errco_reg_8(.CP(n_63612), .D(n_28470), .CD(n_62408), .Q(errco
		[8]));
	notech_ao3 i_11991(.A(n_61094), .B(errco[8]), .C(n_61447), .Z(n_28470)
		);
	notech_reg errco_reg_9(.CP(n_63612), .D(n_28476), .CD(n_62409), .Q(errco
		[9]));
	notech_ao3 i_11999(.A(n_61094), .B(errco[9]), .C(n_61447), .Z(n_28476)
		);
	notech_reg errco_reg_10(.CP(n_63612), .D(n_28482), .CD(n_62409), .Q(errco
		[10]));
	notech_ao3 i_12007(.A(n_61094), .B(errco[10]), .C(n_61447), .Z(n_28482)
		);
	notech_reg errco_reg_11(.CP(n_63612), .D(n_28488), .CD(n_62409), .Q(errco
		[11]));
	notech_ao3 i_12015(.A(n_61094), .B(errco[11]), .C(n_61447), .Z(n_28488)
		);
	notech_reg errco_reg_12(.CP(n_63612), .D(n_28494), .CD(n_62409), .Q(errco
		[12]));
	notech_ao3 i_12023(.A(n_61094), .B(errco[12]), .C(n_61447), .Z(n_28494)
		);
	notech_nand2 i_32263045(.A(sav_ecx[5]), .B(n_61864), .Z(n_1696));
	notech_reg errco_reg_13(.CP(n_63612), .D(n_28500), .CD(n_62409), .Q(errco
		[13]));
	notech_ao3 i_12031(.A(n_61092), .B(errco[13]), .C(n_61447), .Z(n_28500)
		);
	notech_reg errco_reg_14(.CP(n_63610), .D(n_28506), .CD(n_62409), .Q(errco
		[14]));
	notech_ao3 i_12039(.A(n_61091), .B(errco[14]), .C(n_61447), .Z(n_28506)
		);
	notech_reg errco_reg_15(.CP(n_63610), .D(n_28512), .CD(n_62403), .Q(errco
		[15]));
	notech_ao3 i_12047(.A(n_61091), .B(errco[15]), .C(n_61447), .Z(n_28512)
		);
	notech_reg errco_reg_16(.CP(n_63672), .D(n_28518), .CD(n_62403), .Q(errco
		[16]));
	notech_ao3 i_12055(.A(n_61091), .B(errco[16]), .C(n_61447), .Z(n_28518)
		);
	notech_reg errco_reg_17(.CP(n_63672), .D(n_28524), .CD(n_62403), .Q(errco
		[17]));
	notech_ao3 i_12063(.A(n_61092), .B(errco[17]), .C(n_61455), .Z(n_28524)
		);
	notech_reg errco_reg_18(.CP(n_63672), .D(n_28530), .CD(n_62403), .Q(errco
		[18]));
	notech_ao3 i_12071(.A(n_61092), .B(errco[18]), .C(n_61451), .Z(n_28530)
		);
	notech_reg errco_reg_19(.CP(n_63672), .D(n_28538), .CD(n_62403), .Q(errco
		[19]));
	notech_ao3 i_12079(.A(n_61091), .B(errco[19]), .C(n_61451), .Z(n_28538)
		);
	notech_or4 i_29563070(.A(n_24430), .B(n_61052), .C(n_58574), .D(\nbus_11290[4] 
		), .Z(n_168995966));
	notech_reg errco_reg_20(.CP(n_63672), .D(n_28544), .CD(n_62403), .Q(errco
		[20]));
	notech_ao3 i_12087(.A(n_61091), .B(errco[20]), .C(n_61451), .Z(n_28544)
		);
	notech_reg errco_reg_21(.CP(n_63672), .D(n_28550), .CD(n_62403), .Q(errco
		[21]));
	notech_ao3 i_12095(.A(n_61091), .B(errco[21]), .C(n_61451), .Z(n_28550)
		);
	notech_reg errco_reg_22(.CP(n_63672), .D(n_28562), .CD(n_62403), .Q(errco
		[22]));
	notech_ao3 i_12103(.A(n_61091), .B(errco[22]), .C(n_61451), .Z(n_28562)
		);
	notech_reg errco_reg_23(.CP(n_63672), .D(n_28568), .CD(n_62403), .Q(errco
		[23]));
	notech_ao3 i_12111(.A(n_61091), .B(errco[23]), .C(n_61451), .Z(n_28568)
		);
	notech_reg errco_reg_24(.CP(n_63672), .D(n_28575), .CD(n_62403), .Q(errco
		[24]));
	notech_ao3 i_12119(.A(n_61091), .B(errco[24]), .C(n_61451), .Z(n_28575)
		);
	notech_reg errco_reg_25(.CP(n_63672), .D(n_28582), .CD(n_62402), .Q(errco
		[25]));
	notech_ao3 i_12127(.A(n_61092), .B(errco[25]), .C(n_61451), .Z(n_28582)
		);
	notech_reg errco_reg_26(.CP(n_63672), .D(n_28588), .CD(n_62402), .Q(errco
		[26]));
	notech_ao3 i_12135(.A(n_61092), .B(errco[26]), .C(n_61455), .Z(n_28588)
		);
	notech_reg errco_reg_27(.CP(n_63378), .D(n_28594), .CD(n_62402), .Q(errco
		[27]));
	notech_ao3 i_12143(.A(n_61092), .B(errco[27]), .C(n_61455), .Z(n_28594)
		);
	notech_reg errco_reg_28(.CP(n_63672), .D(n_28600), .CD(n_62402), .Q(errco
		[28]));
	notech_ao3 i_12151(.A(n_61092), .B(errco[28]), .C(n_61455), .Z(n_28600)
		);
	notech_reg errco_reg_29(.CP(n_63672), .D(n_28606), .CD(n_62402), .Q(errco
		[29]));
	notech_ao3 i_12159(.A(n_61092), .B(errco[29]), .C(n_61455), .Z(n_28606)
		);
	notech_reg errco_reg_30(.CP(n_63672), .D(n_28612), .CD(n_62403), .Q(errco
		[30]));
	notech_ao3 i_12167(.A(n_61092), .B(errco[30]), .C(n_61451), .Z(n_28612)
		);
	notech_reg errco_reg_31(.CP(n_63672), .D(n_28618), .CD(n_62403), .Q(errco
		[31]));
	notech_ao3 i_12175(.A(n_61092), .B(errco[31]), .C(n_61451), .Z(n_28618)
		);
	notech_reg_set write_data_reg_0(.CP(n_63672), .D(n_28621), .SD(1'b1), .Q
		(write_data[0]));
	notech_mux2 i_12181(.S(n_31326), .A(write_data[0]), .B(n_20844), .Z(n_28621
		));
	notech_reg_set write_data_reg_1(.CP(n_63672), .D(n_28627), .SD(1'b1), .Q
		(write_data[1]));
	notech_mux2 i_12190(.S(n_31326), .A(write_data[1]), .B(n_20849), .Z(n_28627
		));
	notech_reg_set write_data_reg_2(.CP(n_63610), .D(n_28633), .SD(1'b1), .Q
		(write_data[2]));
	notech_mux2 i_12198(.S(n_31326), .A(write_data[2]), .B(n_20854), .Z(n_28633
		));
	notech_nao3 i_31063057(.A(n_3476), .B(n_61279), .C(n_32186), .Z(n_167495980
		));
	notech_reg_set write_data_reg_3(.CP(n_63610), .D(n_28639), .SD(1'b1), .Q
		(write_data[3]));
	notech_mux2 i_12206(.S(n_31326), .A(write_data[3]), .B(n_20859), .Z(n_28639
		));
	notech_reg_set write_data_reg_4(.CP(n_63610), .D(n_28645), .SD(1'b1), .Q
		(write_data[4]));
	notech_mux2 i_12214(.S(n_31326), .A(write_data[4]), .B(n_20864), .Z(n_28645
		));
	notech_reg_set write_data_reg_5(.CP(n_63610), .D(n_28651), .SD(1'b1), .Q
		(write_data[5]));
	notech_mux2 i_12222(.S(n_31326), .A(write_data[5]), .B(n_20869), .Z(n_28651
		));
	notech_reg_set write_data_reg_6(.CP(n_63610), .D(n_28657), .SD(1'b1), .Q
		(write_data[6]));
	notech_mux2 i_12230(.S(n_31326), .A(write_data[6]), .B(n_20874), .Z(n_28657
		));
	notech_reg_set write_data_reg_7(.CP(n_63610), .D(n_28663), .SD(1'b1), .Q
		(write_data[7]));
	notech_mux2 i_12238(.S(n_31326), .A(write_data[7]), .B(n_20879), .Z(n_28663
		));
	notech_reg_set write_data_reg_8(.CP(n_63610), .D(n_28669), .SD(1'b1), .Q
		(write_data[8]));
	notech_mux2 i_12246(.S(n_31326), .A(write_data[8]), .B(n_20884), .Z(n_28669
		));
	notech_reg_set write_data_reg_9(.CP(n_63610), .D(n_28675), .SD(1'b1), .Q
		(write_data[9]));
	notech_mux2 i_12254(.S(n_31326), .A(write_data[9]), .B(n_20889), .Z(n_28675
		));
	notech_reg_set write_data_reg_10(.CP(n_63610), .D(n_28681), .SD(1'b1), .Q
		(write_data[10]));
	notech_mux2 i_12262(.S(n_31326), .A(write_data[10]), .B(n_20894), .Z(n_28681
		));
	notech_reg_set write_data_reg_11(.CP(n_63672), .D(n_28687), .SD(1'b1), .Q
		(write_data[11]));
	notech_mux2 i_12270(.S(n_31326), .A(write_data[11]), .B(n_20899), .Z(n_28687
		));
	notech_reg_set write_data_reg_12(.CP(n_63668), .D(n_28693), .SD(1'b1), .Q
		(write_data[12]));
	notech_mux2 i_12278(.S(n_31326), .A(write_data[12]), .B(n_20904), .Z(n_28693
		));
	notech_reg_set write_data_reg_13(.CP(n_63608), .D(n_28699), .SD(1'b1), .Q
		(write_data[13]));
	notech_mux2 i_12286(.S(n_31326), .A(write_data[13]), .B(n_20909), .Z(n_28699
		));
	notech_reg_set write_data_reg_14(.CP(n_63668), .D(n_28705), .SD(1'b1), .Q
		(write_data[14]));
	notech_mux2 i_12294(.S(n_31326), .A(write_data[14]), .B(n_20914), .Z(n_28705
		));
	notech_reg_set write_data_reg_15(.CP(n_63668), .D(n_28711), .SD(1'b1), .Q
		(write_data[15]));
	notech_mux2 i_12302(.S(n_31326), .A(write_data[15]), .B(n_20919), .Z(n_28711
		));
	notech_nand2 i_17263187(.A(tsc[1]), .B(n_30615), .Z(n_1661));
	notech_reg_set write_data_reg_16(.CP(n_63668), .D(n_28717), .SD(1'b1), .Q
		(write_data[16]));
	notech_mux2 i_12310(.S(n_55289), .A(write_data[16]), .B(n_20924), .Z(n_28717
		));
	notech_reg_set write_data_reg_17(.CP(n_63668), .D(n_28723), .SD(1'b1), .Q
		(write_data[17]));
	notech_mux2 i_12318(.S(n_55289), .A(write_data[17]), .B(n_20929), .Z(n_28723
		));
	notech_reg_set write_data_reg_18(.CP(n_63668), .D(n_28729), .SD(1'b1), .Q
		(write_data[18]));
	notech_mux2 i_12326(.S(n_55289), .A(write_data[18]), .B(n_20934), .Z(n_28729
		));
	notech_reg_set write_data_reg_19(.CP(n_63668), .D(n_28735), .SD(1'b1), .Q
		(write_data[19]));
	notech_mux2 i_12334(.S(n_55289), .A(write_data[19]), .B(n_20939), .Z(n_28735
		));
	notech_reg_set write_data_reg_20(.CP(n_63668), .D(n_28744), .SD(1'b1), .Q
		(write_data[20]));
	notech_mux2 i_12342(.S(n_55289), .A(write_data[20]), .B(n_20944), .Z(n_28744
		));
	notech_ao4 i_93862454(.A(n_63752), .B(n_61958), .C(n_61052), .D(n_28555)
		, .Z(n_165695997));
	notech_reg_set write_data_reg_21(.CP(n_63668), .D(n_28750), .SD(1'b1), .Q
		(write_data[21]));
	notech_mux2 i_12350(.S(n_55289), .A(write_data[21]), .B(n_20949), .Z(n_28750
		));
	notech_reg_set write_data_reg_22(.CP(n_63668), .D(n_28756), .SD(1'b1), .Q
		(write_data[22]));
	notech_mux2 i_12358(.S(n_55289), .A(write_data[22]), .B(n_20954), .Z(n_28756
		));
	notech_reg_set write_data_reg_23(.CP(n_63668), .D(n_28762), .SD(1'b1), .Q
		(write_data[23]));
	notech_mux2 i_12366(.S(n_55289), .A(write_data[23]), .B(n_20959), .Z(n_28762
		));
	notech_reg_set write_data_reg_24(.CP(n_63692), .D(n_28768), .SD(1'b1), .Q
		(write_data[24]));
	notech_mux2 i_12374(.S(n_55289), .A(write_data[24]), .B(n_20964), .Z(n_28768
		));
	notech_ao4 i_11663241(.A(n_60169), .B(n_58229), .C(n_30919), .D(n_30340)
		, .Z(n_165296001));
	notech_reg_set write_data_reg_25(.CP(n_63692), .D(n_28774), .SD(1'b1), .Q
		(write_data[25]));
	notech_mux2 i_12382(.S(n_55289), .A(write_data[25]), .B(n_20969), .Z(n_28774
		));
	notech_reg_set write_data_reg_26(.CP(n_63692), .D(n_28780), .SD(1'b1), .Q
		(write_data[26]));
	notech_mux2 i_12390(.S(n_55289), .A(write_data[26]), .B(n_20974), .Z(n_28780
		));
	notech_ao4 i_11763240(.A(n_60169), .B(n_59005), .C(n_30920), .D(n_30340)
		, .Z(n_165096003));
	notech_reg_set write_data_reg_27(.CP(n_63692), .D(n_28786), .SD(1'b1), .Q
		(write_data[27]));
	notech_mux2 i_12398(.S(n_55289), .A(write_data[27]), .B(n_20979), .Z(n_28786
		));
	notech_reg_set write_data_reg_28(.CP(n_63692), .D(n_28792), .SD(1'b1), .Q
		(write_data[28]));
	notech_mux2 i_12406(.S(n_55289), .A(write_data[28]), .B(n_20984), .Z(n_28792
		));
	notech_mux2 i_15663203(.S(n_32249), .A(n_165296001), .B(n_165096003), .Z
		(n_164896005));
	notech_reg_set write_data_reg_29(.CP(n_63692), .D(n_28798), .SD(1'b1), .Q
		(write_data[29]));
	notech_mux2 i_12414(.S(n_55289), .A(write_data[29]), .B(n_20989), .Z(n_28798
		));
	notech_reg_set write_data_reg_30(.CP(n_63692), .D(n_28804), .SD(1'b1), .Q
		(write_data[30]));
	notech_mux2 i_12422(.S(n_55289), .A(write_data[30]), .B(n_20994), .Z(n_28804
		));
	notech_reg_set write_data_reg_31(.CP(n_63692), .D(n_28810), .SD(1'b1), .Q
		(write_data[31]));
	notech_mux2 i_12430(.S(n_55289), .A(write_data[31]), .B(n_20999), .Z(n_28810
		));
	notech_reg ldtr_reg_0(.CP(n_63692), .D(n_28816), .CD(n_62402), .Q(ldtr[0
		]));
	notech_mux2 i_12438(.S(n_98290349), .A(opb[0]), .B(ldtr[0]), .Z(n_28816)
		);
	notech_and3 i_49063351(.A(n_171460318), .B(n_171660320), .C(n_171060314)
		, .Z(n_30274));
	notech_reg ldtr_reg_1(.CP(n_63692), .D(n_28822), .CD(n_62403), .Q(ldtr[1
		]));
	notech_mux2 i_12446(.S(n_98290349), .A(opb[1]), .B(ldtr[1]), .Z(n_28822)
		);
	notech_or4 i_99663361(.A(n_2383), .B(n_61757), .C(n_61766), .D(n_165695997
		), .Z(n_28554));
	notech_reg ldtr_reg_2(.CP(n_63692), .D(n_28828), .CD(n_62404), .Q(ldtr[2
		]));
	notech_mux2 i_12454(.S(n_98290349), .A(opb[2]), .B(ldtr[2]), .Z(n_28828)
		);
	notech_ao4 i_190964284(.A(n_32243), .B(n_163196017), .C(n_60188), .D(n_27378
		), .Z(n_164496008));
	notech_reg ldtr_reg_3(.CP(n_63692), .D(n_28834), .CD(n_62407), .Q(ldtr[3
		]));
	notech_mux2 i_12462(.S(n_98290349), .A(opb[3]), .B(ldtr[3]), .Z(n_28834)
		);
	notech_reg ldtr_reg_4(.CP(n_63692), .D(n_28840), .CD(n_62404), .Q(ldtr[4
		]));
	notech_mux2 i_12470(.S(n_98290349), .A(opb[4]), .B(ldtr[4]), .Z(n_28840)
		);
	notech_reg ldtr_reg_5(.CP(n_63692), .D(n_28846), .CD(n_62404), .Q(ldtr[5
		]));
	notech_mux2 i_12478(.S(n_98290349), .A(opb[5]), .B(ldtr[5]), .Z(n_28846)
		);
	notech_and3 i_30867(.A(n_61092), .B(n_61660), .C(n_33108), .Z(n_164196010
		));
	notech_reg ldtr_reg_6(.CP(n_63692), .D(n_28853), .CD(n_62407), .Q(ldtr[6
		]));
	notech_mux2 i_12486(.S(n_98290349), .A(opb[6]), .B(ldtr[6]), .Z(n_28853)
		);
	notech_and3 i_30869(.A(n_61092), .B(n_61660), .C(\eflags[10] ), .Z(n_1640
		));
	notech_reg ldtr_reg_7(.CP(n_63692), .D(n_28862), .CD(n_62407), .Q(ldtr[7
		]));
	notech_mux2 i_12494(.S(n_98290349), .A(opb[7]), .B(ldtr[7]), .Z(n_28862)
		);
	notech_reg ldtr_reg_8(.CP(n_63692), .D(n_28871), .CD(n_62407), .Q(ldtr[8
		]));
	notech_mux2 i_12502(.S(n_98290349), .A(opb[8]), .B(ldtr[8]), .Z(n_28871)
		);
	notech_reg ldtr_reg_9(.CP(n_63692), .D(n_28878), .CD(n_62407), .Q(ldtr[9
		]));
	notech_mux2 i_12512(.S(n_98290349), .A(opb[9]), .B(ldtr[9]), .Z(n_28878)
		);
	notech_reg ldtr_reg_10(.CP(n_63668), .D(n_28884), .CD(n_62407), .Q(ldtr[
		10]));
	notech_mux2 i_12520(.S(n_98290349), .A(opb[10]), .B(ldtr[10]), .Z(n_28884
		));
	notech_reg ldtr_reg_11(.CP(n_63692), .D(n_28890), .CD(n_62404), .Q(ldtr[
		11]));
	notech_mux2 i_12528(.S(n_98290349), .A(opb[11]), .B(ldtr[11]), .Z(n_28890
		));
	notech_reg ldtr_reg_12(.CP(n_63670), .D(n_28896), .CD(n_62404), .Q(ldtr[
		12]));
	notech_mux2 i_12536(.S(n_98290349), .A(opb[12]), .B(ldtr[12]), .Z(n_28896
		));
	notech_ao3 i_100565163(.A(n_328160909), .B(n_26624), .C(n_276460613), .Z
		(n_1634));
	notech_reg ldtr_reg_13(.CP(n_63670), .D(n_28902), .CD(n_62404), .Q(ldtr[
		13]));
	notech_mux2 i_12544(.S(n_98290349), .A(opb[13]), .B(ldtr[13]), .Z(n_28902
		));
	notech_nand2 i_100365165(.A(n_28551), .B(n_28552), .Z(n_163396015));
	notech_reg ldtr_reg_14(.CP(n_63670), .D(n_28908), .CD(n_62404), .Q(ldtr[
		14]));
	notech_mux2 i_12552(.S(n_98290349), .A(opb[14]), .B(ldtr[14]), .Z(n_28908
		));
	notech_ao4 i_99765171(.A(n_60169), .B(n_28533), .C(n_60188), .D(n_28007)
		, .Z(n_163296016));
	notech_reg ldtr_reg_15(.CP(n_63670), .D(n_28914), .CD(n_62404), .Q(ldtr[
		15]));
	notech_mux2 i_12560(.S(n_98290349), .A(opb[15]), .B(ldtr[15]), .Z(n_28914
		));
	notech_ao4 i_125066155(.A(n_63752), .B(n_61958), .C(n_61052), .D(n_27378
		), .Z(n_163196017));
	notech_reg ldtr_reg_16(.CP(n_63670), .D(n_28920), .CD(n_62404), .Q(ldtr[
		16]));
	notech_mux2 i_12568(.S(n_55495), .A(opb[16]), .B(ldtr[16]), .Z(n_28920)
		);
	notech_reg ldtr_reg_17(.CP(n_63670), .D(n_28926), .CD(n_62404), .Q(ldtr[
		17]));
	notech_mux2 i_12576(.S(n_55495), .A(opb[17]), .B(ldtr[17]), .Z(n_28926)
		);
	notech_reg ldtr_reg_18(.CP(n_63670), .D(n_28932), .CD(n_62404), .Q(ldtr[
		18]));
	notech_mux2 i_12584(.S(n_55495), .A(opb[18]), .B(ldtr[18]), .Z(n_28932)
		);
	notech_nand3 i_133967997(.A(n_162696022), .B(n_1563), .C(n_1564), .Z(n_162896020
		));
	notech_reg ldtr_reg_19(.CP(n_63670), .D(n_28938), .CD(n_62404), .Q(ldtr[
		19]));
	notech_mux2 i_12592(.S(n_55495), .A(opb[19]), .B(ldtr[19]), .Z(n_28938)
		);
	notech_reg ldtr_reg_20(.CP(n_63670), .D(n_28944), .CD(n_62404), .Q(ldtr[
		20]));
	notech_mux2 i_12600(.S(n_55495), .A(opb[20]), .B(ldtr[20]), .Z(n_28944)
		);
	notech_and4 i_133767999(.A(n_1560), .B(n_327860906), .C(n_1562), .D(n_1561
		), .Z(n_162696022));
	notech_reg ldtr_reg_21(.CP(n_63670), .D(n_28950), .CD(n_62415), .Q(ldtr[
		21]));
	notech_mux2 i_12608(.S(n_55495), .A(opb[21]), .B(ldtr[21]), .Z(n_28950)
		);
	notech_reg ldtr_reg_22(.CP(n_63670), .D(n_28956), .CD(n_62415), .Q(ldtr[
		22]));
	notech_mux2 i_12616(.S(n_55495), .A(opb[22]), .B(ldtr[22]), .Z(n_28956)
		);
	notech_reg ldtr_reg_23(.CP(n_63670), .D(n_28962), .CD(n_62415), .Q(ldtr[
		23]));
	notech_mux2 i_12624(.S(n_55495), .A(opb[23]), .B(ldtr[23]), .Z(n_28962)
		);
	notech_reg ldtr_reg_24(.CP(n_63670), .D(n_28968), .CD(n_62415), .Q(ldtr[
		24]));
	notech_mux2 i_12632(.S(n_55495), .A(opb[24]), .B(ldtr[24]), .Z(n_28968)
		);
	notech_reg ldtr_reg_25(.CP(n_63670), .D(n_28974), .CD(n_62415), .Q(ldtr[
		25]));
	notech_mux2 i_12640(.S(n_55495), .A(opb[25]), .B(ldtr[25]), .Z(n_28974)
		);
	notech_reg ldtr_reg_26(.CP(n_63670), .D(n_28980), .CD(n_62415), .Q(ldtr[
		26]));
	notech_mux2 i_12648(.S(n_55495), .A(opb[26]), .B(ldtr[26]), .Z(n_28980)
		);
	notech_ao3 i_123868088(.A(n_1553), .B(n_1554), .C(n_1618), .Z(n_1620));
	notech_reg ldtr_reg_27(.CP(n_63670), .D(n_28987), .CD(n_62415), .Q(ldtr[
		27]));
	notech_mux2 i_12656(.S(n_55495), .A(opb[27]), .B(ldtr[27]), .Z(n_28987)
		);
	notech_reg ldtr_reg_28(.CP(n_63670), .D(n_28999), .CD(n_62415), .Q(ldtr[
		28]));
	notech_mux2 i_12664(.S(n_55495), .A(opb[28]), .B(ldtr[28]), .Z(n_28999)
		);
	notech_or4 i_123668090(.A(n_1550), .B(n_1551), .C(n_1552), .D(n_1615), .Z
		(n_1618));
	notech_reg ldtr_reg_29(.CP(n_63670), .D(n_29005), .CD(n_62415), .Q(ldtr[
		29]));
	notech_mux2 i_12672(.S(n_55495), .A(opb[29]), .B(ldtr[29]), .Z(n_29005)
		);
	notech_reg ldtr_reg_30(.CP(n_63670), .D(n_29011), .CD(n_62415), .Q(ldtr[
		30]));
	notech_mux2 i_12680(.S(n_55495), .A(opb[30]), .B(ldtr[30]), .Z(n_29011)
		);
	notech_reg ldtr_reg_31(.CP(n_63608), .D(n_29017), .CD(n_62414), .Q(ldtr[
		31]));
	notech_mux2 i_12688(.S(n_55495), .A(n_60629), .B(ldtr[31]), .Z(n_29017)
		);
	notech_or4 i_123368093(.A(n_30917), .B(n_1548), .C(n_1549), .D(n_154796026
		), .Z(n_1615));
	notech_reg gdtr_reg_0(.CP(n_63608), .D(n_29023), .CD(n_62414), .Q(gdtr[0
		]));
	notech_mux2 i_12696(.S(n_98390350), .A(opb[0]), .B(gdtr[0]), .Z(n_29023)
		);
	notech_reg gdtr_reg_1(.CP(n_63608), .D(n_29029), .CD(n_62414), .Q(gdtr[1
		]));
	notech_mux2 i_12704(.S(n_98390350), .A(opb[1]), .B(gdtr[1]), .Z(n_29029)
		);
	notech_reg gdtr_reg_2(.CP(n_63608), .D(n_29035), .CD(n_62414), .Q(gdtr[2
		]));
	notech_mux2 i_12712(.S(n_98390350), .A(opb[2]), .B(gdtr[2]), .Z(n_29035)
		);
	notech_reg gdtr_reg_3(.CP(n_63608), .D(n_29041), .CD(n_62414), .Q(gdtr[3
		]));
	notech_mux2 i_12720(.S(n_98390350), .A(opb[3]), .B(gdtr[3]), .Z(n_29041)
		);
	notech_or4 i_60668684(.A(n_1540), .B(n_1608), .C(n_1541), .D(n_1544), .Z
		(n_1611));
	notech_reg gdtr_reg_4(.CP(n_63608), .D(n_29047), .CD(n_62414), .Q(gdtr[4
		]));
	notech_mux2 i_12728(.S(n_98390350), .A(opb[4]), .B(gdtr[4]), .Z(n_29047)
		);
	notech_reg gdtr_reg_5(.CP(n_63608), .D(n_29053), .CD(n_62414), .Q(gdtr[5
		]));
	notech_mux2 i_12736(.S(n_98390350), .A(opb[5]), .B(gdtr[5]), .Z(n_29053)
		);
	notech_reg gdtr_reg_6(.CP(n_63608), .D(n_29059), .CD(n_62414), .Q(gdtr[6
		]));
	notech_mux2 i_12744(.S(n_98390350), .A(opb[6]), .B(gdtr[6]), .Z(n_29059)
		);
	notech_or4 i_60268688(.A(n_1537), .B(n_1605), .C(n_1538), .D(n_1539), .Z
		(n_1608));
	notech_reg gdtr_reg_7(.CP(n_63608), .D(n_29065), .CD(n_62414), .Q(gdtr[7
		]));
	notech_mux2 i_12752(.S(n_98390350), .A(opb[7]), .B(gdtr[7]), .Z(n_29065)
		);
	notech_reg gdtr_reg_8(.CP(n_63528), .D(n_29071), .CD(n_62418), .Q(gdtr[8
		]));
	notech_mux2 i_12760(.S(n_98390350), .A(opb[8]), .B(gdtr[8]), .Z(n_29071)
		);
	notech_reg gdtr_reg_9(.CP(n_63608), .D(n_29077), .CD(n_62418), .Q(gdtr[9
		]));
	notech_mux2 i_12768(.S(n_98390350), .A(opb[9]), .B(gdtr[9]), .Z(n_29077)
		);
	notech_or4 i_59968691(.A(n_1536), .B(n_1534), .C(n_30634), .D(n_1535), .Z
		(n_1605));
	notech_reg gdtr_reg_10(.CP(n_63614), .D(n_29086), .CD(n_62418), .Q(gdtr[
		10]));
	notech_mux2 i_12776(.S(n_98390350), .A(opb[10]), .B(gdtr[10]), .Z(n_29086
		));
	notech_reg gdtr_reg_11(.CP(n_63530), .D(n_29092), .CD(n_62418), .Q(gdtr[
		11]));
	notech_mux2 i_12784(.S(n_98390350), .A(opb[11]), .B(gdtr[11]), .Z(n_29092
		));
	notech_reg gdtr_reg_12(.CP(n_63530), .D(n_29098), .CD(n_62418), .Q(gdtr[
		12]));
	notech_mux2 i_12792(.S(n_98390350), .A(opb[12]), .B(gdtr[12]), .Z(n_29098
		));
	notech_ao4 i_60568685(.A(n_326760895), .B(n_30002), .C(n_326660894), .D(n_30001
		), .Z(n_1602));
	notech_reg gdtr_reg_13(.CP(n_63530), .D(n_29104), .CD(n_62419), .Q(gdtr[
		13]));
	notech_mux2 i_12800(.S(n_98390350), .A(opb[13]), .B(gdtr[13]), .Z(n_29104
		));
	notech_reg gdtr_reg_14(.CP(n_63530), .D(n_29110), .CD(n_62419), .Q(gdtr[
		14]));
	notech_mux2 i_12808(.S(n_98390350), .A(opb[14]), .B(gdtr[14]), .Z(n_29110
		));
	notech_or4 i_58268708(.A(n_1526), .B(n_1597), .C(n_1527), .D(n_1530), .Z
		(n_1600));
	notech_reg gdtr_reg_15(.CP(n_63530), .D(n_29116), .CD(n_62418), .Q(gdtr[
		15]));
	notech_mux2 i_12816(.S(n_98390350), .A(opb[15]), .B(gdtr[15]), .Z(n_29116
		));
	notech_reg gdtr_reg_16(.CP(n_63530), .D(n_29122), .CD(n_62419), .Q(gdtr[
		16]));
	notech_mux2 i_12824(.S(n_55657), .A(opb[16]), .B(gdtr[16]), .Z(n_29122)
		);
	notech_reg gdtr_reg_17(.CP(n_63530), .D(n_29128), .CD(n_62418), .Q(gdtr[
		17]));
	notech_mux2 i_12832(.S(n_55657), .A(opb[17]), .B(gdtr[17]), .Z(n_29128)
		);
	notech_or4 i_57868712(.A(n_1523), .B(n_1594), .C(n_1524), .D(n_1525), .Z
		(n_1597));
	notech_reg gdtr_reg_18(.CP(n_63530), .D(n_29134), .CD(n_62415), .Q(gdtr[
		18]));
	notech_mux2 i_12840(.S(n_55657), .A(opb[18]), .B(gdtr[18]), .Z(n_29134)
		);
	notech_reg gdtr_reg_19(.CP(n_63530), .D(n_29140), .CD(n_62418), .Q(gdtr[
		19]));
	notech_mux2 i_12848(.S(n_55657), .A(opb[19]), .B(gdtr[19]), .Z(n_29140)
		);
	notech_reg gdtr_reg_20(.CP(n_63616), .D(n_29146), .CD(n_62415), .Q(gdtr[
		20]));
	notech_mux2 i_12856(.S(n_55657), .A(opb[20]), .B(gdtr[20]), .Z(n_29146)
		);
	notech_or4 i_57468715(.A(n_1522), .B(n_1520), .C(n_1521), .D(n_30299), .Z
		(n_1594));
	notech_reg gdtr_reg_21(.CP(n_63616), .D(n_29152), .CD(n_62415), .Q(gdtr[
		21]));
	notech_mux2 i_12864(.S(n_55657), .A(opb[21]), .B(gdtr[21]), .Z(n_29152)
		);
	notech_reg gdtr_reg_22(.CP(n_63616), .D(n_29158), .CD(n_62418), .Q(gdtr[
		22]));
	notech_mux2 i_12873(.S(n_55657), .A(opb[22]), .B(gdtr[22]), .Z(n_29158)
		);
	notech_reg gdtr_reg_23(.CP(n_63616), .D(n_29164), .CD(n_62418), .Q(gdtr[
		23]));
	notech_mux2 i_12881(.S(n_55657), .A(opb[23]), .B(gdtr[23]), .Z(n_29164)
		);
	notech_ao4 i_58168709(.A(n_325760885), .B(n_30002), .C(n_325660884), .D(n_30001
		), .Z(n_1591));
	notech_reg gdtr_reg_24(.CP(n_63616), .D(n_29170), .CD(n_62418), .Q(gdtr[
		24]));
	notech_mux2 i_12889(.S(n_55657), .A(opb[24]), .B(gdtr[24]), .Z(n_29170)
		);
	notech_reg gdtr_reg_25(.CP(n_63616), .D(n_29176), .CD(n_62418), .Q(gdtr[
		25]));
	notech_mux2 i_12897(.S(n_55657), .A(opb[25]), .B(gdtr[25]), .Z(n_29176)
		);
	notech_and4 i_55668732(.A(n_1513), .B(n_1586), .C(n_1514), .D(n_1517), .Z
		(n_1589));
	notech_reg gdtr_reg_26(.CP(n_63616), .D(n_29182), .CD(n_62418), .Q(gdtr[
		26]));
	notech_mux2 i_12905(.S(n_55657), .A(opb[26]), .B(gdtr[26]), .Z(n_29182)
		);
	notech_reg gdtr_reg_27(.CP(n_63616), .D(n_29188), .CD(n_62412), .Q(gdtr[
		27]));
	notech_mux2 i_12913(.S(n_55657), .A(opb[27]), .B(gdtr[27]), .Z(n_29188)
		);
	notech_reg gdtr_reg_28(.CP(n_63616), .D(n_29195), .CD(n_62412), .Q(gdtr[
		28]));
	notech_mux2 i_12921(.S(n_55657), .A(opb[28]), .B(gdtr[28]), .Z(n_29195)
		);
	notech_and4 i_55268736(.A(n_1510), .B(n_1512), .C(n_1511), .D(n_1583), .Z
		(n_1586));
	notech_reg gdtr_reg_29(.CP(n_63616), .D(n_29205), .CD(n_62412), .Q(gdtr[
		29]));
	notech_mux2 i_12929(.S(n_55657), .A(opb[29]), .B(gdtr[29]), .Z(n_29205)
		);
	notech_reg gdtr_reg_30(.CP(n_63616), .D(n_29211), .CD(n_62412), .Q(gdtr[
		30]));
	notech_mux2 i_12937(.S(n_55657), .A(opb[30]), .B(gdtr[30]), .Z(n_29211)
		);
	notech_reg gdtr_reg_31(.CP(n_63616), .D(n_29218), .CD(n_62412), .Q(gdtr[
		31]));
	notech_mux2 i_12945(.S(n_55657), .A(n_60629), .B(gdtr[31]), .Z(n_29218)
		);
	notech_and4 i_54968739(.A(n_1507), .B(n_324860876), .C(n_1508), .D(n_1509
		), .Z(n_1583));
	notech_reg Daddrgs_reg_0(.CP(n_63616), .D(n_17668), .CD(n_62412), .Q(Daddrgs
		[0]));
	notech_reg Daddrgs_reg_1(.CP(n_63616), .D(n_17675), .CD(n_62412), .Q(Daddrgs
		[1]));
	notech_reg Daddrgs_reg_2(.CP(n_63616), .D(n_17682), .CD(n_62412), .Q(Daddrgs
		[2]));
	notech_reg Daddrgs_reg_3(.CP(n_63616), .D(n_17689), .CD(n_62412), .Q(Daddrgs
		[3]));
	notech_reg Daddrgs_reg_4(.CP(n_63616), .D(n_17696), .CD(n_62412), .Q(Daddrgs
		[4]));
	notech_reg Daddrgs_reg_5(.CP(n_63616), .D(n_17703), .CD(n_62410), .Q(Daddrgs
		[5]));
	notech_reg Daddrgs_reg_6(.CP(n_63616), .D(n_17710), .CD(n_62410), .Q(Daddrgs
		[6]));
	notech_reg Daddrgs_reg_7(.CP(n_63674), .D(n_17717), .CD(n_62410), .Q(Daddrgs
		[7]));
	notech_reg Daddrgs_reg_8(.CP(n_63614), .D(n_17724), .CD(n_62410), .Q(Daddrgs
		[8]));
	notech_reg Daddrgs_reg_9(.CP(n_63674), .D(n_17731), .CD(n_62410), .Q(Daddrgs
		[9]));
	notech_reg Daddrgs_reg_10(.CP(n_63674), .D(n_17738), .CD(n_62410), .Q(Daddrgs
		[10]));
	notech_reg Daddrgs_reg_11(.CP(n_63674), .D(n_17745), .CD(n_62412), .Q(Daddrgs
		[11]));
	notech_reg Daddrgs_reg_12(.CP(n_63674), .D(n_17752), .CD(n_62410), .Q(Daddrgs
		[12]));
	notech_reg Daddrgs_reg_13(.CP(n_63674), .D(n_17759), .CD(n_62410), .Q(Daddrgs
		[13]));
	notech_reg Daddrgs_reg_14(.CP(n_63674), .D(n_17766), .CD(n_62413), .Q(Daddrgs
		[14]));
	notech_reg Daddrgs_reg_15(.CP(n_63674), .D(n_17773), .CD(n_62413), .Q(Daddrgs
		[15]));
	notech_reg Daddrgs_reg_16(.CP(n_63674), .D(n_17780), .CD(n_62413), .Q(Daddrgs
		[16]));
	notech_reg Daddrgs_reg_17(.CP(n_63674), .D(n_17787), .CD(n_62413), .Q(Daddrgs
		[17]));
	notech_reg Daddrgs_reg_18(.CP(n_63674), .D(n_17794), .CD(n_62413), .Q(Daddrgs
		[18]));
	notech_reg Daddrgs_reg_19(.CP(n_63674), .D(n_17801), .CD(n_62414), .Q(Daddrgs
		[19]));
	notech_reg Daddrgs_reg_20(.CP(n_63674), .D(n_17808), .CD(n_62414), .Q(Daddrgs
		[20]));
	notech_reg Daddrgs_reg_21(.CP(n_63674), .D(n_17815), .CD(n_62414), .Q(Daddrgs
		[21]));
	notech_reg Daddrgs_reg_22(.CP(n_63674), .D(n_17822), .CD(n_62414), .Q(Daddrgs
		[22]));
	notech_reg Daddrgs_reg_23(.CP(n_63674), .D(n_17829), .CD(n_62413), .Q(Daddrgs
		[23]));
	notech_reg Daddrgs_reg_24(.CP(n_63674), .D(n_17836), .CD(n_62413), .Q(Daddrgs
		[24]));
	notech_reg Daddrgs_reg_25(.CP(n_63674), .D(n_17843), .CD(n_62413), .Q(Daddrgs
		[25]));
	notech_reg Daddrgs_reg_26(.CP(n_63674), .D(n_17850), .CD(n_62412), .Q(Daddrgs
		[26]));
	notech_reg Daddrgs_reg_27(.CP(n_63614), .D(n_17857), .CD(n_62412), .Q(Daddrgs
		[27]));
	notech_reg Daddrgs_reg_28(.CP(n_63614), .D(n_17864), .CD(n_62413), .Q(Daddrgs
		[28]));
	notech_reg Daddrgs_reg_29(.CP(n_63614), .D(n_17871), .CD(n_62413), .Q(Daddrgs
		[29]));
	notech_reg Daddrgs_reg_30(.CP(n_63614), .D(n_17878), .CD(n_62413), .Q(Daddrgs
		[30]));
	notech_reg Daddrgs_reg_31(.CP(n_63614), .D(n_17885), .CD(n_62413), .Q(Daddrgs
		[31]));
	notech_reg idtr_reg_0(.CP(n_63614), .D(n_29293), .CD(n_62413), .Q(idtr[0
		]));
	notech_mux2 i_13081(.S(n_98490351), .A(opb[0]), .B(idtr[0]), .Z(n_29293)
		);
	notech_reg idtr_reg_1(.CP(n_63614), .D(n_29299), .CD(n_62390), .Q(idtr[1
		]));
	notech_mux2 i_13089(.S(n_98490351), .A(opb[1]), .B(idtr[1]), .Z(n_29299)
		);
	notech_reg idtr_reg_2(.CP(n_63614), .D(n_29305), .CD(n_62390), .Q(idtr[2
		]));
	notech_mux2 i_13097(.S(n_98490351), .A(opb[2]), .B(idtr[2]), .Z(n_29305)
		);
	notech_ao4 i_55568733(.A(n_324460872), .B(n_30002), .C(n_324260870), .D(n_30001
		), .Z(n_1580));
	notech_reg idtr_reg_3(.CP(n_63614), .D(n_29311), .CD(n_62390), .Q(idtr[3
		]));
	notech_mux2 i_13105(.S(n_98490351), .A(opb[3]), .B(idtr[3]), .Z(n_29311)
		);
	notech_reg idtr_reg_4(.CP(n_63530), .D(n_29317), .CD(n_62390), .Q(idtr[4
		]));
	notech_mux2 i_13113(.S(n_98490351), .A(opb[4]), .B(idtr[4]), .Z(n_29317)
		);
	notech_and4 i_33868942(.A(n_1503), .B(n_1569), .C(n_1500), .D(n_1575), .Z
		(n_1578));
	notech_reg idtr_reg_5(.CP(n_63530), .D(n_29323), .CD(n_62390), .Q(idtr[5
		]));
	notech_mux2 i_13121(.S(n_98490351), .A(opb[5]), .B(idtr[5]), .Z(n_29323)
		);
	notech_reg idtr_reg_6(.CP(n_63618), .D(n_29329), .CD(n_62390), .Q(idtr[6
		]));
	notech_mux2 i_13129(.S(n_98490351), .A(opb[6]), .B(idtr[6]), .Z(n_29329)
		);
	notech_reg idtr_reg_7(.CP(n_63532), .D(n_29339), .CD(n_62391), .Q(idtr[7
		]));
	notech_mux2 i_13137(.S(n_98490351), .A(opb[7]), .B(idtr[7]), .Z(n_29339)
		);
	notech_and4 i_33468946(.A(n_1497), .B(n_1499), .C(n_1572), .D(n_1498), .Z
		(n_1575));
	notech_reg idtr_reg_8(.CP(n_63532), .D(n_29348), .CD(n_62390), .Q(idtr[8
		]));
	notech_mux2 i_13145(.S(n_98490351), .A(opb[8]), .B(idtr[8]), .Z(n_29348)
		);
	notech_reg idtr_reg_9(.CP(n_63532), .D(n_29354), .CD(n_62390), .Q(idtr[9
		]));
	notech_mux2 i_13153(.S(n_98490351), .A(opb[9]), .B(idtr[9]), .Z(n_29354)
		);
	notech_reg idtr_reg_10(.CP(n_63532), .D(n_29360), .CD(n_62390), .Q(idtr[
		10]));
	notech_mux2 i_13161(.S(n_98490351), .A(opb[10]), .B(idtr[10]), .Z(n_29360
		));
	notech_and3 i_33168949(.A(n_324860876), .B(n_1571), .C(n_1494), .Z(n_1572
		));
	notech_reg idtr_reg_11(.CP(n_63532), .D(n_29366), .CD(n_62389), .Q(idtr[
		11]));
	notech_mux2 i_13169(.S(n_98490351), .A(opb[11]), .B(idtr[11]), .Z(n_29366
		));
	notech_ao4 i_33068950(.A(n_323960867), .B(n_33165), .C(n_100242443), .D(n_323860866
		), .Z(n_1571));
	notech_reg idtr_reg_12(.CP(n_63532), .D(n_29372), .CD(n_62389), .Q(idtr[
		12]));
	notech_mux2 i_13177(.S(n_98490351), .A(opb[12]), .B(idtr[12]), .Z(n_29372
		));
	notech_reg idtr_reg_13(.CP(n_63532), .D(n_29378), .CD(n_62389), .Q(idtr[
		13]));
	notech_mux2 i_13185(.S(n_98490351), .A(opb[13]), .B(idtr[13]), .Z(n_29378
		));
	notech_ao4 i_33668944(.A(n_30391), .B(n_324560873), .C(n_30390), .D(n_324460872
		), .Z(n_1569));
	notech_reg idtr_reg_14(.CP(n_63532), .D(n_29384), .CD(n_62389), .Q(idtr[
		14]));
	notech_mux2 i_13193(.S(n_98490351), .A(opb[14]), .B(idtr[14]), .Z(n_29384
		));
	notech_ao4 i_1069253(.A(n_63698), .B(n_63736), .C(n_60188), .D(n_30212),
		 .Z(n_1568));
	notech_reg idtr_reg_15(.CP(n_63532), .D(n_29390), .CD(n_62389), .Q(idtr[
		15]));
	notech_mux2 i_13201(.S(n_98490351), .A(opb[15]), .B(idtr[15]), .Z(n_29390
		));
	notech_or4 i_121599(.A(n_1565), .B(n_162896020), .C(n_1566), .D(n_1558),
		 .Z(n_1567));
	notech_reg idtr_reg_16(.CP(n_63618), .D(n_29396), .CD(n_62390), .Q(idtr[
		16]));
	notech_mux2 i_13209(.S(n_55646), .A(opb[16]), .B(idtr[16]), .Z(n_29396)
		);
	notech_and2 i_133368003(.A(opb[0]), .B(n_1557), .Z(n_1566));
	notech_reg idtr_reg_17(.CP(n_63618), .D(n_29402), .CD(n_62390), .Q(idtr[
		17]));
	notech_mux2 i_13217(.S(n_55646), .A(opb[17]), .B(idtr[17]), .Z(n_29402)
		);
	notech_nor2 i_133068006(.A(n_3118), .B(n_33169), .Z(n_1565));
	notech_reg idtr_reg_18(.CP(n_63618), .D(n_29408), .CD(n_62389), .Q(idtr[
		18]));
	notech_mux2 i_13225(.S(n_55646), .A(opb[18]), .B(idtr[18]), .Z(n_29408)
		);
	notech_or2 i_132968007(.A(n_26942), .B(n_101142452), .Z(n_1564));
	notech_reg idtr_reg_19(.CP(n_63618), .D(n_29414), .CD(n_62390), .Q(idtr[
		19]));
	notech_mux2 i_13233(.S(n_55646), .A(opb[19]), .B(idtr[19]), .Z(n_29414)
		);
	notech_nao3 i_133168005(.A(n_63752), .B(opc[0]), .C(n_3111), .Z(n_1563)
		);
	notech_reg idtr_reg_20(.CP(n_63618), .D(n_29424), .CD(n_62392), .Q(idtr[
		20]));
	notech_mux2 i_13241(.S(n_55646), .A(opb[20]), .B(idtr[20]), .Z(n_29424)
		);
	notech_nao3 i_133268004(.A(n_63752), .B(opc_10[0]), .C(n_3117), .Z(n_1562
		));
	notech_reg idtr_reg_21(.CP(n_63618), .D(n_29430), .CD(n_62392), .Q(idtr[
		21]));
	notech_mux2 i_13249(.S(n_55646), .A(opb[21]), .B(idtr[21]), .Z(n_29430)
		);
	notech_nand2 i_132868008(.A(n_30665), .B(opd[0]), .Z(n_1561));
	notech_reg idtr_reg_22(.CP(n_63618), .D(n_29436), .CD(n_62391), .Q(idtr[
		22]));
	notech_mux2 i_13257(.S(n_55646), .A(opb[22]), .B(idtr[22]), .Z(n_29436)
		);
	notech_or2 i_132768009(.A(n_57086), .B(n_327560903), .Z(n_1560));
	notech_reg idtr_reg_23(.CP(n_63618), .D(n_29442), .CD(n_62392), .Q(idtr[
		23]));
	notech_mux2 i_13265(.S(n_55646), .A(opb[23]), .B(idtr[23]), .Z(n_29442)
		);
	notech_nand3 i_132668010(.A(n_302744461), .B(n_301744451), .C(n_26935), 
		.Z(n_1559));
	notech_reg idtr_reg_24(.CP(n_63618), .D(n_29448), .CD(n_62392), .Q(idtr[
		24]));
	notech_mux2 i_13273(.S(n_55646), .A(opb[24]), .B(idtr[24]), .Z(n_29448)
		);
	notech_and2 i_133468002(.A(opa[0]), .B(n_1559), .Z(n_1558));
	notech_reg idtr_reg_25(.CP(n_63618), .D(n_29454), .CD(n_62392), .Q(idtr[
		25]));
	notech_mux2 i_13281(.S(n_55646), .A(opb[25]), .B(idtr[25]), .Z(n_29454)
		);
	notech_nand3 i_132468012(.A(n_301844452), .B(n_302844462), .C(n_26940), 
		.Z(n_1557));
	notech_reg idtr_reg_26(.CP(n_63618), .D(n_29460), .CD(n_62392), .Q(idtr[
		26]));
	notech_mux2 i_13289(.S(n_55646), .A(opb[26]), .B(idtr[26]), .Z(n_29460)
		);
	notech_nand3 i_1021608(.A(n_1555), .B(n_1620), .C(n_1546), .Z(n_1556));
	notech_reg idtr_reg_27(.CP(n_63618), .D(n_29466), .CD(n_62392), .Q(idtr[
		27]));
	notech_mux2 i_13297(.S(n_55646), .A(opb[27]), .B(idtr[27]), .Z(n_29466)
		);
	notech_or2 i_122768099(.A(n_26935), .B(n_33168), .Z(n_1555));
	notech_reg idtr_reg_28(.CP(n_63618), .D(n_29472), .CD(n_62392), .Q(idtr[
		28]));
	notech_mux2 i_13305(.S(n_55646), .A(opb[28]), .B(idtr[28]), .Z(n_29472)
		);
	notech_nand2 i_122568101(.A(opa[9]), .B(n_30522), .Z(n_1554));
	notech_reg idtr_reg_29(.CP(n_63618), .D(n_29478), .CD(n_62391), .Q(idtr[
		29]));
	notech_mux2 i_13313(.S(n_55646), .A(opb[29]), .B(idtr[29]), .Z(n_29478)
		);
	notech_or4 i_122668100(.A(n_162262654), .B(n_57406), .C(n_26951), .D(n_99942440
		), .Z(n_1553));
	notech_reg idtr_reg_30(.CP(n_63618), .D(n_29484), .CD(n_62391), .Q(idtr[
		30]));
	notech_mux2 i_13321(.S(n_55646), .A(opb[30]), .B(idtr[30]), .Z(n_29484)
		);
	notech_and3 i_122868098(.A(n_63752), .B(opc[9]), .C(n_26823), .Z(n_1552)
		);
	notech_reg idtr_reg_31(.CP(n_63618), .D(n_29490), .CD(n_62391), .Q(idtr[
		31]));
	notech_mux2 i_13329(.S(n_55646), .A(n_60629), .B(idtr[31]), .Z(n_29490)
		);
	notech_ao3 i_123068096(.A(n_61007), .B(n_26822), .C(n_60188), .Z(n_1551)
		);
	notech_reg tr_reg_3(.CP(n_63618), .D(n_29496), .CD(n_62391), .Q(\tr[3] )
		);
	notech_mux2 i_13337(.S(n_98590352), .A(opb[3]), .B(\tr[3] ), .Z(n_29496)
		);
	notech_nor2 i_122368103(.A(n_303844472), .B(n_327060898), .Z(n_1550));
	notech_reg tr_reg_4(.CP(n_63618), .D(n_29502), .CD(n_62391), .Q(\tr[4] )
		);
	notech_mux2 i_13345(.S(n_98590352), .A(opb[4]), .B(\tr[4] ), .Z(n_29502)
		);
	notech_ao3 i_122968097(.A(n_63752), .B(opc_10[9]), .C(n_26821), .Z(n_1549
		));
	notech_reg tr_reg_5(.CP(n_63532), .D(n_29508), .CD(n_62391), .Q(\tr[5] )
		);
	notech_mux2 i_13353(.S(n_98590352), .A(opb[5]), .B(\tr[5] ), .Z(n_29508)
		);
	notech_and2 i_122268104(.A(n_305144485), .B(opd[9]), .Z(n_1548));
	notech_reg tr_reg_6(.CP(n_63532), .D(n_29514), .CD(n_62391), .Q(\tr[6] )
		);
	notech_mux2 i_13361(.S(n_98590352), .A(opb[6]), .B(\tr[6] ), .Z(n_29514)
		);
	notech_nor2 i_122168105(.A(n_57081), .B(n_326960897), .Z(n_154796026));
	notech_reg tr_reg_7(.CP(n_63534), .D(n_29520), .CD(n_62391), .Q(\tr[7] )
		);
	notech_mux2 i_13369(.S(n_98590352), .A(opb[7]), .B(\tr[7] ), .Z(n_29520)
		);
	notech_nand2 i_122468102(.A(opb[9]), .B(n_30523), .Z(n_1546));
	notech_reg tr_reg_8(.CP(n_63534), .D(n_29526), .CD(n_62391), .Q(\tr[8] )
		);
	notech_mux2 i_13377(.S(n_98590352), .A(opb[8]), .B(\tr[8] ), .Z(n_29526)
		);
	notech_nao3 i_320833(.A(n_1602), .B(n_1533), .C(n_1611), .Z(n_1545));
	notech_reg tr_reg_9(.CP(n_63534), .D(n_29535), .CD(n_62391), .Q(\tr[9] )
		);
	notech_mux2 i_13385(.S(n_98590352), .A(opb[9]), .B(\tr[9] ), .Z(n_29535)
		);
	notech_ao3 i_59268698(.A(n_63752), .B(opc[2]), .C(n_29994), .Z(n_1544)
		);
	notech_reg tr_reg_10(.CP(n_63534), .D(n_29545), .CD(n_62386), .Q(\tr[10] 
		));
	notech_mux2 i_13393(.S(n_98590352), .A(opb[10]), .B(\tr[10] ), .Z(n_29545
		));
	notech_reg tr_reg_11(.CP(n_63534), .D(n_29556), .CD(n_62386), .Q(\tr[11] 
		));
	notech_mux2 i_13401(.S(n_98590352), .A(opb[11]), .B(\tr[11] ), .Z(n_29556
		));
	notech_reg tr_reg_12(.CP(n_63534), .D(n_29564), .CD(n_62386), .Q(\tr[12] 
		));
	notech_mux2 i_13409(.S(n_98590352), .A(opb[12]), .B(\tr[12] ), .Z(n_29564
		));
	notech_nor2 i_59068700(.A(n_100842449), .B(n_30196), .Z(n_1541));
	notech_reg tr_reg_13(.CP(n_63534), .D(n_29570), .CD(n_62386), .Q(\tr[13] 
		));
	notech_mux2 i_13417(.S(n_98590352), .A(opb[13]), .B(\tr[13] ), .Z(n_29570
		));
	notech_nor2 i_58868702(.A(n_1532), .B(n_326160889), .Z(n_1540));
	notech_reg tr_reg_14(.CP(n_63534), .D(n_29577), .CD(n_62386), .Q(\tr[14] 
		));
	notech_mux2 i_13425(.S(n_98590352), .A(opb[14]), .B(\tr[14] ), .Z(n_29577
		));
	notech_and4 i_59168699(.A(n_30212), .B(n_30483), .C(n_63736), .D(opc_10[
		2]), .Z(n_1539));
	notech_reg tr_reg_15(.CP(n_63534), .D(n_29585), .CD(n_62386), .Q(\tr[15] 
		));
	notech_mux2 i_13433(.S(n_98590352), .A(opb[15]), .B(\tr[15] ), .Z(n_29585
		));
	notech_nor2 i_58768703(.A(n_305244486), .B(n_58802), .Z(n_1538));
	notech_reg desc_reg_0(.CP(n_63534), .D(n_29591), .CD(n_62386), .Q(desc[0
		]));
	notech_mux2 i_13441(.S(n_336689251), .A(read_data[0]), .B(desc[0]), .Z(n_29591
		));
	notech_nor2 i_59468696(.A(n_326560893), .B(n_29998), .Z(n_1537));
	notech_reg desc_reg_1(.CP(n_63534), .D(n_29597), .CD(n_62386), .Q(desc[1
		]));
	notech_mux2 i_13449(.S(n_336689251), .A(read_data[1]), .B(desc[1]), .Z(n_29597
		));
	notech_ao3 i_59368697(.A(n_57500), .B(n_323560863), .C(n_326460892), .Z(n_1536
		));
	notech_reg desc_reg_2(.CP(n_63534), .D(n_29603), .CD(n_62386), .Q(desc[2
		]));
	notech_mux2 i_13457(.S(n_336689251), .A(read_data[2]), .B(desc[2]), .Z(n_29603
		));
	notech_nor2 i_58668704(.A(n_57117), .B(n_326060888), .Z(n_1535));
	notech_reg desc_reg_3(.CP(n_63534), .D(n_29609), .CD(n_62386), .Q(desc[3
		]));
	notech_mux2 i_13465(.S(n_336689251), .A(read_data[3]), .B(desc[3]), .Z(n_29609
		));
	notech_nor2 i_58568705(.A(n_325960887), .B(n_30576), .Z(n_1534));
	notech_reg desc_reg_4(.CP(n_63534), .D(n_29615), .CD(n_62385), .Q(desc[4
		]));
	notech_mux2 i_13473(.S(n_336689251), .A(read_data[4]), .B(desc[4]), .Z(n_29615
		));
	notech_nao3 i_58968701(.A(n_30483), .B(\opa_12[2] ), .C(n_304344477), .Z
		(n_1533));
	notech_reg desc_reg_5(.CP(n_63534), .D(n_29621), .CD(n_62385), .Q(desc[5
		]));
	notech_mux2 i_13481(.S(n_336689251), .A(read_data[5]), .B(desc[5]), .Z(n_29621
		));
	notech_nor2 i_81669353(.A(n_30077), .B(n_30428), .Z(n_1532));
	notech_reg desc_reg_6(.CP(n_63534), .D(n_29627), .CD(n_62385), .Q(desc[6
		]));
	notech_mux2 i_13489(.S(n_336689251), .A(read_data[6]), .B(desc[6]), .Z(n_29627
		));
	notech_nao3 i_720837(.A(n_1591), .B(n_1519), .C(n_1600), .Z(n_1531));
	notech_reg desc_reg_7(.CP(n_63534), .D(n_29633), .CD(n_62385), .Q(desc[7
		]));
	notech_mux2 i_13497(.S(n_336689251), .A(read_data[7]), .B(desc[7]), .Z(n_29633
		));
	notech_ao3 i_56668722(.A(n_63752), .B(opc[6]), .C(n_29994), .Z(n_1530)
		);
	notech_reg desc_reg_8(.CP(n_63534), .D(n_29639), .CD(n_62385), .Q(desc[8
		]));
	notech_mux2 i_13505(.S(n_336689251), .A(read_data[8]), .B(desc[8]), .Z(n_29639
		));
	notech_reg desc_reg_9(.CP(n_63534), .D(n_29645), .CD(n_62385), .Q(desc[9
		]));
	notech_mux2 i_13513(.S(n_336689251), .A(read_data[9]), .B(desc[9]), .Z(n_29645
		));
	notech_reg desc_reg_10(.CP(n_63468), .D(n_29651), .CD(n_62386), .Q(desc[
		10]));
	notech_mux2 i_13521(.S(n_336689251), .A(read_data[10]), .B(desc[10]), .Z
		(n_29651));
	notech_nor2 i_56468724(.A(n_100542446), .B(n_30196), .Z(n_1527));
	notech_reg desc_reg_11(.CP(n_63468), .D(n_29657), .CD(n_62385), .Q(desc[
		11]));
	notech_mux2 i_13529(.S(n_336689251), .A(read_data[11]), .B(desc[11]), .Z
		(n_29657));
	notech_nor2 i_56268726(.A(n_1532), .B(n_325160879), .Z(n_1526));
	notech_reg desc_reg_12(.CP(n_63468), .D(n_29663), .CD(n_62385), .Q(desc[
		12]));
	notech_mux2 i_13537(.S(n_336689251), .A(read_data[12]), .B(desc[12]), .Z
		(n_29663));
	notech_and4 i_56568723(.A(n_30212), .B(n_30483), .C(n_63736), .D(opc_10[
		6]), .Z(n_1525));
	notech_reg desc_reg_13(.CP(n_63468), .D(n_29669), .CD(n_62387), .Q(desc[
		13]));
	notech_mux2 i_13545(.S(n_58682), .A(read_data[13]), .B(desc[13]), .Z(n_29669
		));
	notech_nor2 i_56168727(.A(n_305244486), .B(n_31479), .Z(n_1524));
	notech_reg desc_reg_14(.CP(n_63468), .D(n_29675), .CD(n_62389), .Q(desc[
		14]));
	notech_mux2 i_13553(.S(n_58682), .A(read_data[14]), .B(desc[14]), .Z(n_29675
		));
	notech_nor2 i_56868720(.A(n_325560883), .B(n_29998), .Z(n_1523));
	notech_reg desc_reg_15(.CP(n_63468), .D(n_29685), .CD(n_62387), .Q(desc[
		15]));
	notech_mux2 i_13561(.S(n_58682), .A(read_data[15]), .B(desc[15]), .Z(n_29685
		));
	notech_ao3 i_56768721(.A(n_57500), .B(n_323560863), .C(n_325460882), .Z(n_1522
		));
	notech_reg desc_reg_16(.CP(n_63468), .D(n_29691), .CD(n_62387), .Q(desc[
		16]));
	notech_mux2 i_13569(.S(n_58682), .A(read_data[16]), .B(desc[16]), .Z(n_29691
		));
	notech_nor2 i_56068728(.A(n_57117), .B(n_325060878), .Z(n_1521));
	notech_reg desc_reg_17(.CP(n_63468), .D(n_29697), .CD(n_62389), .Q(desc[
		17]));
	notech_mux2 i_13577(.S(n_58682), .A(read_data[17]), .B(desc[17]), .Z(n_29697
		));
	notech_ao3 i_55968729(.A(opa[6]), .B(n_323560863), .C(n_60188), .Z(n_1520
		));
	notech_reg desc_reg_18(.CP(n_63468), .D(n_29703), .CD(n_62389), .Q(desc[
		18]));
	notech_mux2 i_13585(.S(n_58682), .A(read_data[18]), .B(desc[18]), .Z(n_29703
		));
	notech_nao3 i_56368725(.A(n_30483), .B(\opa_12[6] ), .C(n_304344477), .Z
		(n_1519));
	notech_reg desc_reg_19(.CP(n_63378), .D(n_29709), .CD(n_62389), .Q(desc[
		19]));
	notech_mux2 i_13593(.S(n_58682), .A(read_data[19]), .B(desc[19]), .Z(n_29709
		));
	notech_nand3 i_820838(.A(n_1589), .B(n_1580), .C(n_1506), .Z(n_1518));
	notech_reg desc_reg_20(.CP(n_63468), .D(n_29715), .CD(n_62389), .Q(desc[
		20]));
	notech_mux2 i_13601(.S(n_58682), .A(read_data[20]), .B(desc[20]), .Z(n_29715
		));
	notech_nao3 i_54268746(.A(n_63752), .B(opc[7]), .C(n_29994), .Z(n_1517)
		);
	notech_reg desc_reg_21(.CP(n_63566), .D(n_29721), .CD(n_62389), .Q(desc[
		21]));
	notech_mux2 i_13609(.S(n_58682), .A(read_data[21]), .B(desc[21]), .Z(n_29721
		));
	notech_reg desc_reg_22(.CP(n_63420), .D(n_29727), .CD(n_62387), .Q(desc[
		22]));
	notech_mux2 i_13617(.S(n_58682), .A(read_data[22]), .B(desc[22]), .Z(n_29727
		));
	notech_reg desc_reg_23(.CP(n_63420), .D(n_29733), .CD(n_62387), .Q(desc[
		23]));
	notech_mux2 i_13625(.S(n_58682), .A(read_data[23]), .B(desc[23]), .Z(n_29733
		));
	notech_or2 i_54068748(.A(n_100242443), .B(n_30196), .Z(n_1514));
	notech_reg desc_reg_24(.CP(n_63420), .D(n_29739), .CD(n_62387), .Q(desc[
		24]));
	notech_mux2 i_13633(.S(n_115087077), .A(read_data[24]), .B(desc[24]), .Z
		(n_29739));
	notech_or4 i_53868750(.A(n_63698), .B(n_1532), .C(\opcode[2] ), .D(n_58275
		), .Z(n_1513));
	notech_reg desc_reg_25(.CP(n_63494), .D(n_29745), .CD(n_62386), .Q(desc[
		25]));
	notech_mux2 i_13641(.S(n_115087077), .A(read_data[25]), .B(desc[25]), .Z
		(n_29745));
	notech_nao3 i_54168747(.A(n_30212), .B(n_30483), .C(n_324660874), .Z(n_1512
		));
	notech_reg desc_reg_26(.CP(n_63494), .D(n_29751), .CD(n_62387), .Q(desc[
		26]));
	notech_mux2 i_13649(.S(n_115087077), .A(read_data[26]), .B(desc[26]), .Z
		(n_29751));
	notech_or2 i_53768751(.A(n_305244486), .B(n_31480), .Z(n_1511));
	notech_reg desc_reg_27(.CP(n_63494), .D(n_29757), .CD(n_62387), .Q(desc[
		27]));
	notech_mux2 i_13657(.S(n_115087077), .A(read_data[27]), .B(desc[27]), .Z
		(n_29757));
	notech_or4 i_54468744(.A(n_61056), .B(n_57500), .C(n_30576), .D(\nbus_11290[7] 
		), .Z(n_1510));
	notech_reg desc_reg_28(.CP(n_63494), .D(n_29764), .CD(n_62387), .Q(desc[
		28]));
	notech_mux2 i_13665(.S(n_115087077), .A(read_data[28]), .B(desc[28]), .Z
		(n_29764));
	notech_or4 i_54368745(.A(n_61056), .B(n_58275), .C(n_32261), .D(n_30576)
		, .Z(n_1509));
	notech_reg desc_reg_29(.CP(n_63494), .D(n_29770), .CD(n_62387), .Q(desc[
		29]));
	notech_mux2 i_13673(.S(n_115087077), .A(read_data[29]), .B(desc[29]), .Z
		(n_29770));
	notech_or2 i_53668752(.A(n_323760865), .B(n_57112), .Z(n_1508));
	notech_reg desc_reg_30(.CP(n_63494), .D(n_29776), .CD(n_62387), .Q(desc[
		30]));
	notech_mux2 i_13681(.S(n_115087077), .A(read_data[30]), .B(desc[30]), .Z
		(n_29776));
	notech_or4 i_53568753(.A(n_30212), .B(n_1532), .C(n_60188), .D(n_58275),
		 .Z(n_1507));
	notech_reg desc_reg_31(.CP(n_63494), .D(n_29782), .CD(n_62387), .Q(desc[
		31]));
	notech_mux2 i_13689(.S(n_115087077), .A(read_data[31]), .B(desc[31]), .Z
		(n_29782));
	notech_nao3 i_53968749(.A(n_30483), .B(\opa_12[7] ), .C(n_304344477), .Z
		(n_1506));
	notech_reg Daddrs_reg_0(.CP(n_63494), .D(n_29788), .CD(n_62399), .Q(Daddr
		[0]));
	notech_mux2 i_13697(.S(\nbus_11353[0] ), .A(Daddr[0]), .B(n_20628), .Z(n_29788
		));
	notech_nao3 i_820742(.A(n_1504), .B(n_1578), .C(n_1493), .Z(n_1505));
	notech_reg Daddrs_reg_1(.CP(n_63494), .D(n_29794), .CD(n_62399), .Q(Daddr
		[1]));
	notech_mux2 i_13705(.S(\nbus_11353[0] ), .A(Daddr[1]), .B(n_20634), .Z(n_29794
		));
	notech_or2 i_32468956(.A(n_30387), .B(n_324360871), .Z(n_1504));
	notech_reg Daddrs_reg_2(.CP(n_63494), .D(n_29800), .CD(n_62399), .Q(Daddr
		[2]));
	notech_mux2 i_13713(.S(\nbus_11353[0] ), .A(Daddr[2]), .B(n_20640), .Z(n_29800
		));
	notech_or4 i_32268958(.A(n_55831), .B(n_303944473), .C(n_60188), .D(n_58275
		), .Z(n_1503));
	notech_reg Daddrs_reg_3(.CP(n_63494), .D(n_29806), .CD(n_62399), .Q(Daddr
		[3]));
	notech_mux2 i_13721(.S(\nbus_11353[0] ), .A(Daddr[3]), .B(n_20646), .Z(n_29806
		));
	notech_reg Daddrs_reg_4(.CP(n_63494), .D(n_29812), .CD(n_62399), .Q(Daddr
		[4]));
	notech_mux2 i_13729(.S(\nbus_11353[0] ), .A(Daddr[4]), .B(n_20652), .Z(n_29812
		));
	notech_reg Daddrs_reg_5(.CP(n_63494), .D(n_29818), .CD(n_62399), .Q(Daddr
		[5]));
	notech_mux2 i_13737(.S(\nbus_11353[0] ), .A(Daddr[5]), .B(n_20658), .Z(n_29818
		));
	notech_or4 i_32368957(.A(n_303944473), .B(n_60169), .C(n_32266), .D(n_58275
		), .Z(n_1500));
	notech_reg Daddrs_reg_6(.CP(n_63494), .D(n_29824), .CD(n_62401), .Q(Daddr
		[6]));
	notech_mux2 i_13745(.S(\nbus_11353[0] ), .A(Daddr[6]), .B(n_20664), .Z(n_29824
		));
	notech_or4 i_32168959(.A(n_63698), .B(n_303944473), .C(\opcode[2] ), .D(n_58275
		), .Z(n_1499));
	notech_reg Daddrs_reg_7(.CP(n_63494), .D(n_29830), .CD(n_62399), .Q(Daddr
		[7]));
	notech_mux2 i_13753(.S(\nbus_11353[0] ), .A(Daddr[7]), .B(n_20670), .Z(n_29830
		));
	notech_nand2 i_32068960(.A(n_30630), .B(opd[7]), .Z(n_1498));
	notech_reg Daddrs_reg_8(.CP(n_63494), .D(n_29836), .CD(n_62399), .Q(Daddr
		[8]));
	notech_mux2 i_13761(.S(\nbus_11353[0] ), .A(Daddr[8]), .B(n_20676), .Z(n_29836
		));
	notech_nao3 i_32768953(.A(n_55831), .B(n_30484), .C(n_324660874), .Z(n_1497
		));
	notech_reg Daddrs_reg_9(.CP(n_63494), .D(n_29842), .CD(n_62399), .Q(Daddr
		[9]));
	notech_mux2 i_13769(.S(\nbus_11353[0] ), .A(Daddr[9]), .B(n_20682), .Z(n_29842
		));
	notech_reg Daddrs_reg_10(.CP(n_63494), .D(n_29848), .CD(n_62398), .Q(Daddr
		[10]));
	notech_mux2 i_13777(.S(\nbus_11353[0] ), .A(Daddr[10]), .B(n_20688), .Z(n_29848
		));
	notech_reg Daddrs_reg_11(.CP(n_63494), .D(n_29854), .CD(n_62398), .Q(Daddr
		[11]));
	notech_mux2 i_13785(.S(\nbus_11353[0] ), .A(Daddr[11]), .B(n_20694), .Z(n_29854
		));
	notech_or2 i_31768963(.A(n_323760865), .B(n_57163), .Z(n_1494));
	notech_reg Daddrs_reg_12(.CP(n_63566), .D(n_29860), .CD(n_62398), .Q(Daddr
		[12]));
	notech_mux2 i_13793(.S(\nbus_11353[0] ), .A(Daddr[12]), .B(n_20700), .Z(n_29860
		));
	notech_ao3 i_32868952(.A(n_30395), .B(n_57512), .C(n_324760875), .Z(n_1493
		));
	notech_reg Daddrs_reg_13(.CP(n_63492), .D(n_29866), .CD(n_62398), .Q(Daddr
		[13]));
	notech_mux2 i_13801(.S(\nbus_11353[0] ), .A(Daddr[13]), .B(n_20706), .Z(n_29866
		));
	notech_nao3 i_13569129(.A(n_57406), .B(n_30662), .C(n_26949), .Z(n_1492)
		);
	notech_reg Daddrs_reg_14(.CP(n_63566), .D(n_29872), .CD(n_62398), .Q(Daddr
		[14]));
	notech_mux2 i_13809(.S(\nbus_11353[0] ), .A(Daddr[14]), .B(n_20712), .Z(n_29872
		));
	notech_nand2 i_10769156(.A(n_115442595), .B(n_32208), .Z(n_1491));
	notech_reg Daddrs_reg_15(.CP(n_63566), .D(n_29878), .CD(n_62399), .Q(Daddr
		[15]));
	notech_mux2 i_13817(.S(\nbus_11353[0] ), .A(Daddr[15]), .B(n_20718), .Z(n_29878
		));
	notech_nand2 i_10569158(.A(n_115942600), .B(n_125342694), .Z(n_1490));
	notech_reg Daddrs_reg_16(.CP(n_63566), .D(n_29884), .CD(n_62399), .Q(Daddr
		[16]));
	notech_mux2 i_13825(.S(n_56279), .A(Daddr[16]), .B(n_20724), .Z(n_29884)
		);
	notech_nand2 i_10369160(.A(n_115942600), .B(n_32220), .Z(n_1489));
	notech_reg Daddrs_reg_17(.CP(n_63566), .D(n_29894), .CD(n_62399), .Q(Daddr
		[17]));
	notech_mux2 i_13833(.S(n_56279), .A(Daddr[17]), .B(n_20730), .Z(n_29894)
		);
	notech_reg Daddrs_reg_18(.CP(n_63566), .D(n_29900), .CD(n_62399), .Q(Daddr
		[18]));
	notech_mux2 i_13841(.S(n_56279), .A(Daddr[18]), .B(n_20736), .Z(n_29900)
		);
	notech_reg Daddrs_reg_19(.CP(n_63566), .D(n_29907), .CD(n_62402), .Q(Daddr
		[19]));
	notech_mux2 i_13849(.S(n_56279), .A(Daddr[19]), .B(n_20742), .Z(n_29907)
		);
	notech_ao4 i_26069366(.A(n_57566), .B(n_57637), .C(n_125342694), .D(n_30316
		), .Z(n_1486));
	notech_reg Daddrs_reg_20(.CP(n_63566), .D(n_29913), .CD(n_62402), .Q(Daddr
		[20]));
	notech_mux2 i_13857(.S(n_56279), .A(Daddr[20]), .B(n_20748), .Z(n_29913)
		);
	notech_reg Daddrs_reg_21(.CP(n_63566), .D(n_29920), .CD(n_62401), .Q(Daddr
		[21]));
	notech_mux2 i_13865(.S(n_56279), .A(Daddr[21]), .B(n_20754), .Z(n_29920)
		);
	notech_or4 i_8569178(.A(n_61819), .B(n_57535), .C(n_57662), .D(n_125342694
		), .Z(n_1484));
	notech_reg Daddrs_reg_22(.CP(n_63566), .D(n_29926), .CD(n_62401), .Q(Daddr
		[22]));
	notech_mux2 i_13873(.S(n_56279), .A(Daddr[22]), .B(n_20760), .Z(n_29926)
		);
	notech_reg Daddrs_reg_23(.CP(n_63566), .D(n_29932), .CD(n_62402), .Q(Daddr
		[23]));
	notech_mux2 i_13881(.S(n_56279), .A(Daddr[23]), .B(n_20766), .Z(n_29932)
		);
	notech_reg Daddrs_reg_24(.CP(n_63566), .D(n_29938), .CD(n_62402), .Q(Daddr
		[24]));
	notech_mux2 i_13889(.S(n_56279), .A(Daddr[24]), .B(n_20772), .Z(n_29938)
		);
	notech_ao4 i_83869305(.A(n_63728), .B(n_61958), .C(n_61052), .D(n_30212)
		, .Z(n_1481));
	notech_reg Daddrs_reg_25(.CP(n_63566), .D(n_29944), .CD(n_62402), .Q(Daddr
		[25]));
	notech_mux2 i_13897(.S(n_56279), .A(Daddr[25]), .B(n_20778), .Z(n_29944)
		);
	notech_reg Daddrs_reg_26(.CP(n_63566), .D(n_29950), .CD(n_62402), .Q(Daddr
		[26]));
	notech_mux2 i_13905(.S(n_56279), .A(Daddr[26]), .B(n_20784), .Z(n_29950)
		);
	notech_reg Daddrs_reg_27(.CP(n_63566), .D(n_29956), .CD(n_62402), .Q(Daddr
		[27]));
	notech_mux2 i_13913(.S(n_56279), .A(Daddr[27]), .B(n_20790), .Z(n_29956)
		);
	notech_or4 i_28671693(.A(n_1453), .B(n_1454), .C(n_1452), .D(n_1475), .Z
		(n_1478));
	notech_reg Daddrs_reg_28(.CP(n_63566), .D(n_29962), .CD(n_62401), .Q(Daddr
		[28]));
	notech_mux2 i_13921(.S(n_56279), .A(Daddr[28]), .B(n_20796), .Z(n_29962)
		);
	notech_reg Daddrs_reg_29(.CP(n_63566), .D(n_29968), .CD(n_62401), .Q(Daddr
		[29]));
	notech_mux2 i_13929(.S(n_56279), .A(Daddr[29]), .B(n_20802), .Z(n_29968)
		);
	notech_reg Daddrs_reg_30(.CP(n_63566), .D(n_29974), .CD(n_62401), .Q(Daddr
		[30]));
	notech_mux2 i_13937(.S(n_56279), .A(Daddr[30]), .B(n_20808), .Z(n_29974)
		);
	notech_nand3 i_28371696(.A(n_1449), .B(n_1472), .C(n_1474), .Z(n_1475)
		);
	notech_reg Daddrs_reg_31(.CP(n_63420), .D(n_29980), .CD(n_62401), .Q(Daddr
		[31]));
	notech_mux2 i_13945(.S(n_56279), .A(Daddr[31]), .B(n_20814), .Z(n_29980)
		);
	notech_ao4 i_28271697(.A(n_30257), .B(n_2383), .C(n_30240), .D(n_322460852
		), .Z(n_1474));
	notech_reg read_req_reg(.CP(n_63492), .D(n_29986), .CD(n_62401), .Q(read_reqs
		));
	notech_mux2 i_13953(.S(n_18351), .A(read_reqs), .B(n_31360), .Z(n_29986)
		);
	notech_reg writeio_req_reg(.CP(n_63492), .D(n_29992), .CD(n_62401), .Q(writeio_req
		));
	notech_mux2 i_13961(.S(n_17446), .A(writeio_req), .B(n_61660), .Z(n_29992
		));
	notech_ao4 i_28071699(.A(n_61092), .B(n_30759), .C(n_59099), .D(n_114845640
		), .Z(n_1472));
	notech_reg flush_tlb_reg(.CP(n_63492), .D(n_30004), .CD(n_62401), .Q(flush_tlb
		));
	notech_mux2 i_13969(.S(n_31361), .A(flush_tlb), .B(n_61660), .Z(n_30004)
		);
	notech_or2 i_25571724(.A(n_322460852), .B(n_323260860), .Z(n_1471));
	notech_reg flush_Dtlb_reg(.CP(n_63420), .D(n_30010), .CD(n_62401), .Q(flush_Dtlb
		));
	notech_mux2 i_13977(.S(n_14262), .A(flush_Dtlb), .B(n_311392439), .Z(n_30010
		));
	notech_reg_set terms_reg(.CP(n_63492), .D(n_30016), .SD(n_62401), .Q(terminate
		));
	notech_mux2 i_13985(.S(n_11332), .A(terminate), .B(n_11335), .Z(n_30016)
		);
	notech_reg writeio_data_reg_0(.CP(n_63496), .D(n_30022), .CD(n_62401), .Q
		(writeio_data[0]));
	notech_mux2 i_13993(.S(n_113490501), .A(n_60953), .B(writeio_data[0]), .Z
		(n_30022));
	notech_reg writeio_data_reg_1(.CP(n_63448), .D(n_30028), .CD(n_62396), .Q
		(writeio_data[1]));
	notech_mux2 i_14001(.S(n_113490501), .A(opa[1]), .B(writeio_data[1]), .Z
		(n_30028));
	notech_ao4 i_25871721(.A(n_1466), .B(n_30922), .C(n_1465), .D(n_30921), 
		.Z(n_1467));
	notech_reg writeio_data_reg_2(.CP(n_63448), .D(n_30034), .CD(n_62396), .Q
		(writeio_data[2]));
	notech_mux2 i_14009(.S(n_113490501), .A(opa[2]), .B(writeio_data[2]), .Z
		(n_30034));
	notech_nao3 i_6271902(.A(instrc[89]), .B(n_322260850), .C(instrc[91]), .Z
		(n_1466));
	notech_reg writeio_data_reg_3(.CP(n_63448), .D(n_30040), .CD(n_62396), .Q
		(writeio_data[3]));
	notech_mux2 i_14017(.S(n_113490501), .A(opa[3]), .B(writeio_data[3]), .Z
		(n_30040));
	notech_nao3 i_6171903(.A(instrc[93]), .B(n_33141), .C(n_321960847), .Z(n_1465
		));
	notech_reg writeio_data_reg_4(.CP(n_63496), .D(n_30046), .CD(n_62396), .Q
		(writeio_data[4]));
	notech_mux2 i_14025(.S(n_113490501), .A(opa[4]), .B(writeio_data[4]), .Z
		(n_30046));
	notech_and4 i_4871916(.A(n_30829), .B(instrc[105]), .C(n_30869), .D(n_30785
		), .Z(n_1464));
	notech_reg writeio_data_reg_5(.CP(n_63496), .D(n_30052), .CD(n_62396), .Q
		(writeio_data[5]));
	notech_mux2 i_14033(.S(n_113490501), .A(opa[5]), .B(writeio_data[5]), .Z
		(n_30052));
	notech_reg writeio_data_reg_6(.CP(n_63496), .D(n_30058), .CD(n_62396), .Q
		(writeio_data[6]));
	notech_mux2 i_14041(.S(n_113490501), .A(n_60989), .B(writeio_data[6]), .Z
		(n_30058));
	notech_or2 i_4371921(.A(n_322060848), .B(n_33161), .Z(n_1462));
	notech_reg writeio_data_reg_7(.CP(n_63496), .D(n_30064), .CD(n_62397), .Q
		(writeio_data[7]));
	notech_mux2 i_14049(.S(n_113490501), .A(n_60998), .B(writeio_data[7]), .Z
		(n_30064));
	notech_reg writeio_data_reg_8(.CP(n_63496), .D(n_30070), .CD(n_62396), .Q
		(writeio_data[8]));
	notech_mux2 i_14057(.S(n_113490501), .A(opa[8]), .B(writeio_data[8]), .Z
		(n_30070));
	notech_or4 i_1771947(.A(n_32484), .B(n_30618), .C(n_30343), .D(n_61661),
		 .Z(n_1460));
	notech_reg writeio_data_reg_9(.CP(n_63496), .D(n_30080), .CD(n_62396), .Q
		(writeio_data[9]));
	notech_mux2 i_14065(.S(n_113490501), .A(n_61007), .B(writeio_data[9]), .Z
		(n_30080));
	notech_reg writeio_data_reg_10(.CP(n_63496), .D(n_30086), .CD(n_62396), 
		.Q(writeio_data[10]));
	notech_mux2 i_14073(.S(n_113490501), .A(opa[10]), .B(writeio_data[10]), 
		.Z(n_30086));
	notech_reg writeio_data_reg_11(.CP(n_63496), .D(n_30092), .CD(n_62392), 
		.Q(writeio_data[11]));
	notech_mux2 i_14081(.S(n_113490501), .A(opa[11]), .B(writeio_data[11]), 
		.Z(n_30092));
	notech_or4 i_51750(.A(n_1455), .B(n_1478), .C(n_1446), .D(n_1456), .Z(n_1457
		));
	notech_reg writeio_data_reg_12(.CP(n_63496), .D(n_30098), .CD(n_62392), 
		.Q(writeio_data[12]));
	notech_mux2 i_14089(.S(n_113490501), .A(n_61016), .B(writeio_data[12]), 
		.Z(n_30098));
	notech_and2 i_27871701(.A(n_59099), .B(n_33324), .Z(n_1456));
	notech_reg writeio_data_reg_13(.CP(n_63496), .D(n_30104), .CD(n_62392), 
		.Q(writeio_data[13]));
	notech_mux2 i_14097(.S(n_113490501), .A(n_61025), .B(writeio_data[13]), 
		.Z(n_30104));
	notech_and2 i_27671703(.A(n_241746909), .B(n_33325), .Z(n_1455));
	notech_reg writeio_data_reg_14(.CP(n_63496), .D(n_30110), .CD(n_62392), 
		.Q(writeio_data[14]));
	notech_mux2 i_14105(.S(n_113490501), .A(opa[14]), .B(writeio_data[14]), 
		.Z(n_30110));
	notech_and2 i_27471705(.A(n_241346905), .B(n_28555), .Z(n_1454));
	notech_reg writeio_data_reg_15(.CP(n_63496), .D(n_30116), .CD(n_62392), 
		.Q(writeio_data[15]));
	notech_mux2 i_14113(.S(n_113490501), .A(n_61034), .B(writeio_data[15]), 
		.Z(n_30116));
	notech_and4 i_27571704(.A(instrc[104]), .B(instrc[106]), .C(n_33157), .D
		(n_1464), .Z(n_1453));
	notech_reg writeio_data_reg_16(.CP(n_63496), .D(n_30122), .CD(n_62396), 
		.Q(writeio_data[16]));
	notech_mux2 i_14121(.S(n_61043), .A(opa[16]), .B(writeio_data[16]), .Z(n_30122
		));
	notech_ao3 i_27771702(.A(n_63728), .B(n_28555), .C(n_1444), .Z(n_1452)
		);
	notech_reg writeio_data_reg_17(.CP(n_63496), .D(n_30128), .CD(n_62396), 
		.Q(writeio_data[17]));
	notech_mux2 i_14129(.S(n_61043), .A(opa[17]), .B(writeio_data[17]), .Z(n_30128
		));
	notech_reg writeio_data_reg_18(.CP(n_63448), .D(n_30134), .CD(n_62396), 
		.Q(writeio_data[18]));
	notech_mux2 i_14137(.S(n_61043), .A(opa[18]), .B(writeio_data[18]), .Z(n_30134
		));
	notech_reg writeio_data_reg_19(.CP(n_63496), .D(n_30140), .CD(n_62396), 
		.Q(writeio_data[19]));
	notech_mux2 i_14145(.S(n_61043), .A(opa[19]), .B(writeio_data[19]), .Z(n_30140
		));
	notech_nand3 i_27171708(.A(n_171160315), .B(n_61092), .C(n_61661), .Z(n_1449
		));
	notech_reg writeio_data_reg_20(.CP(n_63496), .D(n_30146), .CD(n_62398), 
		.Q(writeio_data[20]));
	notech_mux2 i_14153(.S(n_61043), .A(opa[20]), .B(writeio_data[20]), .Z(n_30146
		));
	notech_reg writeio_data_reg_21(.CP(n_63496), .D(n_30152), .CD(n_62398), 
		.Q(writeio_data[21]));
	notech_mux2 i_14161(.S(n_61043), .A(opa[21]), .B(writeio_data[21]), .Z(n_30152
		));
	notech_nao3 i_26971710(.A(n_1467), .B(n_144260310), .C(n_144160309), .Z(n_1447
		));
	notech_reg writeio_data_reg_22(.CP(n_63448), .D(n_30158), .CD(n_62397), 
		.Q(writeio_data[22]));
	notech_mux2 i_14169(.S(n_61043), .A(opa[22]), .B(writeio_data[22]), .Z(n_30158
		));
	notech_and4 i_27971700(.A(n_32481), .B(n_30869), .C(n_32353), .D(n_1447)
		, .Z(n_1446));
	notech_reg writeio_data_reg_23(.CP(n_63496), .D(n_30164), .CD(n_62398), 
		.Q(writeio_data[23]));
	notech_mux2 i_14177(.S(n_61043), .A(opa[23]), .B(writeio_data[23]), .Z(n_30164
		));
	notech_ao4 i_26171718(.A(n_114845640), .B(n_1443), .C(n_322560853), .D(n_30441
		), .Z(n_1445));
	notech_reg writeio_data_reg_24(.CP(n_63448), .D(n_30170), .CD(n_62398), 
		.Q(writeio_data[24]));
	notech_mux2 i_14185(.S(n_61043), .A(opa[24]), .B(writeio_data[24]), .Z(n_30170
		));
	notech_ao4 i_25671723(.A(n_57637), .B(n_2810), .C(n_30798), .D(n_32548),
		 .Z(n_1444));
	notech_reg writeio_data_reg_25(.CP(n_63448), .D(n_30176), .CD(n_62398), 
		.Q(writeio_data[25]));
	notech_mux2 i_14193(.S(n_61043), .A(opa[25]), .B(writeio_data[25]), .Z(n_30176
		));
	notech_ao4 i_2771937(.A(n_165695997), .B(n_57412), .C(n_30310), .D(n_1471
		), .Z(n_1443));
	notech_reg writeio_data_reg_26(.CP(n_63448), .D(n_30182), .CD(n_62398), 
		.Q(writeio_data[26]));
	notech_mux2 i_14201(.S(n_113490501), .A(opa[26]), .B(writeio_data[26]), 
		.Z(n_30182));
	notech_or4 i_26671713(.A(n_322660854), .B(n_33159), .C(instrc[99]), .D(n_33178
		), .Z(n_144260310));
	notech_reg writeio_data_reg_27(.CP(n_63448), .D(n_30188), .CD(n_62398), 
		.Q(writeio_data[27]));
	notech_mux2 i_14209(.S(n_61043), .A(opa[27]), .B(writeio_data[27]), .Z(n_30188
		));
	notech_ao3 i_26571714(.A(instrc[102]), .B(n_33142), .C(n_1462), .Z(n_144160309
		));
	notech_reg writeio_data_reg_28(.CP(n_63448), .D(n_30195), .CD(n_62398), 
		.Q(writeio_data[28]));
	notech_mux2 i_14217(.S(n_61043), .A(opa[28]), .B(writeio_data[28]), .Z(n_30195
		));
	notech_reg writeio_data_reg_29(.CP(n_63448), .D(n_30204), .CD(n_62397), 
		.Q(writeio_data[29]));
	notech_mux2 i_14225(.S(n_61043), .A(opa[29]), .B(writeio_data[29]), .Z(n_30204
		));
	notech_reg writeio_data_reg_30(.CP(n_63448), .D(n_30211), .CD(n_62397), 
		.Q(writeio_data[30]));
	notech_mux2 i_14233(.S(n_61043), .A(opa[30]), .B(writeio_data[30]), .Z(n_30211
		));
	notech_reg writeio_data_reg_31(.CP(n_63448), .D(n_30218), .CD(n_62397), 
		.Q(writeio_data[31]));
	notech_mux2 i_14241(.S(n_61043), .A(opa[31]), .B(writeio_data[31]), .Z(n_30218
		));
	notech_reg write_req_reg(.CP(n_63448), .D(n_30224), .CD(n_62397), .Q(write_reqs
		));
	notech_mux2 i_14249(.S(n_9187), .A(write_reqs), .B(n_31364), .Z(n_30224)
		);
	notech_reg pc_req_reg(.CP(n_63448), .D(n_30230), .CD(n_62397), .Q(pc_req
		));
	notech_mux2 i_14257(.S(n_8737), .A(pc_req), .B(n_61661), .Z(n_30230));
	notech_reg had_lgjmp_reg(.CP(n_63448), .D(n_30239), .CD(n_62397), .Q(had_lgjmp
		));
	notech_mux2 i_14265(.S(n_310992437), .A(\nbus_14542[31] ), .B(had_lgjmp)
		, .Z(n_30239));
	notech_and2 i_22515(.A(instrc[94]), .B(instrc[92]), .Z(n_143460302));
	notech_reg readio_req_reg(.CP(n_63448), .D(n_30246), .CD(n_62397), .Q(readio_req
		));
	notech_mux2 i_14273(.S(n_7488), .A(readio_req), .B(n_61661), .Z(n_30246)
		);
	notech_and2 i_22516(.A(instrc[90]), .B(instrc[88]), .Z(n_143360301));
	notech_reg write_sz_reg_0(.CP(n_63448), .D(n_30255), .CD(n_62397), .Q(write_sz
		[0]));
	notech_mux2 i_14281(.S(\nbus_11272[0] ), .A(write_sz[0]), .B(n_311292438
		), .Z(n_30255));
	notech_reg_set write_sz_reg_1(.CP(n_63448), .D(n_30262), .SD(n_62397), .Q
		(write_sz[1]));
	notech_mux2 i_14289(.S(\nbus_11272[0] ), .A(write_sz[1]), .B(n_31366), .Z
		(n_30262));
	notech_inv i_30315(.A(n_29557), .Z(n_30269));
	notech_inv i_30316(.A(n_27829), .Z(n_30270));
	notech_inv i_30320(.A(n_105014667), .Z(n_30271));
	notech_inv i_30321(.A(n_57887), .Z(n_30272));
	notech_inv i_30322(.A(n_57745), .Z(n_30273));
	notech_inv i_30323(.A(n_328360911), .Z(n_30275));
	notech_inv i_30324(.A(n_83839558), .Z(n_30276));
	notech_inv i_30325(.A(n_117276238), .Z(n_30277));
	notech_inv i_30326(.A(n_140576471), .Z(n_30278));
	notech_inv i_30327(.A(n_140776473), .Z(n_30279));
	notech_inv i_30328(.A(n_140976475), .Z(n_30281));
	notech_inv i_30329(.A(n_29560), .Z(n_30282));
	notech_inv i_30330(.A(n_386764398), .Z(n_30283));
	notech_inv i_30331(.A(n_216073528), .Z(n_30284));
	notech_inv i_30332(.A(n_212873496), .Z(n_30285));
	notech_inv i_30333(.A(n_170176767), .Z(n_30286));
	notech_inv i_30334(.A(n_1855), .Z(n_30287));
	notech_inv i_30335(.A(n_193776995), .Z(n_30288));
	notech_inv i_30336(.A(n_223277284), .Z(n_30289));
	notech_inv i_30337(.A(n_223977291), .Z(n_30290));
	notech_inv i_30338(.A(n_224677298), .Z(n_30291));
	notech_inv i_30339(.A(n_233777389), .Z(n_30292));
	notech_inv i_30340(.A(n_278577796), .Z(n_30293));
	notech_inv i_30341(.A(n_305978069), .Z(n_30294));
	notech_inv i_30342(.A(n_306678076), .Z(n_30295));
	notech_inv i_30343(.A(n_307378083), .Z(n_30296));
	notech_inv i_30344(.A(n_308078090), .Z(n_30297));
	notech_inv i_30345(.A(n_320678216), .Z(n_30298));
	notech_inv i_30346(.A(n_325860886), .Z(n_30299));
	notech_inv i_30347(.A(n_323578244), .Z(n_30300));
	notech_inv i_30348(.A(n_336678371), .Z(n_30301));
	notech_inv i_30349(.A(n_340378407), .Z(n_30302));
	notech_inv i_30351(.A(n_32520), .Z(n_30304));
	notech_inv i_30352(.A(n_32388), .Z(n_30305));
	notech_inv i_30353(.A(n_1852), .Z(n_30306));
	notech_inv i_30354(.A(n_19725), .Z(n_30307));
	notech_inv i_30355(.A(n_57501), .Z(n_30308));
	notech_inv i_30356(.A(n_32315), .Z(n_30309));
	notech_inv i_30357(.A(n_322360851), .Z(n_30310));
	notech_inv i_30358(.A(n_353378536), .Z(n_30311));
	notech_inv i_30359(.A(n_355078553), .Z(n_30312));
	notech_inv i_30360(.A(n_57385), .Z(n_30313));
	notech_inv i_30361(.A(n_24736), .Z(n_30314));
	notech_inv i_30362(.A(n_58279), .Z(n_30315));
	notech_inv i_30363(.A(n_57382), .Z(n_30316));
	notech_inv i_30364(.A(n_58058), .Z(n_30317));
	notech_inv i_30365(.A(n_193276990), .Z(n_30318));
	notech_inv i_30366(.A(n_29214), .Z(n_30319));
	notech_inv i_30367(.A(n_57129), .Z(n_30320));
	notech_inv i_30368(.A(n_63212389), .Z(n_30321));
	notech_inv i_30369(.A(n_57950), .Z(n_30322));
	notech_inv i_30370(.A(n_32508), .Z(n_30323));
	notech_inv i_30371(.A(n_19663), .Z(n_30324));
	notech_inv i_30372(.A(n_300322028), .Z(n_30325));
	notech_inv i_30373(.A(n_5680), .Z(n_30326));
	notech_inv i_30377(.A(n_32487), .Z(n_30330));
	notech_inv i_30378(.A(n_72012477), .Z(n_30331));
	notech_inv i_30379(.A(n_30864), .Z(n_30332));
	notech_inv i_30380(.A(n_30855), .Z(n_30333));
	notech_inv i_30381(.A(n_322260850), .Z(n_30334));
	notech_inv i_30382(.A(n_30829), .Z(n_30335));
	notech_inv i_30383(.A(n_19595), .Z(n_30336));
	notech_inv i_30385(.A(n_23763), .Z(n_30340));
	notech_inv i_30386(.A(n_63012387), .Z(n_30341));
	notech_inv i_30387(.A(n_56572), .Z(n_30342));
	notech_inv i_30388(.A(n_32481), .Z(n_30343));
	notech_inv i_30389(.A(n_379364324), .Z(n_30344));
	notech_inv i_30390(.A(n_317071143), .Z(n_30345));
	notech_inv i_30391(.A(n_313471111), .Z(n_30346));
	notech_inv i_30392(.A(n_223980740), .Z(n_30347));
	notech_inv i_30393(.A(n_235880859), .Z(n_30348));
	notech_inv i_30394(.A(n_236080861), .Z(n_30349));
	notech_inv i_30396(.A(n_333878344), .Z(n_30351));
	notech_inv i_30397(.A(n_271781206), .Z(n_30352));
	notech_inv i_30398(.A(n_271981208), .Z(n_30353));
	notech_inv i_30399(.A(n_441968003), .Z(n_30354));
	notech_inv i_30400(.A(n_61928), .Z(\opcode[2] ));
	notech_inv i_30401(.A(n_38705), .Z(n_30356));
	notech_inv i_30402(.A(n_338981856), .Z(n_30357));
	notech_inv i_30403(.A(n_19620), .Z(n_30358));
	notech_inv i_30404(.A(n_55975), .Z(n_30359));
	notech_inv i_30405(.A(n_384382274), .Z(n_30360));
	notech_inv i_30406(.A(n_396382340), .Z(n_30361));
	notech_inv i_30408(.A(n_32247), .Z(n_30363));
	notech_inv i_30410(.A(n_19548), .Z(n_30364));
	notech_inv i_30411(.A(n_4056), .Z(n_30365));
	notech_inv i_30412(.A(n_322960857), .Z(n_30366));
	notech_inv i_30414(.A(n_391364444), .Z(n_30367));
	notech_inv i_30415(.A(n_96629667), .Z(n_30368));
	notech_inv i_30416(.A(n_27798), .Z(n_30369));
	notech_inv i_30417(.A(n_414582401), .Z(n_30370));
	notech_inv i_30418(.A(n_309271075), .Z(n_30371));
	notech_inv i_30419(.A(n_56661), .Z(n_30372));
	notech_inv i_30420(.A(n_19637), .Z(n_30374));
	notech_inv i_30421(.A(n_4128), .Z(n_30375));
	notech_inv i_30422(.A(n_2081), .Z(n_30377));
	notech_inv i_30423(.A(n_347771364), .Z(n_30381));
	notech_inv i_30424(.A(n_347971365), .Z(n_30382));
	notech_inv i_30425(.A(n_59560), .Z(n_30383));
	notech_inv i_30426(.A(n_214080643), .Z(n_30384));
	notech_inv i_30427(.A(n_215180654), .Z(n_30385));
	notech_inv i_30428(.A(n_217580676), .Z(n_30388));
	notech_inv i_30429(.A(n_329360921), .Z(n_30389));
	notech_inv i_30430(.A(n_4375), .Z(n_30392));
	notech_inv i_30431(.A(n_4378), .Z(n_30396));
	notech_inv i_30432(.A(n_4380), .Z(n_30397));
	notech_inv i_30433(.A(n_4382), .Z(n_30398));
	notech_inv i_30434(.A(n_4383), .Z(n_30399));
	notech_inv i_30435(.A(n_4384), .Z(n_30400));
	notech_inv i_30436(.A(n_4386), .Z(n_30401));
	notech_inv i_30437(.A(n_4388), .Z(n_30402));
	notech_inv i_30438(.A(n_4389), .Z(n_30403));
	notech_inv i_30439(.A(n_4390), .Z(n_30404));
	notech_inv i_30440(.A(n_4392), .Z(n_30405));
	notech_inv i_30441(.A(n_4398), .Z(n_30406));
	notech_inv i_30442(.A(n_4399), .Z(n_30407));
	notech_inv i_30443(.A(\add_len_pc[2] ), .Z(n_30408));
	notech_inv i_30444(.A(\add_len_pc[3] ), .Z(n_30409));
	notech_inv i_30445(.A(\add_len_pc[4] ), .Z(n_30410));
	notech_inv i_30446(.A(n_4411), .Z(n_30411));
	notech_inv i_30447(.A(\add_len_pc[9] ), .Z(n_30412));
	notech_inv i_30448(.A(n_4430), .Z(n_30413));
	notech_inv i_30449(.A(n_1850), .Z(n_30414));
	notech_inv i_30450(.A(n_4434), .Z(n_30415));
	notech_inv i_30451(.A(n_56832), .Z(n_30416));
	notech_inv i_30452(.A(n_56904), .Z(n_30417));
	notech_inv i_30453(.A(n_383382264), .Z(n_30418));
	notech_inv i_30454(.A(n_446868052), .Z(n_30419));
	notech_inv i_30455(.A(n_342578429), .Z(n_30420));
	notech_inv i_30456(.A(n_4443), .Z(n_30421));
	notech_inv i_30457(.A(n_4446), .Z(n_30422));
	notech_inv i_30458(.A(n_446768051), .Z(n_30423));
	notech_inv i_30459(.A(n_4448), .Z(n_30424));
	notech_inv i_30460(.A(n_56930), .Z(n_30425));
	notech_inv i_30461(.A(n_30076), .Z(n_30426));
	notech_inv i_30462(.A(n_4454), .Z(n_30427));
	notech_inv i_30463(.A(n_30201), .Z(n_30428));
	notech_inv i_30464(.A(n_336860996), .Z(n_30429));
	notech_inv i_30465(.A(\add_len_pc[15] ), .Z(n_30430));
	notech_inv i_30466(.A(n_4463), .Z(n_30431));
	notech_inv i_30467(.A(\add_len_pc[12] ), .Z(n_30432));
	notech_inv i_30468(.A(\add_len_pc[11] ), .Z(n_30433));
	notech_inv i_30469(.A(n_4469), .Z(n_30434));
	notech_inv i_30471(.A(n_337060998), .Z(n_30436));
	notech_inv i_30472(.A(n_440967993), .Z(n_30437));
	notech_inv i_30473(.A(n_440767991), .Z(n_30438));
	notech_inv i_30474(.A(n_440467988), .Z(n_30439));
	notech_inv i_30475(.A(n_439867982), .Z(n_30440));
	notech_inv i_30476(.A(n_28555), .Z(n_30441));
	notech_inv i_30477(.A(n_439067974), .Z(n_30442));
	notech_inv i_30478(.A(n_438367967), .Z(n_30443));
	notech_inv i_30479(.A(n_438267966), .Z(n_30444));
	notech_inv i_30480(.A(n_438167965), .Z(n_30445));
	notech_inv i_30481(.A(n_135483810), .Z(n_30446));
	notech_inv i_30482(.A(n_188566312), .Z(n_30447));
	notech_inv i_30483(.A(n_171366155), .Z(n_30448));
	notech_inv i_30484(.A(n_436767951), .Z(n_30449));
	notech_inv i_30485(.A(n_436667950), .Z(n_30450));
	notech_inv i_30486(.A(n_139683852), .Z(n_30451));
	notech_inv i_30487(.A(n_139783853), .Z(n_30452));
	notech_inv i_30489(.A(n_142583881), .Z(n_30454));
	notech_inv i_30490(.A(n_142783883), .Z(n_30455));
	notech_inv i_30491(.A(n_153183987), .Z(n_30456));
	notech_inv i_30492(.A(n_170184157), .Z(n_30457));
	notech_inv i_30493(.A(n_427367857), .Z(n_30458));
	notech_inv i_30494(.A(n_171684168), .Z(n_30459));
	notech_inv i_30495(.A(n_172584175), .Z(n_30460));
	notech_inv i_30496(.A(n_176584199), .Z(n_30461));
	notech_inv i_30498(.A(n_195184378), .Z(n_30463));
	notech_inv i_30499(.A(n_215984579), .Z(n_30464));
	notech_inv i_30500(.A(n_217084590), .Z(n_30465));
	notech_inv i_30501(.A(n_218184601), .Z(n_30466));
	notech_inv i_30502(.A(n_218884608), .Z(n_30467));
	notech_inv i_30503(.A(n_219584615), .Z(n_30469));
	notech_inv i_30504(.A(n_220284622), .Z(n_30470));
	notech_inv i_30505(.A(n_220984629), .Z(n_30471));
	notech_inv i_30506(.A(n_223784657), .Z(n_30472));
	notech_inv i_30507(.A(n_32210), .Z(n_30473));
	notech_inv i_30508(.A(n_260885025), .Z(n_30475));
	notech_inv i_30509(.A(n_261985036), .Z(n_30476));
	notech_inv i_30510(.A(n_263085047), .Z(n_30477));
	notech_inv i_30511(.A(n_264185058), .Z(n_30478));
	notech_inv i_30512(.A(n_265285069), .Z(n_30479));
	notech_inv i_30513(.A(n_266085077), .Z(n_30480));
	notech_inv i_30514(.A(n_266885085), .Z(n_30481));
	notech_inv i_30515(.A(n_267685093), .Z(n_30482));
	notech_inv i_30516(.A(n_305844492), .Z(n_30483));
	notech_inv i_30517(.A(n_328060908), .Z(n_30484));
	notech_inv i_30518(.A(n_282185235), .Z(n_30485));
	notech_inv i_30519(.A(n_282385237), .Z(n_30486));
	notech_inv i_30520(.A(n_282585239), .Z(n_30487));
	notech_inv i_30521(.A(n_293485348), .Z(n_30488));
	notech_inv i_30522(.A(n_294585359), .Z(n_30489));
	notech_inv i_30524(.A(n_345785866), .Z(n_30491));
	notech_inv i_30525(.A(n_344785856), .Z(n_30492));
	notech_inv i_30527(.A(n_348285890), .Z(n_30494));
	notech_inv i_30528(.A(n_382764358), .Z(n_30495));
	notech_inv i_30529(.A(n_310267479), .Z(n_30497));
	notech_inv i_30532(.A(n_310167478), .Z(n_30498));
	notech_inv i_30533(.A(n_310067477), .Z(n_30500));
	notech_inv i_30534(.A(n_170584161), .Z(n_30502));
	notech_inv i_30535(.A(n_384964380), .Z(n_30504));
	notech_inv i_30536(.A(n_384864379), .Z(n_30505));
	notech_inv i_30538(.A(n_216384583), .Z(n_30506));
	notech_inv i_30539(.A(n_217484594), .Z(n_30507));
	notech_inv i_30540(.A(n_304167418), .Z(n_30508));
	notech_inv i_30541(.A(n_303667413), .Z(n_30509));
	notech_inv i_30543(.A(n_261285029), .Z(n_30510));
	notech_inv i_30544(.A(n_262385040), .Z(n_30511));
	notech_inv i_30545(.A(n_263485051), .Z(n_30512));
	notech_inv i_30547(.A(n_264585062), .Z(n_30513));
	notech_inv i_30548(.A(n_293885352), .Z(n_30514));
	notech_inv i_30549(.A(n_194866375), .Z(n_30515));
	notech_inv i_30550(.A(n_323260860), .Z(n_30516));
	notech_inv i_30551(.A(n_290067277), .Z(n_30517));
	notech_inv i_30552(.A(n_289867275), .Z(n_30518));
	notech_inv i_30553(.A(n_124545737), .Z(n_30519));
	notech_inv i_30554(.A(n_251347005), .Z(n_30520));
	notech_inv i_30555(.A(n_58532), .Z(n_30521));
	notech_inv i_30556(.A(n_303144465), .Z(n_30522));
	notech_inv i_30557(.A(n_303244466), .Z(n_30523));
	notech_inv i_30558(.A(n_19680), .Z(n_30524));
	notech_inv i_30559(.A(n_289167268), .Z(n_30525));
	notech_inv i_30560(.A(n_4450), .Z(n_30526));
	notech_inv i_30561(.A(n_288967266), .Z(n_30527));
	notech_inv i_30562(.A(n_336360991), .Z(n_30528));
	notech_inv i_30563(.A(n_119587122), .Z(n_30529));
	notech_inv i_30564(.A(n_121287139), .Z(n_30530));
	notech_inv i_30565(.A(n_122187148), .Z(n_30531));
	notech_inv i_30566(.A(n_123087157), .Z(n_30532));
	notech_inv i_30567(.A(n_123987166), .Z(n_30533));
	notech_inv i_30568(.A(n_124887175), .Z(n_30534));
	notech_inv i_30569(.A(n_125787184), .Z(n_30535));
	notech_inv i_30570(.A(n_126687193), .Z(n_30536));
	notech_inv i_30571(.A(n_127587202), .Z(n_30537));
	notech_inv i_30572(.A(n_4338), .Z(n_30538));
	notech_inv i_30573(.A(n_130987236), .Z(n_30539));
	notech_inv i_30574(.A(n_57688), .Z(n_30540));
	notech_inv i_30575(.A(n_131387240), .Z(n_30541));
	notech_inv i_30576(.A(n_140087327), .Z(n_30542));
	notech_inv i_30577(.A(n_140987336), .Z(n_30543));
	notech_inv i_30578(.A(n_141887345), .Z(n_30544));
	notech_inv i_30579(.A(n_142787354), .Z(n_30545));
	notech_inv i_30580(.A(n_143687363), .Z(n_30546));
	notech_inv i_30581(.A(n_30798), .Z(n_30547));
	notech_inv i_30583(.A(n_27378), .Z(n_30549));
	notech_inv i_30584(.A(n_30869), .Z(n_30550));
	notech_inv i_30585(.A(n_30785), .Z(n_30551));
	notech_inv i_30586(.A(n_29582), .Z(n_30552));
	notech_inv i_30587(.A(n_25121), .Z(n_30553));
	notech_inv i_30588(.A(n_29906), .Z(n_30554));
	notech_inv i_30589(.A(n_160487531), .Z(n_30555));
	notech_inv i_30590(.A(n_160987536), .Z(n_30556));
	notech_inv i_30591(.A(n_161287539), .Z(n_30557));
	notech_inv i_30592(.A(n_377364304), .Z(n_30558));
	notech_inv i_30593(.A(n_30468), .Z(n_30559));
	notech_inv i_30594(.A(n_32368), .Z(n_30560));
	notech_inv i_30595(.A(n_268667071), .Z(n_30561));
	notech_inv i_30596(.A(n_268467069), .Z(n_30562));
	notech_inv i_30597(.A(n_267767062), .Z(n_30563));
	notech_inv i_30598(.A(n_267567060), .Z(n_30564));
	notech_inv i_30599(.A(n_266667053), .Z(n_30565));
	notech_inv i_30600(.A(n_266067051), .Z(n_30566));
	notech_inv i_30601(.A(n_240488314), .Z(n_30567));
	notech_inv i_30602(.A(n_240788317), .Z(n_30568));
	notech_inv i_30603(.A(n_240988319), .Z(n_30569));
	notech_inv i_30604(.A(n_246488366), .Z(n_30570));
	notech_inv i_30605(.A(n_247288373), .Z(n_30571));
	notech_inv i_30606(.A(n_248688387), .Z(n_30572));
	notech_inv i_30607(.A(n_249388394), .Z(n_30573));
	notech_inv i_30608(.A(n_65029351), .Z(n_30574));
	notech_inv i_30609(.A(n_234966749), .Z(n_30575));
	notech_inv i_30610(.A(n_323560863), .Z(n_30576));
	notech_inv i_30612(.A(n_30395), .Z(n_30578));
	notech_inv i_30614(.A(n_234066740), .Z(n_30580));
	notech_inv i_30615(.A(n_264688547), .Z(n_30581));
	notech_inv i_30616(.A(n_265388554), .Z(n_30582));
	notech_inv i_30617(.A(n_233166731), .Z(n_30583));
	notech_inv i_30618(.A(n_266088561), .Z(n_30584));
	notech_inv i_30619(.A(n_266788568), .Z(n_30585));
	notech_inv i_30620(.A(n_2322), .Z(n_30586));
	notech_inv i_30621(.A(n_271388614), .Z(n_30587));
	notech_inv i_30622(.A(n_272088621), .Z(n_30588));
	notech_inv i_30623(.A(n_272788628), .Z(n_30589));
	notech_inv i_30624(.A(n_32219), .Z(n_30590));
	notech_inv i_30626(.A(n_26823), .Z(n_30592));
	notech_inv i_30627(.A(n_26822), .Z(n_30593));
	notech_inv i_30629(.A(n_56896), .Z(n_30595));
	notech_inv i_30633(.A(n_29417), .Z(n_30599));
	notech_inv i_30635(.A(n_442082451), .Z(n_30601));
	notech_inv i_30636(.A(n_284588745), .Z(n_30602));
	notech_inv i_30637(.A(n_288788787), .Z(n_30603));
	notech_inv i_30639(.A(n_26316138), .Z(n_30605));
	notech_inv i_30640(.A(n_26116136), .Z(n_30606));
	notech_inv i_30641(.A(n_222566626), .Z(n_30607));
	notech_inv i_30642(.A(n_221466615), .Z(n_30608));
	notech_inv i_30644(.A(n_22746), .Z(n_30610));
	notech_inv i_30645(.A(n_23351), .Z(n_30611));
	notech_inv i_30646(.A(n_23330), .Z(n_30612));
	notech_inv i_30647(.A(n_185866285), .Z(n_30613));
	notech_inv i_30648(.A(n_179566227), .Z(n_30614));
	notech_inv i_30649(.A(n_56035), .Z(n_30615));
	notech_inv i_30651(.A(n_78412540), .Z(n_30617));
	notech_inv i_30652(.A(n_32353), .Z(n_30618));
	notech_inv i_30653(.A(n_182666258), .Z(n_30619));
	notech_inv i_30654(.A(n_182466256), .Z(n_30620));
	notech_inv i_30655(.A(n_172766169), .Z(n_30621));
	notech_inv i_30656(.A(n_343489317), .Z(n_30622));
	notech_inv i_30657(.A(n_181966251), .Z(n_30623));
	notech_inv i_30658(.A(n_2025), .Z(n_30624));
	notech_inv i_30659(.A(n_344289324), .Z(n_30625));
	notech_inv i_30660(.A(n_344589327), .Z(n_30626));
	notech_inv i_30661(.A(n_3469), .Z(n_30627));
	notech_inv i_30662(.A(n_26086), .Z(n_30628));
	notech_inv i_30663(.A(n_58682), .Z(n_30629));
	notech_inv i_30664(.A(n_305344487), .Z(n_30630));
	notech_inv i_30665(.A(n_303044464), .Z(n_30631));
	notech_inv i_30666(.A(n_175266188), .Z(n_30632));
	notech_inv i_30667(.A(n_28552), .Z(n_30633));
	notech_inv i_30668(.A(n_326860896), .Z(n_30634));
	notech_inv i_30669(.A(n_365964190), .Z(n_30635));
	notech_inv i_30670(.A(n_19645), .Z(n_30636));
	notech_inv i_30671(.A(n_389664427), .Z(n_30637));
	notech_inv i_30672(.A(\add_len_pc[13] ), .Z(n_30638));
	notech_inv i_30673(.A(\add_len_pc[10] ), .Z(n_30639));
	notech_inv i_30674(.A(n_383364364), .Z(n_30640));
	notech_inv i_30675(.A(n_387164402), .Z(n_30641));
	notech_inv i_30676(.A(n_285763759), .Z(n_30642));
	notech_inv i_30677(.A(n_384664377), .Z(n_30643));
	notech_inv i_30678(.A(n_384564376), .Z(n_30644));
	notech_inv i_30679(.A(n_384464375), .Z(n_30645));
	notech_inv i_30680(.A(n_256563512), .Z(n_30646));
	notech_inv i_30681(.A(n_256763514), .Z(n_30647));
	notech_inv i_30682(.A(n_1849), .Z(n_30648));
	notech_inv i_30683(.A(n_83245324), .Z(n_30649));
	notech_inv i_30684(.A(n_2091), .Z(n_30650));
	notech_inv i_30685(.A(n_2178), .Z(n_30651));
	notech_inv i_30686(.A(n_210833639), .Z(n_30652));
	notech_inv i_30687(.A(n_1816), .Z(n_30653));
	notech_inv i_30688(.A(n_353728636), .Z(n_30654));
	notech_inv i_30690(.A(n_380664337), .Z(n_30656));
	notech_inv i_30691(.A(n_380364334), .Z(n_30657));
	notech_inv i_30692(.A(n_232463321), .Z(n_30658));
	notech_inv i_30693(.A(n_377864309), .Z(n_30659));
	notech_inv i_30694(.A(n_179862826), .Z(n_30660));
	notech_inv i_30695(.A(n_61819), .Z(\opcode[3] ));
	notech_inv i_30696(.A(n_162262654), .Z(n_30662));
	notech_inv i_30698(.A(n_32241), .Z(n_30664));
	notech_inv i_30699(.A(n_305544489), .Z(n_30665));
	notech_inv i_30700(.A(n_375464285), .Z(n_30666));
	notech_inv i_30701(.A(n_128990656), .Z(n_30667));
	notech_inv i_30702(.A(n_351785925), .Z(n_30668));
	notech_inv i_30703(.A(n_125390620), .Z(n_30669));
	notech_inv i_30704(.A(n_57041), .Z(n_30670));
	notech_inv i_30705(.A(n_56583), .Z(n_30671));
	notech_inv i_30706(.A(n_57717), .Z(n_30672));
	notech_inv i_30708(.A(n_3298), .Z(n_30674));
	notech_inv i_30709(.A(n_152690893), .Z(n_30675));
	notech_inv i_30710(.A(n_179291159), .Z(n_30676));
	notech_inv i_30711(.A(n_352864060), .Z(n_30677));
	notech_inv i_30712(.A(n_32323), .Z(n_30678));
	notech_inv i_30713(.A(n_32215), .Z(n_30679));
	notech_inv i_30714(.A(n_347271361), .Z(n_30680));
	notech_inv i_30715(.A(n_349671381), .Z(n_30681));
	notech_inv i_30716(.A(n_212433655), .Z(n_30682));
	notech_inv i_30717(.A(n_211833649), .Z(n_30683));
	notech_inv i_30718(.A(n_223191585), .Z(n_30684));
	notech_inv i_30719(.A(n_223491588), .Z(n_30685));
	notech_inv i_30720(.A(n_223691590), .Z(n_30686));
	notech_inv i_30721(.A(n_27842), .Z(n_30687));
	notech_inv i_30722(.A(n_27826), .Z(n_30688));
	notech_inv i_30723(.A(n_27823), .Z(n_30691));
	notech_inv i_30724(.A(n_231291666), .Z(n_30692));
	notech_inv i_30725(.A(n_27923), .Z(n_30696));
	notech_inv i_30726(.A(n_32321), .Z(n_30698));
	notech_inv i_30727(.A(n_231891672), .Z(n_30699));
	notech_inv i_30728(.A(n_57206), .Z(n_30700));
	notech_inv i_30729(.A(n_23845), .Z(n_30701));
	notech_inv i_30730(.A(n_3274), .Z(n_30702));
	notech_inv i_30731(.A(n_3260), .Z(n_30703));
	notech_inv i_30732(.A(n_3248), .Z(n_30704));
	notech_inv i_30733(.A(n_3241), .Z(n_30705));
	notech_inv i_30734(.A(n_3214), .Z(n_30706));
	notech_inv i_30735(.A(n_3127), .Z(n_30707));
	notech_inv i_30736(.A(n_3108), .Z(n_30708));
	notech_inv i_30740(.A(n_61119), .Z(n_30712));
	notech_inv i_30742(.A(n_19629), .Z(n_30714));
	notech_inv i_30743(.A(n_57724), .Z(n_30715));
	notech_inv i_30744(.A(n_295663854), .Z(n_30716));
	notech_inv i_30745(.A(n_294963847), .Z(n_30717));
	notech_inv i_30746(.A(n_294263840), .Z(n_30718));
	notech_inv i_30747(.A(n_59599), .Z(n_30720));
	notech_inv i_30748(.A(n_3456), .Z(n_30722));
	notech_inv i_30749(.A(n_115290519), .Z(n_30724));
	notech_inv i_30750(.A(n_54327), .Z(n_30726));
	notech_inv i_30751(.A(n_61775), .Z(\opcode[0] ));
	notech_inv i_30752(.A(n_315792476), .Z(n_30730));
	notech_inv i_30753(.A(n_290763807), .Z(n_30731));
	notech_inv i_30754(.A(n_286163763), .Z(n_30732));
	notech_inv i_30755(.A(n_286063762), .Z(n_30733));
	notech_inv i_30756(.A(n_281863720), .Z(n_30734));
	notech_inv i_30757(.A(n_281763719), .Z(n_30735));
	notech_inv i_30758(.A(n_2111), .Z(n_30736));
	notech_inv i_30759(.A(n_340061028), .Z(n_30737));
	notech_inv i_30760(.A(n_340161029), .Z(n_30738));
	notech_inv i_30761(.A(n_339761025), .Z(n_30739));
	notech_inv i_30762(.A(n_278663690), .Z(n_30740));
	notech_inv i_30763(.A(n_156694049), .Z(n_30741));
	notech_inv i_30764(.A(n_163194114), .Z(n_30742));
	notech_inv i_30765(.A(n_29229), .Z(n_30743));
	notech_inv i_30766(.A(n_340261030), .Z(n_30744));
	notech_inv i_30767(.A(n_2765), .Z(n_30745));
	notech_inv i_30768(.A(n_2756), .Z(n_30746));
	notech_inv i_30769(.A(n_256363510), .Z(n_30747));
	notech_inv i_30770(.A(n_54405), .Z(n_30748));
	notech_inv i_30771(.A(n_280595278), .Z(n_30749));
	notech_inv i_30772(.A(n_248763435), .Z(n_30750));
	notech_inv i_30773(.A(n_30865), .Z(n_30751));
	notech_inv i_30775(.A(n_20902), .Z(n_30753));
	notech_inv i_30776(.A(n_222663225), .Z(n_30754));
	notech_inv i_30777(.A(n_222463223), .Z(n_30755));
	notech_inv i_30778(.A(n_197963006), .Z(n_30756));
	notech_inv i_30779(.A(n_197863005), .Z(n_30757));
	notech_inv i_30780(.A(n_326695682), .Z(n_30758));
	notech_inv i_30781(.A(fecx), .Z(n_30759));
	notech_inv i_30782(.A(sav_ecx[0]), .Z(n_30760));
	notech_inv i_30783(.A(sav_ecx[1]), .Z(n_30761));
	notech_inv i_30784(.A(sav_ecx[3]), .Z(n_30762));
	notech_inv i_30785(.A(sav_ecx[4]), .Z(n_30763));
	notech_inv i_30786(.A(sav_ecx[7]), .Z(n_30764));
	notech_inv i_30787(.A(sav_ecx[8]), .Z(n_30765));
	notech_inv i_30788(.A(sav_ecx[9]), .Z(n_30766));
	notech_inv i_30789(.A(sav_ecx[10]), .Z(n_30767));
	notech_inv i_30790(.A(sav_ecx[11]), .Z(n_30768));
	notech_inv i_30791(.A(sav_ecx[12]), .Z(n_30769));
	notech_inv i_30792(.A(sav_ecx[13]), .Z(n_30770));
	notech_inv i_30793(.A(sav_ecx[14]), .Z(n_30771));
	notech_inv i_30794(.A(sav_ecx[15]), .Z(n_30772));
	notech_inv i_30795(.A(sav_ecx[21]), .Z(n_30773));
	notech_inv i_30796(.A(sav_ecx[22]), .Z(n_30774));
	notech_inv i_30797(.A(fesp), .Z(n_30775));
	notech_inv i_30798(.A(sav_esp[0]), .Z(n_30776));
	notech_inv i_30799(.A(sav_esp[1]), .Z(n_30777));
	notech_inv i_30800(.A(sav_esp[2]), .Z(n_30778));
	notech_inv i_30801(.A(sav_esp[3]), .Z(n_30779));
	notech_inv i_30802(.A(sav_esp[4]), .Z(n_30781));
	notech_inv i_30803(.A(sav_esp[5]), .Z(n_30782));
	notech_inv i_30804(.A(sav_esp[6]), .Z(n_30783));
	notech_inv i_30805(.A(sav_esp[8]), .Z(n_30784));
	notech_inv i_30806(.A(sav_esp[9]), .Z(n_30787));
	notech_inv i_30807(.A(sav_esp[10]), .Z(n_30789));
	notech_inv i_30808(.A(sav_esp[11]), .Z(n_30790));
	notech_inv i_30809(.A(sav_esp[12]), .Z(n_30791));
	notech_inv i_30810(.A(sav_esp[14]), .Z(n_30793));
	notech_inv i_30811(.A(sav_esp[15]), .Z(n_30794));
	notech_inv i_30812(.A(sav_esp[16]), .Z(n_30795));
	notech_inv i_30813(.A(sav_esp[17]), .Z(n_30797));
	notech_inv i_30814(.A(sav_esp[18]), .Z(n_30799));
	notech_inv i_30815(.A(sav_esp[19]), .Z(n_30801));
	notech_inv i_30816(.A(sav_esp[26]), .Z(n_30802));
	notech_inv i_30817(.A(sav_esp[27]), .Z(n_30805));
	notech_inv i_30818(.A(sav_esp[28]), .Z(n_30806));
	notech_inv i_30819(.A(sav_esp[29]), .Z(n_30807));
	notech_inv i_30820(.A(sav_esp[30]), .Z(n_30808));
	notech_inv i_30821(.A(sav_esp[31]), .Z(n_30809));
	notech_inv i_30822(.A(sav_esi[0]), .Z(n_30810));
	notech_inv i_30823(.A(sav_esi[1]), .Z(n_30811));
	notech_inv i_30824(.A(sav_esi[3]), .Z(n_30812));
	notech_inv i_30825(.A(sav_esi[8]), .Z(n_30813));
	notech_inv i_30826(.A(sav_esi[9]), .Z(n_30814));
	notech_inv i_30827(.A(sav_esi[10]), .Z(n_30816));
	notech_inv i_30828(.A(sav_esi[11]), .Z(n_30818));
	notech_inv i_30829(.A(sav_esi[12]), .Z(n_30819));
	notech_inv i_30830(.A(sav_esi[13]), .Z(n_30820));
	notech_inv i_30831(.A(sav_esi[15]), .Z(n_30821));
	notech_inv i_30832(.A(sav_esi[20]), .Z(n_30824));
	notech_inv i_30833(.A(sav_esi[21]), .Z(n_30825));
	notech_inv i_30834(.A(sav_esi[22]), .Z(n_30826));
	notech_inv i_30835(.A(sav_esi[23]), .Z(n_30827));
	notech_inv i_30836(.A(sav_esi[24]), .Z(n_30830));
	notech_inv i_30837(.A(sav_esi[25]), .Z(n_30831));
	notech_inv i_30838(.A(sav_edi[0]), .Z(n_30832));
	notech_inv i_30839(.A(sav_edi[1]), .Z(n_30833));
	notech_inv i_30840(.A(sav_edi[2]), .Z(n_30834));
	notech_inv i_30841(.A(sav_edi[3]), .Z(n_30836));
	notech_inv i_30843(.A(sav_edi[4]), .Z(n_30837));
	notech_inv i_30844(.A(sav_edi[5]), .Z(n_30838));
	notech_inv i_30845(.A(sav_edi[6]), .Z(n_30840));
	notech_inv i_30846(.A(sav_edi[7]), .Z(n_30841));
	notech_inv i_30847(.A(sav_edi[8]), .Z(n_30843));
	notech_inv i_30848(.A(sav_edi[9]), .Z(n_30844));
	notech_inv i_30850(.A(sav_edi[10]), .Z(n_30845));
	notech_inv i_30851(.A(sav_edi[11]), .Z(n_30846));
	notech_inv i_30852(.A(sav_edi[12]), .Z(n_30847));
	notech_inv i_30853(.A(sav_edi[13]), .Z(n_30848));
	notech_inv i_30854(.A(sav_edi[15]), .Z(n_30850));
	notech_inv i_30855(.A(sav_edi[20]), .Z(n_30851));
	notech_inv i_30856(.A(sav_edi[21]), .Z(n_30852));
	notech_inv i_30857(.A(sav_edi[22]), .Z(n_30853));
	notech_inv i_30858(.A(sav_edi[23]), .Z(n_30854));
	notech_inv i_30859(.A(sav_edi[24]), .Z(n_30856));
	notech_inv i_30860(.A(sav_edi[25]), .Z(n_30857));
	notech_inv i_30861(.A(sav_edi[30]), .Z(n_30859));
	notech_inv i_30862(.A(sav_epc[0]), .Z(n_30860));
	notech_inv i_30863(.A(sav_epc[1]), .Z(n_30861));
	notech_inv i_30864(.A(sav_epc[2]), .Z(n_30862));
	notech_inv i_30865(.A(sav_epc[3]), .Z(n_30863));
	notech_inv i_30866(.A(sav_epc[4]), .Z(n_30866));
	notech_inv i_30871(.A(sav_epc[5]), .Z(n_30870));
	notech_inv i_30872(.A(sav_epc[6]), .Z(n_30871));
	notech_inv i_30873(.A(sav_epc[7]), .Z(n_30872));
	notech_inv i_30874(.A(sav_epc[8]), .Z(n_30873));
	notech_inv i_30875(.A(sav_epc[9]), .Z(n_30874));
	notech_inv i_30876(.A(sav_epc[10]), .Z(n_30875));
	notech_inv i_30877(.A(sav_epc[11]), .Z(n_30876));
	notech_inv i_30878(.A(sav_epc[12]), .Z(n_30877));
	notech_inv i_30879(.A(sav_epc[13]), .Z(n_30878));
	notech_inv i_30880(.A(sav_epc[14]), .Z(n_30879));
	notech_inv i_30881(.A(sav_epc[15]), .Z(n_30880));
	notech_inv i_30882(.A(n_158062612), .Z(n_30881));
	notech_inv i_30883(.A(sav_epc[16]), .Z(n_30882));
	notech_inv i_30884(.A(sav_epc[17]), .Z(n_30883));
	notech_inv i_30885(.A(sav_epc[18]), .Z(n_30884));
	notech_inv i_30886(.A(sav_epc[19]), .Z(n_30885));
	notech_inv i_30887(.A(n_157162603), .Z(n_30886));
	notech_inv i_30888(.A(sav_epc[26]), .Z(n_30887));
	notech_inv i_30889(.A(sav_epc[27]), .Z(n_30888));
	notech_inv i_30890(.A(sav_epc[28]), .Z(n_30889));
	notech_inv i_30891(.A(n_155562587), .Z(n_30890));
	notech_inv i_30892(.A(sav_epc[29]), .Z(n_30892));
	notech_inv i_30893(.A(sav_epc[31]), .Z(n_30893));
	notech_inv i_30894(.A(\nbus_11287[0] ), .Z(n_30894));
	notech_inv i_30895(.A(n_156062592), .Z(n_30895));
	notech_inv i_30896(.A(n_8327), .Z(n_30897));
	notech_inv i_30897(.A(n_32394), .Z(n_30898));
	notech_inv i_30898(.A(n_309860726), .Z(n_30899));
	notech_inv i_30899(.A(n_61806), .Z(n_30900));
	notech_inv i_30900(.A(n_312460752), .Z(n_30901));
	notech_inv i_30901(.A(n_61958), .Z(\opcode[1] ));
	notech_inv i_30902(.A(n_275660605), .Z(n_30903));
	notech_inv i_30903(.A(n_336260990), .Z(n_30904));
	notech_inv i_30904(.A(n_338261010), .Z(n_30905));
	notech_inv i_30905(.A(n_330960937), .Z(n_30906));
	notech_inv i_30906(.A(n_333960967), .Z(n_30907));
	notech_inv i_30907(.A(n_333860966), .Z(n_30908));
	notech_inv i_30908(.A(n_333760965), .Z(n_30909));
	notech_inv i_30909(.A(n_165695997), .Z(n_30910));
	notech_inv i_30910(.A(n_163196017), .Z(n_30911));
	notech_inv i_30911(.A(n_329060918), .Z(n_30912));
	notech_inv i_30912(.A(n_19364), .Z(n_30913));
	notech_inv i_30913(.A(n_1634), .Z(n_30915));
	notech_inv i_30914(.A(n_327460902), .Z(n_30917));
	notech_inv i_30915(.A(n_1457), .Z(n_30918));
	notech_inv i_30916(.A(n_143460302), .Z(n_30921));
	notech_inv i_30917(.A(n_143360301), .Z(n_30922));
	notech_inv i_30918(.A(n_1464), .Z(n_30923));
	notech_inv i_30919(.A(n_18524), .Z(n_30924));
	notech_inv i_30920(.A(n_16223), .Z(n_30925));
	notech_inv i_30921(.A(n_317260800), .Z(n_30926));
	notech_inv i_30922(.A(n_16397), .Z(n_30927));
	notech_inv i_30923(.A(n_15874), .Z(n_30928));
	notech_inv i_30924(.A(n_15880), .Z(n_30929));
	notech_inv i_30925(.A(n_15898), .Z(n_30930));
	notech_inv i_30926(.A(n_15904), .Z(n_30931));
	notech_inv i_30927(.A(n_15910), .Z(n_30932));
	notech_inv i_30928(.A(n_15916), .Z(n_30933));
	notech_inv i_30929(.A(n_15958), .Z(n_30934));
	notech_inv i_30930(.A(pipe_mul[0]), .Z(n_30935));
	notech_inv i_30931(.A(eval_flag), .Z(n_30936));
	notech_inv i_30932(.A(rep_en1), .Z(n_30937));
	notech_inv i_30933(.A(rep_en4), .Z(n_30938));
	notech_inv i_30934(.A(nCF), .Z(n_30939));
	notech_inv i_30935(.A(n_7415), .Z(n_30940));
	notech_inv i_30936(.A(n_8508), .Z(n_30941));
	notech_inv i_30937(.A(nAF), .Z(n_30942));
	notech_inv i_30938(.A(nSF), .Z(n_30943));
	notech_inv i_30939(.A(n_364350916), .Z(n_30944));
	notech_inv i_30940(.A(n_14232), .Z(n_30945));
	notech_inv i_30941(.A(n_14229), .Z(n_30946));
	notech_inv i_30942(.A(n_20384), .Z(n_30947));
	notech_inv i_30943(.A(n_20420), .Z(n_30948));
	notech_inv i_30944(.A(\nbus_11352[9] ), .Z(n_30949));
	notech_inv i_30945(.A(\nbus_11352[10] ), .Z(n_30950));
	notech_inv i_30946(.A(n_15522), .Z(n_30951));
	notech_inv i_30947(.A(n_15528), .Z(n_30952));
	notech_inv i_30948(.A(n_15534), .Z(n_30953));
	notech_inv i_30949(.A(n_15540), .Z(n_30954));
	notech_inv i_30950(.A(n_15546), .Z(n_30955));
	notech_inv i_30951(.A(n_15552), .Z(n_30956));
	notech_inv i_30952(.A(n_15558), .Z(n_30957));
	notech_inv i_30953(.A(n_15564), .Z(n_30958));
	notech_inv i_30954(.A(n_15606), .Z(n_30959));
	notech_inv i_30955(.A(n_304560674), .Z(n_30960));
	notech_inv i_30956(.A(\nbus_11326[0] ), .Z(n_30961));
	notech_inv i_30957(.A(n_303260661), .Z(n_30962));
	notech_inv i_30958(.A(n_302460653), .Z(n_30963));
	notech_inv i_30959(.A(n_302560654), .Z(n_30964));
	notech_inv i_30960(.A(n_2844), .Z(n_30965));
	notech_inv i_30961(.A(n_14337), .Z(n_30966));
	notech_inv i_30962(.A(temp_sp[0]), .Z(n_30967));
	notech_inv i_30963(.A(n_14342), .Z(n_30968));
	notech_inv i_30964(.A(temp_sp[1]), .Z(n_30969));
	notech_inv i_30965(.A(n_14347), .Z(n_30970));
	notech_inv i_30966(.A(temp_sp[2]), .Z(n_30971));
	notech_inv i_30967(.A(n_14352), .Z(n_30972));
	notech_inv i_30968(.A(temp_sp[3]), .Z(n_30973));
	notech_inv i_30969(.A(n_14357), .Z(n_30974));
	notech_inv i_30970(.A(temp_sp[4]), .Z(n_30975));
	notech_inv i_30971(.A(n_14362), .Z(n_30976));
	notech_inv i_30972(.A(temp_sp[5]), .Z(n_30977));
	notech_inv i_30973(.A(n_14367), .Z(n_30978));
	notech_inv i_30974(.A(temp_sp[6]), .Z(n_30979));
	notech_inv i_30975(.A(n_14372), .Z(n_30980));
	notech_inv i_30976(.A(temp_sp[7]), .Z(n_30981));
	notech_inv i_30977(.A(n_14377), .Z(n_30982));
	notech_inv i_30978(.A(temp_sp[8]), .Z(n_30983));
	notech_inv i_30979(.A(n_14382), .Z(n_30984));
	notech_inv i_30980(.A(temp_sp[9]), .Z(n_30985));
	notech_inv i_30981(.A(n_14387), .Z(n_30986));
	notech_inv i_30982(.A(temp_sp[10]), .Z(n_30987));
	notech_inv i_30983(.A(n_14392), .Z(n_30988));
	notech_inv i_30984(.A(temp_sp[11]), .Z(n_30989));
	notech_inv i_30985(.A(n_14397), .Z(n_30990));
	notech_inv i_30986(.A(temp_sp[12]), .Z(n_30991));
	notech_inv i_30987(.A(n_14402), .Z(n_30992));
	notech_inv i_30988(.A(temp_sp[13]), .Z(n_30993));
	notech_inv i_30989(.A(n_14407), .Z(n_30994));
	notech_inv i_30990(.A(temp_sp[14]), .Z(n_30995));
	notech_inv i_30991(.A(n_14412), .Z(n_30996));
	notech_inv i_30992(.A(temp_sp[15]), .Z(n_30997));
	notech_inv i_30993(.A(n_14417), .Z(n_30998));
	notech_inv i_30994(.A(temp_sp[16]), .Z(n_30999));
	notech_inv i_30995(.A(n_2823), .Z(n_31000));
	notech_inv i_30996(.A(n_14422), .Z(n_31001));
	notech_inv i_30997(.A(temp_sp[17]), .Z(n_31002));
	notech_inv i_30998(.A(n_14427), .Z(n_31003));
	notech_inv i_30999(.A(temp_sp[18]), .Z(n_31004));
	notech_inv i_31000(.A(n_14432), .Z(n_31005));
	notech_inv i_31001(.A(temp_sp[19]), .Z(n_31006));
	notech_inv i_31002(.A(n_14437), .Z(n_31007));
	notech_inv i_31003(.A(temp_sp[20]), .Z(n_31008));
	notech_inv i_31004(.A(n_14442), .Z(n_31009));
	notech_inv i_31005(.A(temp_sp[21]), .Z(n_31010));
	notech_inv i_31006(.A(n_14447), .Z(n_31011));
	notech_inv i_31007(.A(temp_sp[22]), .Z(n_31012));
	notech_inv i_31008(.A(n_14452), .Z(n_31013));
	notech_inv i_31009(.A(temp_sp[23]), .Z(n_31014));
	notech_inv i_31010(.A(n_14457), .Z(n_31015));
	notech_inv i_31011(.A(temp_sp[24]), .Z(n_31016));
	notech_inv i_31012(.A(n_14462), .Z(n_31017));
	notech_inv i_31013(.A(temp_sp[25]), .Z(n_31018));
	notech_inv i_31014(.A(n_14467), .Z(n_31019));
	notech_inv i_31015(.A(temp_sp[26]), .Z(n_31020));
	notech_inv i_31016(.A(n_14472), .Z(n_31021));
	notech_inv i_31017(.A(temp_sp[27]), .Z(n_31022));
	notech_inv i_31018(.A(n_14477), .Z(n_31023));
	notech_inv i_31019(.A(temp_sp[28]), .Z(n_31024));
	notech_inv i_31020(.A(n_14482), .Z(n_31025));
	notech_inv i_31021(.A(temp_sp[29]), .Z(n_31026));
	notech_inv i_31022(.A(n_14487), .Z(n_31027));
	notech_inv i_31023(.A(temp_sp[30]), .Z(n_31028));
	notech_inv i_31024(.A(n_14492), .Z(n_31029));
	notech_inv i_31025(.A(temp_sp[31]), .Z(n_31030));
	notech_inv i_31026(.A(n_15170), .Z(n_31031));
	notech_inv i_31027(.A(n_15194), .Z(n_31032));
	notech_inv i_31028(.A(n_15200), .Z(n_31033));
	notech_inv i_31029(.A(n_15206), .Z(n_31034));
	notech_inv i_31032(.A(n_15212), .Z(n_31035));
	notech_inv i_31034(.A(n_275560604), .Z(n_31036));
	notech_inv i_31035(.A(n_12644), .Z(n_31037));
	notech_inv i_31036(.A(n_12650), .Z(n_31038));
	notech_inv i_31037(.A(n_12692), .Z(n_31039));
	notech_inv i_31038(.A(n_12728), .Z(n_31040));
	notech_inv i_31039(.A(n_12746), .Z(n_31041));
	notech_inv i_31040(.A(n_12752), .Z(n_31042));
	notech_inv i_31041(.A(n_12758), .Z(n_31043));
	notech_inv i_31042(.A(n_12776), .Z(n_31044));
	notech_inv i_31043(.A(n_12800), .Z(n_31045));
	notech_inv i_31044(.A(n_12812), .Z(n_31046));
	notech_inv i_31045(.A(n_12818), .Z(n_31049));
	notech_inv i_31046(.A(n_12824), .Z(n_31050));
	notech_inv i_31047(.A(\nbus_14542[1] ), .Z(n_31051));
	notech_inv i_31049(.A(\nbus_14542[3] ), .Z(n_31052));
	notech_inv i_31050(.A(\nbus_14542[4] ), .Z(n_31053));
	notech_inv i_31051(.A(\nbus_14542[6] ), .Z(n_31054));
	notech_inv i_31052(.A(\nbus_14542[7] ), .Z(n_31055));
	notech_inv i_31053(.A(\nbus_14542[8] ), .Z(n_31056));
	notech_inv i_31054(.A(\nbus_14542[9] ), .Z(n_31057));
	notech_inv i_31055(.A(\nbus_14542[10] ), .Z(n_31058));
	notech_inv i_31056(.A(\nbus_14542[11] ), .Z(n_31059));
	notech_inv i_31057(.A(\nbus_14542[12] ), .Z(n_31060));
	notech_inv i_31058(.A(\nbus_14542[13] ), .Z(n_31061));
	notech_inv i_31059(.A(\nbus_14542[14] ), .Z(n_31062));
	notech_inv i_31060(.A(\nbus_14542[15] ), .Z(n_31063));
	notech_inv i_31061(.A(n_11275), .Z(n_31064));
	notech_inv i_31063(.A(n_11281), .Z(n_31065));
	notech_inv i_31064(.A(mask8b[1]), .Z(n_31066));
	notech_inv i_31065(.A(mask8b[2]), .Z(n_31069));
	notech_inv i_31066(.A(\nbus_11301[0] ), .Z(n_31070));
	notech_inv i_31067(.A(n_13617), .Z(n_31073));
	notech_inv i_31068(.A(n_13623), .Z(n_31076));
	notech_inv i_31069(.A(n_13629), .Z(n_31077));
	notech_inv i_31070(.A(n_13665), .Z(n_31078));
	notech_inv i_31071(.A(n_13671), .Z(n_31079));
	notech_inv i_31072(.A(n_13701), .Z(n_31080));
	notech_inv i_31073(.A(n_13719), .Z(n_31081));
	notech_inv i_31074(.A(n_13725), .Z(n_31082));
	notech_inv i_31075(.A(n_12310), .Z(n_31083));
	notech_inv i_31076(.A(n_12316), .Z(n_31084));
	notech_inv i_31077(.A(n_12328), .Z(n_31085));
	notech_inv i_31078(.A(n_12376), .Z(n_31086));
	notech_inv i_31079(.A(n_12394), .Z(n_31087));
	notech_inv i_31080(.A(n_12406), .Z(n_31088));
	notech_inv i_31081(.A(n_12448), .Z(n_31089));
	notech_inv i_31082(.A(n_12460), .Z(n_31090));
	notech_inv i_31083(.A(n_12478), .Z(n_31091));
	notech_inv i_31084(.A(n_11941), .Z(n_31092));
	notech_inv i_31085(.A(n_11953), .Z(n_31093));
	notech_inv i_31086(.A(n_11971), .Z(n_31094));
	notech_inv i_31087(.A(n_12019), .Z(n_31095));
	notech_inv i_31088(.A(n_12037), .Z(n_31096));
	notech_inv i_31089(.A(n_12049), .Z(n_31097));
	notech_inv i_31090(.A(n_12103), .Z(n_31100));
	notech_inv i_31091(.A(n_12121), .Z(n_31101));
	notech_inv i_31092(.A(n_7949), .Z(n_31102));
	notech_inv i_31093(.A(n_7954), .Z(n_31103));
	notech_inv i_31094(.A(n_7959), .Z(n_31104));
	notech_inv i_31095(.A(n_7964), .Z(n_31105));
	notech_inv i_31096(.A(n_7969), .Z(n_31106));
	notech_inv i_31097(.A(n_7974), .Z(n_31107));
	notech_inv i_31098(.A(n_7979), .Z(n_31108));
	notech_inv i_31099(.A(n_7984), .Z(n_31109));
	notech_inv i_31100(.A(n_7989), .Z(n_31110));
	notech_inv i_31101(.A(n_7994), .Z(n_31111));
	notech_inv i_31102(.A(n_7999), .Z(n_31112));
	notech_inv i_31103(.A(n_8004), .Z(n_31113));
	notech_inv i_31104(.A(n_8009), .Z(n_31114));
	notech_inv i_31105(.A(n_8014), .Z(n_31115));
	notech_inv i_31106(.A(n_8019), .Z(n_31116));
	notech_inv i_31107(.A(n_8024), .Z(n_31117));
	notech_inv i_31108(.A(n_8029), .Z(n_31120));
	notech_inv i_31109(.A(n_8034), .Z(n_31121));
	notech_inv i_31110(.A(n_8039), .Z(n_31124));
	notech_inv i_31111(.A(n_8044), .Z(n_31127));
	notech_inv i_31112(.A(n_8049), .Z(n_31128));
	notech_inv i_31113(.A(n_8054), .Z(n_31129));
	notech_inv i_31114(.A(n_8059), .Z(n_31130));
	notech_inv i_31115(.A(n_8064), .Z(n_31131));
	notech_inv i_31116(.A(n_8069), .Z(n_31132));
	notech_inv i_31117(.A(n_8074), .Z(n_31133));
	notech_inv i_31118(.A(n_8079), .Z(n_31134));
	notech_inv i_31119(.A(n_8084), .Z(n_31135));
	notech_inv i_31120(.A(n_8089), .Z(n_31136));
	notech_inv i_31121(.A(n_8094), .Z(n_31137));
	notech_inv i_31124(.A(n_9821), .Z(n_31140));
	notech_inv i_31125(.A(n_9831), .Z(n_31141));
	notech_inv i_31126(.A(\nbus_11289[5] ), .Z(n_31142));
	notech_inv i_31127(.A(n_9896), .Z(n_31143));
	notech_inv i_31128(.A(n_9901), .Z(n_31144));
	notech_inv i_31129(.A(n_9906), .Z(n_31145));
	notech_inv i_31130(.A(n_9911), .Z(n_31146));
	notech_inv i_31131(.A(n_9916), .Z(n_31147));
	notech_inv i_31132(.A(n_9921), .Z(n_31148));
	notech_inv i_31133(.A(n_9926), .Z(n_31149));
	notech_inv i_31134(.A(n_9931), .Z(n_31150));
	notech_inv i_31135(.A(n_9936), .Z(n_31151));
	notech_inv i_31136(.A(n_9941), .Z(n_31152));
	notech_inv i_31137(.A(n_9946), .Z(n_31153));
	notech_inv i_31138(.A(n_9951), .Z(n_31154));
	notech_inv i_31139(.A(n_9956), .Z(n_31155));
	notech_inv i_31140(.A(n_9961), .Z(n_31156));
	notech_inv i_31141(.A(n_9966), .Z(n_31157));
	notech_inv i_31142(.A(n_9971), .Z(n_31158));
	notech_inv i_31143(.A(\nbus_11289[16] ), .Z(n_31159));
	notech_inv i_31144(.A(nZF), .Z(n_31160));
	notech_inv i_31145(.A(n_11662), .Z(n_31161));
	notech_inv i_31148(.A(n_11674), .Z(n_31162));
	notech_inv i_31149(.A(n_11680), .Z(n_31163));
	notech_inv i_31150(.A(n_11686), .Z(n_31164));
	notech_inv i_31151(.A(n_11698), .Z(n_31165));
	notech_inv i_31152(.A(n_11710), .Z(n_31166));
	notech_inv i_31153(.A(n_11722), .Z(n_31167));
	notech_inv i_31154(.A(n_11728), .Z(n_31168));
	notech_inv i_31155(.A(n_11734), .Z(n_31169));
	notech_inv i_31156(.A(n_11746), .Z(n_31170));
	notech_inv i_31157(.A(n_11752), .Z(n_31171));
	notech_inv i_31158(.A(nbus_14541[0]), .Z(n_31172));
	notech_inv i_31159(.A(nbus_14541[1]), .Z(n_31173));
	notech_inv i_31161(.A(nbus_14541[2]), .Z(n_31174));
	notech_inv i_31162(.A(nbus_14541[3]), .Z(n_31175));
	notech_inv i_31163(.A(nbus_14541[4]), .Z(n_31176));
	notech_inv i_31164(.A(nbus_14541[5]), .Z(n_31177));
	notech_inv i_31165(.A(nbus_14541[6]), .Z(n_31178));
	notech_inv i_31166(.A(nbus_14541[8]), .Z(n_31179));
	notech_inv i_31167(.A(nbus_14541[9]), .Z(n_31180));
	notech_inv i_31168(.A(nbus_14541[10]), .Z(n_31181));
	notech_inv i_31169(.A(nbus_14541[11]), .Z(n_31182));
	notech_inv i_31170(.A(nbus_14541[12]), .Z(n_31183));
	notech_inv i_31171(.A(nbus_14541[16]), .Z(n_31184));
	notech_inv i_31172(.A(nbus_14541[17]), .Z(n_31185));
	notech_inv i_31173(.A(nbus_14541[18]), .Z(n_31186));
	notech_inv i_31174(.A(nbus_14541[19]), .Z(n_31187));
	notech_inv i_31175(.A(nbus_14541[20]), .Z(n_31188));
	notech_inv i_31177(.A(nbus_14541[21]), .Z(n_31189));
	notech_inv i_31178(.A(nbus_14541[22]), .Z(n_31190));
	notech_inv i_31179(.A(nbus_14541[23]), .Z(n_31191));
	notech_inv i_31180(.A(nbus_14541[24]), .Z(n_31192));
	notech_inv i_31181(.A(nbus_14541[25]), .Z(n_31193));
	notech_inv i_31182(.A(nbus_14541[26]), .Z(n_31194));
	notech_inv i_31183(.A(nbus_14541[27]), .Z(n_31195));
	notech_inv i_31184(.A(nbus_14541[28]), .Z(n_31196));
	notech_inv i_31185(.A(nbus_14541[29]), .Z(n_31197));
	notech_inv i_31186(.A(nbus_14541[30]), .Z(n_31198));
	notech_inv i_31187(.A(nbus_14541[31]), .Z(n_31199));
	notech_inv i_31188(.A(cr2_reg[0]), .Z(n_31200));
	notech_inv i_31189(.A(cr2_reg[1]), .Z(n_31201));
	notech_inv i_31190(.A(cr2_reg[2]), .Z(n_31202));
	notech_inv i_31191(.A(cr2_reg[3]), .Z(n_31203));
	notech_inv i_31193(.A(cr2_reg[4]), .Z(n_31204));
	notech_inv i_31194(.A(cr2_reg[6]), .Z(n_31205));
	notech_inv i_31195(.A(cr2_reg[7]), .Z(n_31206));
	notech_inv i_31196(.A(cr2_reg[8]), .Z(n_31207));
	notech_inv i_31197(.A(cr2_reg[9]), .Z(n_31208));
	notech_inv i_31198(.A(cr2_reg[10]), .Z(n_31209));
	notech_inv i_31199(.A(cr2_reg[11]), .Z(n_31210));
	notech_inv i_31200(.A(cr2_reg[12]), .Z(n_31211));
	notech_inv i_31201(.A(cr2_reg[13]), .Z(n_31212));
	notech_inv i_31202(.A(cr2_reg[14]), .Z(n_31213));
	notech_inv i_31203(.A(cr2_reg[15]), .Z(n_31214));
	notech_inv i_31204(.A(cr2_reg[16]), .Z(n_31215));
	notech_inv i_31205(.A(cr2_reg[21]), .Z(n_31216));
	notech_inv i_31206(.A(\nbus_14540[0] ), .Z(n_31217));
	notech_inv i_31207(.A(\nbus_14540[1] ), .Z(n_31219));
	notech_inv i_31209(.A(\nbus_14540[2] ), .Z(n_31221));
	notech_inv i_31210(.A(\nbus_14540[3] ), .Z(n_31222));
	notech_inv i_31211(.A(\nbus_14540[4] ), .Z(n_31223));
	notech_inv i_31212(.A(\nbus_14540[5] ), .Z(n_31224));
	notech_inv i_31213(.A(\nbus_14540[6] ), .Z(n_31225));
	notech_inv i_31214(.A(\nbus_14540[7] ), .Z(n_31226));
	notech_inv i_31215(.A(\nbus_14540[8] ), .Z(n_31227));
	notech_inv i_31216(.A(\nbus_14540[9] ), .Z(n_31228));
	notech_inv i_31217(.A(\nbus_14540[10] ), .Z(n_31229));
	notech_inv i_31218(.A(\nbus_14540[11] ), .Z(n_31230));
	notech_inv i_31219(.A(n_17048), .Z(n_31231));
	notech_inv i_31220(.A(n_17054), .Z(n_31233));
	notech_inv i_31221(.A(n_17060), .Z(n_31234));
	notech_inv i_31222(.A(n_17066), .Z(n_31235));
	notech_inv i_31223(.A(n_17072), .Z(n_31236));
	notech_inv i_31224(.A(n_17084), .Z(n_31237));
	notech_inv i_31225(.A(n_17090), .Z(n_31238));
	notech_inv i_31226(.A(\nbus_11337[0] ), .Z(n_31239));
	notech_inv i_31227(.A(n_17096), .Z(n_31240));
	notech_inv i_31228(.A(n_17102), .Z(n_31241));
	notech_inv i_31229(.A(n_17108), .Z(n_31242));
	notech_inv i_31230(.A(n_17114), .Z(n_31243));
	notech_inv i_31231(.A(n_17120), .Z(n_31244));
	notech_inv i_31232(.A(n_17126), .Z(n_31245));
	notech_inv i_31233(.A(n_17132), .Z(n_31246));
	notech_inv i_31234(.A(n_17138), .Z(n_31247));
	notech_inv i_31235(.A(\nbus_11337[16] ), .Z(n_31248));
	notech_inv i_31236(.A(tcmp), .Z(n_31249));
	notech_inv i_31237(.A(n_18288), .Z(n_31250));
	notech_inv i_31238(.A(n_61898), .Z(n_31251));
	notech_inv i_31239(.A(fsm[2]), .Z(n_31252));
	notech_inv i_31241(.A(n_13955), .Z(n_31253));
	notech_inv i_31242(.A(fsm[3]), .Z(n_31254));
	notech_inv i_31243(.A(n_13961), .Z(n_31255));
	notech_inv i_31244(.A(vliw_pc[0]), .Z(n_31256));
	notech_inv i_31245(.A(vliw_pc[3]), .Z(n_31257));
	notech_inv i_31246(.A(vliw_pc[4]), .Z(n_31258));
	notech_inv i_31247(.A(n_21312), .Z(n_31259));
	notech_inv i_31248(.A(\nbus_11355[0] ), .Z(n_31260));
	notech_inv i_31249(.A(temp_ss[0]), .Z(n_31261));
	notech_inv i_31250(.A(temp_ss[1]), .Z(n_31262));
	notech_inv i_31251(.A(temp_ss[2]), .Z(n_31263));
	notech_inv i_31252(.A(temp_ss[3]), .Z(n_31264));
	notech_inv i_31253(.A(temp_ss[4]), .Z(n_31265));
	notech_inv i_31254(.A(temp_ss[5]), .Z(n_31266));
	notech_inv i_31255(.A(temp_ss[6]), .Z(n_31267));
	notech_inv i_31257(.A(temp_ss[7]), .Z(n_31268));
	notech_inv i_31258(.A(temp_ss[8]), .Z(n_31269));
	notech_inv i_31259(.A(temp_ss[9]), .Z(n_31270));
	notech_inv i_31260(.A(temp_ss[10]), .Z(n_31271));
	notech_inv i_31261(.A(temp_ss[11]), .Z(n_31272));
	notech_inv i_31262(.A(temp_ss[12]), .Z(n_31273));
	notech_inv i_31264(.A(temp_ss[13]), .Z(n_31274));
	notech_inv i_31265(.A(temp_ss[14]), .Z(n_31275));
	notech_inv i_31267(.A(temp_ss[15]), .Z(n_31276));
	notech_inv i_31268(.A(temp_ss[16]), .Z(n_31277));
	notech_inv i_31269(.A(temp_ss[17]), .Z(n_31278));
	notech_inv i_31270(.A(temp_ss[18]), .Z(n_31279));
	notech_inv i_31271(.A(temp_ss[19]), .Z(n_31280));
	notech_inv i_31272(.A(temp_ss[20]), .Z(n_31281));
	notech_inv i_31273(.A(temp_ss[21]), .Z(n_31282));
	notech_inv i_31275(.A(temp_ss[22]), .Z(n_31283));
	notech_inv i_31276(.A(temp_ss[23]), .Z(n_31284));
	notech_inv i_31277(.A(temp_ss[24]), .Z(n_31285));
	notech_inv i_31279(.A(temp_ss[25]), .Z(n_31286));
	notech_inv i_31280(.A(temp_ss[26]), .Z(n_31287));
	notech_inv i_31281(.A(temp_ss[27]), .Z(n_31288));
	notech_inv i_31282(.A(temp_ss[28]), .Z(n_31289));
	notech_inv i_31283(.A(temp_ss[29]), .Z(n_31290));
	notech_inv i_31284(.A(temp_ss[30]), .Z(n_31291));
	notech_inv i_31285(.A(temp_ss[31]), .Z(n_31292));
	notech_inv i_31286(.A(\nbus_11345[0] ), .Z(n_31293));
	notech_inv i_31287(.A(errco[0]), .Z(n_31294));
	notech_inv i_31288(.A(errco[1]), .Z(n_31295));
	notech_inv i_31289(.A(errco[2]), .Z(n_31296));
	notech_inv i_31290(.A(errco[3]), .Z(n_31297));
	notech_inv i_31291(.A(errco[4]), .Z(n_31298));
	notech_inv i_31292(.A(errco[5]), .Z(n_31299));
	notech_inv i_31293(.A(errco[6]), .Z(n_31300));
	notech_inv i_31296(.A(errco[7]), .Z(n_31301));
	notech_inv i_31297(.A(errco[8]), .Z(n_31302));
	notech_inv i_31298(.A(errco[9]), .Z(n_31303));
	notech_inv i_31299(.A(errco[10]), .Z(n_31304));
	notech_inv i_31300(.A(errco[11]), .Z(n_31305));
	notech_inv i_31301(.A(errco[12]), .Z(n_31306));
	notech_inv i_31302(.A(errco[13]), .Z(n_31307));
	notech_inv i_31303(.A(errco[14]), .Z(n_31308));
	notech_inv i_31304(.A(errco[15]), .Z(n_31309));
	notech_inv i_31305(.A(errco[16]), .Z(n_31310));
	notech_inv i_31306(.A(errco[17]), .Z(n_31311));
	notech_inv i_31307(.A(errco[18]), .Z(n_31312));
	notech_inv i_31308(.A(errco[19]), .Z(n_31313));
	notech_inv i_31310(.A(errco[20]), .Z(n_31314));
	notech_inv i_31311(.A(errco[21]), .Z(n_31315));
	notech_inv i_31312(.A(errco[22]), .Z(n_31316));
	notech_inv i_31313(.A(errco[23]), .Z(n_31317));
	notech_inv i_31314(.A(errco[24]), .Z(n_31318));
	notech_inv i_31315(.A(errco[25]), .Z(n_31319));
	notech_inv i_31317(.A(errco[26]), .Z(n_31320));
	notech_inv i_31318(.A(errco[27]), .Z(n_31321));
	notech_inv i_31319(.A(errco[28]), .Z(n_31322));
	notech_inv i_31320(.A(errco[29]), .Z(n_31323));
	notech_inv i_31321(.A(errco[30]), .Z(n_31324));
	notech_inv i_31322(.A(errco[31]), .Z(n_31325));
	notech_inv i_31323(.A(\nbus_11354[0] ), .Z(n_31326));
	notech_inv i_31324(.A(n_1862), .Z(n_31327));
	notech_inv i_31325(.A(Daddrgs[0]), .Z(n_31328));
	notech_inv i_31326(.A(Daddrgs[1]), .Z(n_31329));
	notech_inv i_31327(.A(Daddrgs[2]), .Z(n_31330));
	notech_inv i_31328(.A(Daddrgs[3]), .Z(n_31331));
	notech_inv i_31329(.A(Daddrgs[4]), .Z(n_31332));
	notech_inv i_31330(.A(Daddrgs[5]), .Z(n_31333));
	notech_inv i_31331(.A(Daddrgs[6]), .Z(n_31334));
	notech_inv i_31332(.A(Daddrgs[7]), .Z(n_31335));
	notech_inv i_31333(.A(Daddrgs[8]), .Z(n_31336));
	notech_inv i_31334(.A(Daddrgs[9]), .Z(n_31337));
	notech_inv i_31335(.A(Daddrgs[10]), .Z(n_31338));
	notech_inv i_31336(.A(Daddrgs[11]), .Z(n_31339));
	notech_inv i_31337(.A(Daddrgs[12]), .Z(n_31340));
	notech_inv i_31338(.A(Daddrgs[13]), .Z(n_31341));
	notech_inv i_31339(.A(Daddrgs[14]), .Z(n_31342));
	notech_inv i_31340(.A(Daddrgs[15]), .Z(n_31343));
	notech_inv i_31341(.A(Daddrgs[16]), .Z(n_31344));
	notech_inv i_31342(.A(Daddrgs[17]), .Z(n_31345));
	notech_inv i_31343(.A(Daddrgs[18]), .Z(n_31346));
	notech_inv i_31344(.A(Daddrgs[19]), .Z(n_31347));
	notech_inv i_31345(.A(Daddrgs[20]), .Z(n_31348));
	notech_inv i_31346(.A(Daddrgs[21]), .Z(n_31349));
	notech_inv i_31347(.A(Daddrgs[22]), .Z(n_31350));
	notech_inv i_31348(.A(Daddrgs[23]), .Z(n_31351));
	notech_inv i_31349(.A(Daddrgs[24]), .Z(n_31352));
	notech_inv i_31350(.A(Daddrgs[25]), .Z(n_31353));
	notech_inv i_31351(.A(Daddrgs[26]), .Z(n_31354));
	notech_inv i_31352(.A(Daddrgs[27]), .Z(n_31355));
	notech_inv i_31353(.A(Daddrgs[28]), .Z(n_31356));
	notech_inv i_31354(.A(Daddrgs[29]), .Z(n_31357));
	notech_inv i_31355(.A(Daddrgs[30]), .Z(n_31358));
	notech_inv i_31356(.A(Daddrgs[31]), .Z(n_31359));
	notech_inv i_31357(.A(n_18354), .Z(n_31360));
	notech_inv i_31358(.A(n_16862), .Z(n_31361));
	notech_inv i_31359(.A(n_171360317), .Z(n_31362));
	notech_inv i_31360(.A(n_164496008), .Z(n_31363));
	notech_inv i_31361(.A(n_9190), .Z(n_31364));
	notech_inv i_31362(.A(n_61661), .Z(n_31365));
	notech_inv i_31363(.A(n_7469), .Z(n_31366));
	notech_inv i_31364(.A(cs[0]), .Z(n_31367));
	notech_inv i_31365(.A(cs[1]), .Z(n_31368));
	notech_inv i_31366(.A(all_cnt[0]), .Z(n_31369));
	notech_inv i_31367(.A(all_cnt[1]), .Z(n_31370));
	notech_inv i_31368(.A(all_cnt[2]), .Z(n_31371));
	notech_inv i_31369(.A(all_cnt[3]), .Z(n_31372));
	notech_inv i_31370(.A(calc_sz[0]), .Z(n_31373));
	notech_inv i_31371(.A(calc_sz[2]), .Z(n_31374));
	notech_inv i_31372(.A(n_60953), .Z(nbus_11273[0]));
	notech_inv i_31373(.A(opa[1]), .Z(nbus_11273[1]));
	notech_inv i_31374(.A(n_60962), .Z(nbus_11273[2]));
	notech_inv i_31375(.A(n_60971), .Z(nbus_11273[3]));
	notech_inv i_31376(.A(opa[4]), .Z(nbus_11273[4]));
	notech_inv i_31377(.A(n_60980), .Z(nbus_11273[5]));
	notech_inv i_31378(.A(n_60989), .Z(nbus_11273[6]));
	notech_inv i_31379(.A(n_60998), .Z(nbus_11273[7]));
	notech_inv i_31380(.A(opa[8]), .Z(nbus_11273[8]));
	notech_inv i_31381(.A(n_61007), .Z(nbus_11273[9]));
	notech_inv i_31382(.A(opa[10]), .Z(nbus_11273[10]));
	notech_inv i_31383(.A(opa[11]), .Z(nbus_11273[11]));
	notech_inv i_31384(.A(n_61016), .Z(nbus_11273[12]));
	notech_inv i_31385(.A(n_61025), .Z(nbus_11273[13]));
	notech_inv i_31386(.A(opa[14]), .Z(nbus_11273[14]));
	notech_inv i_31387(.A(n_61034), .Z(nbus_11273[15]));
	notech_inv i_31388(.A(opa[16]), .Z(\nbus_11283[16] ));
	notech_inv i_31389(.A(opa[17]), .Z(\nbus_11283[17] ));
	notech_inv i_31391(.A(opa[18]), .Z(\nbus_11283[18] ));
	notech_inv i_31392(.A(opa[19]), .Z(\nbus_11283[19] ));
	notech_inv i_31393(.A(opa[20]), .Z(\nbus_11283[20] ));
	notech_inv i_31394(.A(opa[21]), .Z(\nbus_11283[21] ));
	notech_inv i_31398(.A(opa[22]), .Z(\nbus_11283[22] ));
	notech_inv i_31399(.A(opa[23]), .Z(\nbus_11283[23] ));
	notech_inv i_31401(.A(opa[24]), .Z(\nbus_11283[24] ));
	notech_inv i_31402(.A(opa[25]), .Z(\nbus_11283[25] ));
	notech_inv i_31403(.A(opa[26]), .Z(\nbus_11283[26] ));
	notech_inv i_31404(.A(opa[27]), .Z(\nbus_11283[27] ));
	notech_inv i_31405(.A(opa[28]), .Z(\nbus_11283[28] ));
	notech_inv i_31406(.A(opa[29]), .Z(\nbus_11283[29] ));
	notech_inv i_31407(.A(opa[30]), .Z(\nbus_11283[30] ));
	notech_inv i_31408(.A(opa[31]), .Z(\nbus_11283[31] ));
	notech_inv i_31409(.A(reps[2]), .Z(n_31407));
	notech_inv i_31411(.A(ecx[0]), .Z(n_31408));
	notech_inv i_31412(.A(ecx[1]), .Z(n_31409));
	notech_inv i_31413(.A(ecx[2]), .Z(n_31410));
	notech_inv i_31414(.A(ecx[3]), .Z(n_31411));
	notech_inv i_31415(.A(ecx[4]), .Z(n_31412));
	notech_inv i_31418(.A(ecx[5]), .Z(n_31413));
	notech_inv i_31419(.A(ecx[6]), .Z(n_31414));
	notech_inv i_31420(.A(ecx[7]), .Z(n_31415));
	notech_inv i_31421(.A(ecx[8]), .Z(n_31416));
	notech_inv i_31423(.A(ecx[9]), .Z(n_31417));
	notech_inv i_31424(.A(ecx[10]), .Z(n_31418));
	notech_inv i_31426(.A(ecx[11]), .Z(n_31419));
	notech_inv i_31427(.A(ecx[12]), .Z(n_31420));
	notech_inv i_31428(.A(ecx[13]), .Z(n_31421));
	notech_inv i_31430(.A(ecx[14]), .Z(n_31422));
	notech_inv i_31431(.A(ecx[15]), .Z(n_31423));
	notech_inv i_31432(.A(ecx[16]), .Z(n_31424));
	notech_inv i_31433(.A(ecx[17]), .Z(n_31425));
	notech_inv i_31435(.A(ecx[18]), .Z(n_31426));
	notech_inv i_31436(.A(ecx[19]), .Z(n_31427));
	notech_inv i_31437(.A(ecx[20]), .Z(n_31428));
	notech_inv i_31438(.A(ecx[21]), .Z(n_31429));
	notech_inv i_31439(.A(ecx[22]), .Z(n_31430));
	notech_inv i_31440(.A(ecx[23]), .Z(n_31431));
	notech_inv i_31441(.A(ecx[24]), .Z(n_31432));
	notech_inv i_31442(.A(ecx[25]), .Z(n_31433));
	notech_inv i_31443(.A(ecx[26]), .Z(n_31434));
	notech_inv i_31444(.A(ecx[27]), .Z(n_31435));
	notech_inv i_31445(.A(ecx[28]), .Z(n_31436));
	notech_inv i_31446(.A(ecx[29]), .Z(n_31437));
	notech_inv i_31447(.A(ecx[30]), .Z(n_31438));
	notech_inv i_31448(.A(ecx[31]), .Z(n_31439));
	notech_inv i_31449(.A(opb[0]), .Z(\nbus_11290[0] ));
	notech_inv i_31450(.A(opb[1]), .Z(\nbus_11290[1] ));
	notech_inv i_31451(.A(opb[2]), .Z(\nbus_11290[2] ));
	notech_inv i_31452(.A(opb[3]), .Z(\nbus_11290[3] ));
	notech_inv i_31453(.A(opb[4]), .Z(\nbus_11290[4] ));
	notech_inv i_31454(.A(opb[5]), .Z(\nbus_11290[5] ));
	notech_inv i_31455(.A(opb[6]), .Z(\nbus_11290[6] ));
	notech_inv i_31456(.A(opb[7]), .Z(\nbus_11290[7] ));
	notech_inv i_31457(.A(opb[8]), .Z(\nbus_11290[8] ));
	notech_inv i_31458(.A(opb[9]), .Z(\nbus_11290[9] ));
	notech_inv i_31459(.A(opb[10]), .Z(\nbus_11290[10] ));
	notech_inv i_31460(.A(opb[11]), .Z(\nbus_11290[11] ));
	notech_inv i_31461(.A(opb[12]), .Z(\nbus_11290[12] ));
	notech_inv i_31462(.A(opb[13]), .Z(\nbus_11290[13] ));
	notech_inv i_31463(.A(opb[14]), .Z(\nbus_11290[14] ));
	notech_inv i_31464(.A(opb[15]), .Z(\nbus_11290[15] ));
	notech_inv i_31465(.A(opb[16]), .Z(\nbus_11290[16] ));
	notech_inv i_31467(.A(opb[17]), .Z(\nbus_11290[17] ));
	notech_inv i_31468(.A(opb[18]), .Z(\nbus_11290[18] ));
	notech_inv i_31469(.A(opb[19]), .Z(\nbus_11290[19] ));
	notech_inv i_31470(.A(opb[20]), .Z(\nbus_11290[20] ));
	notech_inv i_31471(.A(opb[21]), .Z(\nbus_11290[21] ));
	notech_inv i_31472(.A(opb[22]), .Z(\nbus_11290[22] ));
	notech_inv i_31473(.A(opb[23]), .Z(\nbus_11290[23] ));
	notech_inv i_31474(.A(opb[24]), .Z(\nbus_11290[24] ));
	notech_inv i_31475(.A(opb[25]), .Z(\nbus_11290[25] ));
	notech_inv i_31476(.A(opb[26]), .Z(\nbus_11290[26] ));
	notech_inv i_31477(.A(opb[27]), .Z(\nbus_11290[27] ));
	notech_inv i_31478(.A(opb[28]), .Z(\nbus_11290[28] ));
	notech_inv i_31479(.A(opb[29]), .Z(\nbus_11290[29] ));
	notech_inv i_31480(.A(opb[30]), .Z(\nbus_11290[30] ));
	notech_inv i_31481(.A(n_60629), .Z(\nbus_11290[31] ));
	notech_inv i_31482(.A(opd[0]), .Z(n_31472));
	notech_inv i_31483(.A(opd[1]), .Z(n_31473));
	notech_inv i_31484(.A(opd[2]), .Z(n_31474));
	notech_inv i_31486(.A(opd[3]), .Z(n_31476));
	notech_inv i_31487(.A(opd[4]), .Z(n_31477));
	notech_inv i_31488(.A(opd[5]), .Z(n_31478));
	notech_inv i_31490(.A(opd[6]), .Z(n_31479));
	notech_inv i_31491(.A(opd[7]), .Z(n_31480));
	notech_inv i_31492(.A(opd[8]), .Z(n_31481));
	notech_inv i_31493(.A(opd[9]), .Z(n_31482));
	notech_inv i_31494(.A(opd[10]), .Z(n_31483));
	notech_inv i_31495(.A(opd[11]), .Z(n_31484));
	notech_inv i_31496(.A(opd[12]), .Z(n_31485));
	notech_inv i_31497(.A(opd[13]), .Z(n_31486));
	notech_inv i_31498(.A(opd[14]), .Z(n_31487));
	notech_inv i_31499(.A(opd[15]), .Z(n_31488));
	notech_inv i_31500(.A(opd[16]), .Z(n_31489));
	notech_inv i_31501(.A(opd[17]), .Z(n_31490));
	notech_inv i_31502(.A(opd[18]), .Z(n_31491));
	notech_inv i_31503(.A(opd[19]), .Z(n_31492));
	notech_inv i_31504(.A(opd[20]), .Z(n_31493));
	notech_inv i_31505(.A(opd[21]), .Z(n_31494));
	notech_inv i_31506(.A(opd[22]), .Z(n_31496));
	notech_inv i_31507(.A(opd[23]), .Z(n_31499));
	notech_inv i_31508(.A(opd[24]), .Z(n_31500));
	notech_inv i_31509(.A(opd[25]), .Z(n_31501));
	notech_inv i_31510(.A(n_57965), .Z(n_31502));
	notech_inv i_31511(.A(n_57956), .Z(n_31503));
	notech_inv i_31512(.A(n_57946), .Z(n_31504));
	notech_inv i_31513(.A(n_57937), .Z(n_31505));
	notech_inv i_31514(.A(opd[30]), .Z(n_31506));
	notech_inv i_31515(.A(n_58018), .Z(n_31507));
	notech_inv i_31516(.A(read_data[0]), .Z(n_31508));
	notech_inv i_31517(.A(read_data[1]), .Z(n_31509));
	notech_inv i_31518(.A(read_data[2]), .Z(n_31510));
	notech_inv i_31519(.A(read_data[3]), .Z(n_31511));
	notech_inv i_31520(.A(read_data[4]), .Z(n_31512));
	notech_inv i_31521(.A(read_data[5]), .Z(n_31513));
	notech_inv i_31522(.A(read_data[6]), .Z(n_31514));
	notech_inv i_31523(.A(read_data[7]), .Z(n_31515));
	notech_inv i_31524(.A(read_data[8]), .Z(n_31516));
	notech_inv i_31525(.A(read_data[9]), .Z(n_31517));
	notech_inv i_31526(.A(read_data[10]), .Z(n_31518));
	notech_inv i_31527(.A(read_data[11]), .Z(n_31519));
	notech_inv i_31528(.A(read_data[12]), .Z(n_31520));
	notech_inv i_31529(.A(read_data[13]), .Z(n_31521));
	notech_inv i_31530(.A(read_data[14]), .Z(n_31522));
	notech_inv i_31531(.A(read_data[15]), .Z(n_31523));
	notech_inv i_31532(.A(read_data[16]), .Z(n_31524));
	notech_inv i_31533(.A(read_data[17]), .Z(n_31525));
	notech_inv i_31534(.A(read_data[18]), .Z(n_31526));
	notech_inv i_31535(.A(read_data[19]), .Z(n_31527));
	notech_inv i_31536(.A(read_data[20]), .Z(n_31528));
	notech_inv i_31537(.A(read_data[21]), .Z(n_31529));
	notech_inv i_31538(.A(read_data[22]), .Z(n_31530));
	notech_inv i_31539(.A(read_data[23]), .Z(n_31531));
	notech_inv i_31540(.A(read_data[24]), .Z(n_31532));
	notech_inv i_31541(.A(read_data[25]), .Z(n_31533));
	notech_inv i_31542(.A(read_data[26]), .Z(n_31534));
	notech_inv i_31543(.A(read_data[27]), .Z(n_31535));
	notech_inv i_31544(.A(read_data[28]), .Z(n_31536));
	notech_inv i_31545(.A(read_data[29]), .Z(n_31537));
	notech_inv i_31546(.A(read_data[30]), .Z(n_31538));
	notech_inv i_31547(.A(read_data[31]), .Z(n_31539));
	notech_inv i_31548(.A(opc[0]), .Z(nbus_11271[0]));
	notech_inv i_31549(.A(opc[1]), .Z(nbus_11271[1]));
	notech_inv i_31550(.A(opc[2]), .Z(nbus_11271[2]));
	notech_inv i_31551(.A(opc[3]), .Z(nbus_11271[3]));
	notech_inv i_31552(.A(opc[4]), .Z(nbus_11271[4]));
	notech_inv i_31553(.A(opc[5]), .Z(nbus_11271[5]));
	notech_inv i_31554(.A(opc[6]), .Z(nbus_11271[6]));
	notech_inv i_31555(.A(opc[7]), .Z(nbus_11271[7]));
	notech_inv i_31556(.A(opc[8]), .Z(nbus_11271[8]));
	notech_inv i_31557(.A(opc[9]), .Z(nbus_11271[9]));
	notech_inv i_31558(.A(opc[10]), .Z(nbus_11271[10]));
	notech_inv i_31559(.A(opc[11]), .Z(nbus_11271[11]));
	notech_inv i_31560(.A(opc[12]), .Z(nbus_11271[12]));
	notech_inv i_31561(.A(opc[13]), .Z(nbus_11271[13]));
	notech_inv i_31562(.A(opc[14]), .Z(nbus_11271[14]));
	notech_inv i_31563(.A(opc[15]), .Z(nbus_11271[15]));
	notech_inv i_31564(.A(opc[16]), .Z(nbus_11271[16]));
	notech_inv i_31565(.A(opc[17]), .Z(nbus_11271[17]));
	notech_inv i_31566(.A(opc[18]), .Z(nbus_11271[18]));
	notech_inv i_31567(.A(opc[19]), .Z(nbus_11271[19]));
	notech_inv i_31568(.A(opc[20]), .Z(nbus_11271[20]));
	notech_inv i_31569(.A(opc[21]), .Z(nbus_11271[21]));
	notech_inv i_31570(.A(opc[22]), .Z(nbus_11271[22]));
	notech_inv i_31571(.A(opc[23]), .Z(nbus_11271[23]));
	notech_inv i_31573(.A(opc[24]), .Z(nbus_11271[24]));
	notech_inv i_31574(.A(opc[25]), .Z(nbus_11271[25]));
	notech_inv i_31575(.A(opc[26]), .Z(nbus_11271[26]));
	notech_inv i_31576(.A(opc[27]), .Z(nbus_11271[27]));
	notech_inv i_31577(.A(opc[28]), .Z(nbus_11271[28]));
	notech_inv i_31578(.A(opc[29]), .Z(nbus_11271[29]));
	notech_inv i_31579(.A(opc[30]), .Z(nbus_11271[30]));
	notech_inv i_31580(.A(n_60602), .Z(nbus_11271[31]));
	notech_inv i_31581(.A(regs_14[0]), .Z(n_31572));
	notech_inv i_31582(.A(regs_14[1]), .Z(n_31573));
	notech_inv i_31583(.A(regs_14[2]), .Z(n_31574));
	notech_inv i_31585(.A(regs_14[3]), .Z(n_31575));
	notech_inv i_31586(.A(regs_14[4]), .Z(n_31576));
	notech_inv i_31587(.A(regs_14[5]), .Z(n_31577));
	notech_inv i_31588(.A(regs_14[6]), .Z(n_31578));
	notech_inv i_31589(.A(regs_14[7]), .Z(n_31579));
	notech_inv i_31590(.A(regs_14[8]), .Z(n_31580));
	notech_inv i_31591(.A(regs_14[9]), .Z(n_31581));
	notech_inv i_31592(.A(regs_14[10]), .Z(n_31582));
	notech_inv i_31593(.A(regs_14[11]), .Z(n_31583));
	notech_inv i_31594(.A(regs_14[12]), .Z(n_31584));
	notech_inv i_31595(.A(regs_14[13]), .Z(n_31585));
	notech_inv i_31596(.A(regs_14[14]), .Z(n_31586));
	notech_inv i_31597(.A(regs_14[15]), .Z(n_31587));
	notech_inv i_31598(.A(regs_14[16]), .Z(n_31588));
	notech_inv i_31599(.A(regs_14[17]), .Z(n_31589));
	notech_inv i_31600(.A(regs_14[18]), .Z(n_31590));
	notech_inv i_31601(.A(regs_14[19]), .Z(n_31591));
	notech_inv i_31602(.A(regs_14[20]), .Z(n_31592));
	notech_inv i_31603(.A(regs_14[21]), .Z(n_31593));
	notech_inv i_31604(.A(regs_14[22]), .Z(n_31594));
	notech_inv i_31605(.A(regs_14[23]), .Z(n_31595));
	notech_inv i_31606(.A(regs_14[24]), .Z(n_31596));
	notech_inv i_31607(.A(regs_14[25]), .Z(n_31597));
	notech_inv i_31608(.A(regs_14[26]), .Z(n_31598));
	notech_inv i_31609(.A(regs_14[27]), .Z(n_31599));
	notech_inv i_31610(.A(regs_14[28]), .Z(n_31600));
	notech_inv i_31611(.A(regs_14[29]), .Z(n_31601));
	notech_inv i_31612(.A(regs_14[30]), .Z(n_31602));
	notech_inv i_31613(.A(regs_14[31]), .Z(n_31603));
	notech_inv i_31614(.A(opz[0]), .Z(n_31604));
	notech_inv i_31615(.A(opz[1]), .Z(n_31605));
	notech_inv i_31616(.A(opz[2]), .Z(n_31606));
	notech_inv i_31617(.A(cr3[12]), .Z(n_31607));
	notech_inv i_31618(.A(cr3[13]), .Z(n_31608));
	notech_inv i_31619(.A(cr3[14]), .Z(n_31609));
	notech_inv i_31620(.A(cr3[15]), .Z(n_31610));
	notech_inv i_31621(.A(opc_10[0]), .Z(n_31611));
	notech_inv i_31622(.A(opc_10[1]), .Z(n_31612));
	notech_inv i_31623(.A(opc_10[2]), .Z(n_31613));
	notech_inv i_31624(.A(opc_10[3]), .Z(n_31614));
	notech_inv i_31625(.A(opc_10[4]), .Z(n_31615));
	notech_inv i_31626(.A(opc_10[5]), .Z(n_31616));
	notech_inv i_31627(.A(opc_10[6]), .Z(n_31617));
	notech_inv i_31628(.A(opc_10[7]), .Z(n_31618));
	notech_inv i_31629(.A(opc_10[8]), .Z(n_31619));
	notech_inv i_31630(.A(opc_10[9]), .Z(n_31620));
	notech_inv i_31631(.A(opc_10[10]), .Z(n_31621));
	notech_inv i_31632(.A(opc_10[11]), .Z(n_31622));
	notech_inv i_31633(.A(opc_10[12]), .Z(n_31623));
	notech_inv i_31634(.A(opc_10[13]), .Z(n_31624));
	notech_inv i_31636(.A(opc_10[14]), .Z(n_31625));
	notech_inv i_31637(.A(opc_10[15]), .Z(n_31626));
	notech_inv i_31638(.A(opc_10[16]), .Z(n_31627));
	notech_inv i_31639(.A(opc_10[17]), .Z(n_31628));
	notech_inv i_31640(.A(opc_10[18]), .Z(n_31629));
	notech_inv i_31641(.A(opc_10[19]), .Z(n_31630));
	notech_inv i_31642(.A(opc_10[20]), .Z(n_31631));
	notech_inv i_31643(.A(opc_10[21]), .Z(n_31632));
	notech_inv i_31646(.A(opc_10[22]), .Z(n_31633));
	notech_inv i_31647(.A(opc_10[23]), .Z(n_31634));
	notech_inv i_31648(.A(opc_10[24]), .Z(n_31635));
	notech_inv i_31649(.A(opc_10[25]), .Z(n_31636));
	notech_inv i_31651(.A(opc_10[26]), .Z(n_31637));
	notech_inv i_31652(.A(opc_10[27]), .Z(n_31638));
	notech_inv i_31654(.A(opc_10[28]), .Z(n_31639));
	notech_inv i_31655(.A(opc_10[29]), .Z(n_31640));
	notech_inv i_31656(.A(opc_10[30]), .Z(n_31641));
	notech_inv i_31657(.A(opc_10[31]), .Z(n_31642));
	notech_inv i_31658(.A(regs_6[0]), .Z(n_31643));
	notech_inv i_31659(.A(regs_6[1]), .Z(n_31644));
	notech_inv i_31660(.A(regs_6[2]), .Z(n_31645));
	notech_inv i_31661(.A(regs_6[3]), .Z(n_31646));
	notech_inv i_31662(.A(regs_6[4]), .Z(n_31647));
	notech_inv i_31663(.A(regs_6[5]), .Z(n_31648));
	notech_inv i_31664(.A(regs_6[6]), .Z(n_31649));
	notech_inv i_31665(.A(regs_6[7]), .Z(n_31650));
	notech_inv i_31666(.A(regs_6[8]), .Z(n_31651));
	notech_inv i_31667(.A(regs_6[9]), .Z(n_31652));
	notech_inv i_31668(.A(regs_6[10]), .Z(n_31653));
	notech_inv i_31669(.A(regs_6[11]), .Z(n_31654));
	notech_inv i_31670(.A(regs_6[12]), .Z(n_31655));
	notech_inv i_31671(.A(regs_6[13]), .Z(n_31656));
	notech_inv i_31672(.A(regs_6[14]), .Z(n_31657));
	notech_inv i_31673(.A(regs_6[15]), .Z(n_31658));
	notech_inv i_31674(.A(regs_6[16]), .Z(n_31659));
	notech_inv i_31675(.A(regs_6[17]), .Z(n_31660));
	notech_inv i_31676(.A(regs_6[18]), .Z(n_31661));
	notech_inv i_31677(.A(regs_6[19]), .Z(n_31662));
	notech_inv i_31678(.A(regs_6[20]), .Z(n_31663));
	notech_inv i_31679(.A(regs_6[21]), .Z(n_31664));
	notech_inv i_31680(.A(regs_6[22]), .Z(n_31665));
	notech_inv i_31681(.A(regs_6[23]), .Z(n_31666));
	notech_inv i_31682(.A(regs_6[24]), .Z(n_31667));
	notech_inv i_31683(.A(regs_6[25]), .Z(n_31668));
	notech_inv i_31684(.A(regs_6[26]), .Z(n_31669));
	notech_inv i_31685(.A(regs_6[27]), .Z(n_31670));
	notech_inv i_31686(.A(regs_6[28]), .Z(n_31671));
	notech_inv i_31687(.A(regs_6[29]), .Z(n_31672));
	notech_inv i_31688(.A(regs_6[30]), .Z(n_31673));
	notech_inv i_31689(.A(regs_6[31]), .Z(n_31674));
	notech_inv i_31690(.A(regs_10[0]), .Z(n_31675));
	notech_inv i_31691(.A(regs_10[1]), .Z(n_31676));
	notech_inv i_31692(.A(regs_10[2]), .Z(n_31677));
	notech_inv i_31693(.A(regs_10[3]), .Z(n_31678));
	notech_inv i_31694(.A(regs_10[4]), .Z(n_31679));
	notech_inv i_31695(.A(regs_10[5]), .Z(n_31680));
	notech_inv i_31696(.A(regs_10[6]), .Z(n_31681));
	notech_inv i_31697(.A(regs_10[7]), .Z(n_31682));
	notech_inv i_31698(.A(regs_10[8]), .Z(n_31683));
	notech_inv i_31699(.A(regs_10[9]), .Z(n_31684));
	notech_inv i_31700(.A(regs_10[10]), .Z(n_31685));
	notech_inv i_31701(.A(regs_10[11]), .Z(n_31686));
	notech_inv i_31702(.A(regs_10[12]), .Z(n_31687));
	notech_inv i_31703(.A(regs_10[13]), .Z(n_31688));
	notech_inv i_31704(.A(regs_10[14]), .Z(n_31689));
	notech_inv i_31705(.A(regs_10[15]), .Z(n_31690));
	notech_inv i_31706(.A(regs_10[16]), .Z(n_31691));
	notech_inv i_31707(.A(regs_10[17]), .Z(n_31692));
	notech_inv i_31708(.A(regs_10[18]), .Z(n_31693));
	notech_inv i_31709(.A(regs_10[19]), .Z(n_31694));
	notech_inv i_31710(.A(regs_10[20]), .Z(n_31695));
	notech_inv i_31711(.A(regs_10[21]), .Z(n_31696));
	notech_inv i_31712(.A(regs_10[22]), .Z(n_31697));
	notech_inv i_31713(.A(regs_10[23]), .Z(n_31698));
	notech_inv i_31714(.A(regs_10[24]), .Z(n_31699));
	notech_inv i_31715(.A(regs_10[25]), .Z(n_31700));
	notech_inv i_31716(.A(regs_10[26]), .Z(n_31701));
	notech_inv i_31717(.A(regs_10[27]), .Z(n_31702));
	notech_inv i_31718(.A(regs_10[28]), .Z(n_31703));
	notech_inv i_31719(.A(regs_10[29]), .Z(n_31704));
	notech_inv i_31720(.A(regs_10[30]), .Z(n_31705));
	notech_inv i_31721(.A(regs_10[31]), .Z(n_31706));
	notech_inv i_31722(.A(regs_8[0]), .Z(n_31707));
	notech_inv i_31723(.A(regs_8[1]), .Z(n_31708));
	notech_inv i_31724(.A(regs_8[2]), .Z(n_31709));
	notech_inv i_31725(.A(regs_8[3]), .Z(n_31710));
	notech_inv i_31726(.A(regs_8[4]), .Z(n_31711));
	notech_inv i_31727(.A(regs_8[5]), .Z(n_31712));
	notech_inv i_31728(.A(regs_8[6]), .Z(n_31713));
	notech_inv i_31729(.A(regs_8[7]), .Z(n_31714));
	notech_inv i_31730(.A(regs_8[8]), .Z(n_31715));
	notech_inv i_31731(.A(regs_8[9]), .Z(n_31716));
	notech_inv i_31732(.A(regs_8[10]), .Z(n_31717));
	notech_inv i_31733(.A(regs_8[11]), .Z(n_31718));
	notech_inv i_31734(.A(regs_8[12]), .Z(n_31719));
	notech_inv i_31735(.A(regs_8[13]), .Z(n_31720));
	notech_inv i_31736(.A(regs_8[14]), .Z(n_31721));
	notech_inv i_31737(.A(regs_8[15]), .Z(n_31722));
	notech_inv i_31738(.A(regs_8[16]), .Z(n_31723));
	notech_inv i_31739(.A(regs_8[17]), .Z(n_31724));
	notech_inv i_31740(.A(regs_8[18]), .Z(n_31725));
	notech_inv i_31741(.A(regs_8[19]), .Z(n_31726));
	notech_inv i_31742(.A(regs_8[20]), .Z(n_31727));
	notech_inv i_31743(.A(regs_8[21]), .Z(n_31728));
	notech_inv i_31744(.A(regs_8[22]), .Z(n_31729));
	notech_inv i_31745(.A(regs_8[23]), .Z(n_31730));
	notech_inv i_31746(.A(regs_8[24]), .Z(n_31731));
	notech_inv i_31747(.A(regs_8[25]), .Z(n_31732));
	notech_inv i_31748(.A(regs_8[26]), .Z(n_31733));
	notech_inv i_31749(.A(regs_8[27]), .Z(n_31734));
	notech_inv i_31750(.A(regs_8[28]), .Z(n_31735));
	notech_inv i_31751(.A(regs_8[29]), .Z(n_31736));
	notech_inv i_31752(.A(regs_8[30]), .Z(n_31737));
	notech_inv i_31753(.A(regs_8[31]), .Z(n_31738));
	notech_inv i_31754(.A(regs_11[0]), .Z(n_31739));
	notech_inv i_31755(.A(regs_11[1]), .Z(n_31740));
	notech_inv i_31756(.A(regs_11[2]), .Z(n_31741));
	notech_inv i_31757(.A(regs_11[3]), .Z(n_31742));
	notech_inv i_31758(.A(regs_11[4]), .Z(n_31743));
	notech_inv i_31759(.A(regs_11[5]), .Z(n_31744));
	notech_inv i_31760(.A(regs_11[6]), .Z(n_31745));
	notech_inv i_31761(.A(regs_11[7]), .Z(n_31746));
	notech_inv i_31766(.A(regs_11[8]), .Z(n_31747));
	notech_inv i_31767(.A(regs_11[9]), .Z(n_31748));
	notech_inv i_31768(.A(regs_11[10]), .Z(n_31749));
	notech_inv i_31770(.A(regs_11[11]), .Z(n_31750));
	notech_inv i_31772(.A(regs_11[12]), .Z(n_31751));
	notech_inv i_31773(.A(regs_11[13]), .Z(n_31752));
	notech_inv i_31774(.A(regs_11[14]), .Z(n_31753));
	notech_inv i_31775(.A(regs_11[15]), .Z(n_31754));
	notech_inv i_31776(.A(regs_11[16]), .Z(n_31755));
	notech_inv i_31777(.A(regs_11[17]), .Z(n_31756));
	notech_inv i_31778(.A(regs_11[18]), .Z(n_31757));
	notech_inv i_31779(.A(regs_11[19]), .Z(n_31758));
	notech_inv i_31780(.A(regs_11[20]), .Z(n_31759));
	notech_inv i_31781(.A(regs_11[21]), .Z(n_31760));
	notech_inv i_31782(.A(regs_11[22]), .Z(n_31761));
	notech_inv i_31783(.A(regs_11[23]), .Z(n_31762));
	notech_inv i_31784(.A(regs_11[24]), .Z(n_31763));
	notech_inv i_31785(.A(regs_11[25]), .Z(n_31764));
	notech_inv i_31786(.A(regs_11[26]), .Z(n_31765));
	notech_inv i_31787(.A(regs_11[27]), .Z(n_31766));
	notech_inv i_31788(.A(regs_11[28]), .Z(n_31767));
	notech_inv i_31789(.A(regs_11[29]), .Z(n_31768));
	notech_inv i_31790(.A(regs_11[30]), .Z(n_31769));
	notech_inv i_31791(.A(regs_11[31]), .Z(n_31770));
	notech_inv i_31792(.A(regs_12[0]), .Z(n_31771));
	notech_inv i_31793(.A(regs_12[1]), .Z(n_31772));
	notech_inv i_31794(.A(regs_12[2]), .Z(n_31773));
	notech_inv i_31795(.A(regs_12[3]), .Z(n_31774));
	notech_inv i_31796(.A(regs_12[4]), .Z(n_31775));
	notech_inv i_31798(.A(regs_12[5]), .Z(n_31776));
	notech_inv i_31799(.A(regs_12[6]), .Z(n_31777));
	notech_inv i_31800(.A(regs_12[7]), .Z(n_31778));
	notech_inv i_31801(.A(regs_12[8]), .Z(n_31779));
	notech_inv i_31802(.A(regs_12[9]), .Z(n_31780));
	notech_inv i_31803(.A(regs_12[10]), .Z(n_31781));
	notech_inv i_31804(.A(regs_12[11]), .Z(n_31782));
	notech_inv i_31805(.A(regs_12[12]), .Z(n_31783));
	notech_inv i_31806(.A(regs_12[13]), .Z(n_31784));
	notech_inv i_31807(.A(regs_12[14]), .Z(n_31785));
	notech_inv i_31809(.A(regs_12[15]), .Z(n_31786));
	notech_inv i_31810(.A(regs_12[16]), .Z(n_31787));
	notech_inv i_31811(.A(regs_12[17]), .Z(n_31788));
	notech_inv i_31813(.A(regs_12[18]), .Z(n_31789));
	notech_inv i_31814(.A(regs_12[19]), .Z(n_31790));
	notech_inv i_31815(.A(regs_12[20]), .Z(n_31791));
	notech_inv i_31816(.A(regs_12[21]), .Z(n_31792));
	notech_inv i_31817(.A(regs_12[22]), .Z(n_31793));
	notech_inv i_31818(.A(regs_12[23]), .Z(n_31794));
	notech_inv i_31819(.A(regs_12[24]), .Z(n_31795));
	notech_inv i_31820(.A(regs_12[25]), .Z(n_31796));
	notech_inv i_31821(.A(regs_12[26]), .Z(n_31797));
	notech_inv i_31823(.A(regs_12[27]), .Z(n_31798));
	notech_inv i_31824(.A(regs_12[28]), .Z(n_31799));
	notech_inv i_31825(.A(regs_12[29]), .Z(n_31800));
	notech_inv i_31826(.A(regs_12[30]), .Z(n_31801));
	notech_inv i_31827(.A(regs_12[31]), .Z(n_31802));
	notech_inv i_31828(.A(regs_3[0]), .Z(n_31803));
	notech_inv i_31829(.A(regs_3[1]), .Z(n_31804));
	notech_inv i_31830(.A(regs_3[2]), .Z(n_31805));
	notech_inv i_31831(.A(regs_3[3]), .Z(n_31806));
	notech_inv i_31832(.A(regs_3[4]), .Z(n_31807));
	notech_inv i_31833(.A(regs_3[5]), .Z(n_31808));
	notech_inv i_31834(.A(regs_3[6]), .Z(n_31809));
	notech_inv i_31835(.A(regs_3[7]), .Z(n_31810));
	notech_inv i_31836(.A(regs_3[8]), .Z(n_31811));
	notech_inv i_31837(.A(regs_3[9]), .Z(n_31812));
	notech_inv i_31838(.A(regs_3[10]), .Z(n_31813));
	notech_inv i_31839(.A(regs_3[11]), .Z(n_31814));
	notech_inv i_31840(.A(regs_3[12]), .Z(n_31815));
	notech_inv i_31841(.A(regs_3[13]), .Z(n_31816));
	notech_inv i_31842(.A(regs_3[14]), .Z(n_31817));
	notech_inv i_31843(.A(regs_3[15]), .Z(n_31818));
	notech_inv i_31844(.A(regs_3[16]), .Z(n_31819));
	notech_inv i_31845(.A(regs_3[17]), .Z(n_31820));
	notech_inv i_31846(.A(regs_3[18]), .Z(n_31821));
	notech_inv i_31847(.A(regs_3[19]), .Z(n_31822));
	notech_inv i_31848(.A(regs_3[20]), .Z(n_31823));
	notech_inv i_31849(.A(regs_3[21]), .Z(n_31824));
	notech_inv i_31850(.A(regs_3[22]), .Z(n_31825));
	notech_inv i_31851(.A(regs_3[23]), .Z(n_31826));
	notech_inv i_31852(.A(regs_3[24]), .Z(n_31827));
	notech_inv i_31853(.A(regs_3[25]), .Z(n_31828));
	notech_inv i_31854(.A(regs_3[26]), .Z(n_31829));
	notech_inv i_31855(.A(regs_3[27]), .Z(n_31830));
	notech_inv i_31856(.A(regs_3[28]), .Z(n_31831));
	notech_inv i_31857(.A(regs_3[29]), .Z(n_31832));
	notech_inv i_31858(.A(regs_3[30]), .Z(n_31833));
	notech_inv i_31859(.A(regs_3[31]), .Z(n_31834));
	notech_inv i_31860(.A(gs[0]), .Z(n_31835));
	notech_inv i_31861(.A(gs[1]), .Z(n_31836));
	notech_inv i_31862(.A(n_56951), .Z(n_31837));
	notech_inv i_31863(.A(gs[3]), .Z(n_31838));
	notech_inv i_31864(.A(gs[4]), .Z(n_31839));
	notech_inv i_31865(.A(gs[5]), .Z(n_31840));
	notech_inv i_31866(.A(gs[6]), .Z(n_31841));
	notech_inv i_31867(.A(gs[7]), .Z(n_31842));
	notech_inv i_31868(.A(gs[8]), .Z(n_31843));
	notech_inv i_31869(.A(gs[9]), .Z(n_31844));
	notech_inv i_31870(.A(gs[10]), .Z(n_31845));
	notech_inv i_31871(.A(gs[11]), .Z(n_31846));
	notech_inv i_31872(.A(gs[12]), .Z(n_31847));
	notech_inv i_31873(.A(gs[13]), .Z(n_31848));
	notech_inv i_31874(.A(gs[14]), .Z(n_31849));
	notech_inv i_31875(.A(gs[15]), .Z(n_31850));
	notech_inv i_31876(.A(gs[16]), .Z(n_31851));
	notech_inv i_31877(.A(gs[17]), .Z(n_31852));
	notech_inv i_31878(.A(gs[18]), .Z(n_31853));
	notech_inv i_31879(.A(gs[19]), .Z(n_31854));
	notech_inv i_31880(.A(gs[20]), .Z(n_31855));
	notech_inv i_31881(.A(gs[21]), .Z(n_31856));
	notech_inv i_31882(.A(gs[22]), .Z(n_31857));
	notech_inv i_31883(.A(gs[23]), .Z(n_31858));
	notech_inv i_31884(.A(gs[24]), .Z(n_31859));
	notech_inv i_31885(.A(gs[25]), .Z(n_31860));
	notech_inv i_31886(.A(gs[26]), .Z(n_31861));
	notech_inv i_31887(.A(gs[27]), .Z(n_31862));
	notech_inv i_31892(.A(gs[28]), .Z(n_31863));
	notech_inv i_31893(.A(gs[29]), .Z(n_31864));
	notech_inv i_31896(.A(gs[30]), .Z(n_31865));
	notech_inv i_31897(.A(gs[31]), .Z(n_31866));
	notech_inv i_31899(.A(regs_5[0]), .Z(n_31867));
	notech_inv i_31902(.A(regs_5[1]), .Z(n_31868));
	notech_inv i_31903(.A(regs_5[2]), .Z(n_31869));
	notech_inv i_31904(.A(regs_5[3]), .Z(n_31870));
	notech_inv i_31905(.A(regs_5[4]), .Z(n_31871));
	notech_inv i_31906(.A(regs_5[5]), .Z(n_31872));
	notech_inv i_31907(.A(regs_5[6]), .Z(n_31873));
	notech_inv i_31908(.A(regs_5[7]), .Z(n_31874));
	notech_inv i_31909(.A(regs_5[8]), .Z(n_31875));
	notech_inv i_31910(.A(regs_5[9]), .Z(n_31876));
	notech_inv i_31911(.A(regs_5[10]), .Z(n_31877));
	notech_inv i_31912(.A(regs_5[11]), .Z(n_31878));
	notech_inv i_31913(.A(regs_5[12]), .Z(n_31879));
	notech_inv i_31914(.A(regs_5[13]), .Z(n_31880));
	notech_inv i_31915(.A(regs_5[14]), .Z(n_31881));
	notech_inv i_31916(.A(regs_5[15]), .Z(n_31882));
	notech_inv i_31917(.A(regs_5[16]), .Z(n_31883));
	notech_inv i_31918(.A(regs_5[17]), .Z(n_31884));
	notech_inv i_31919(.A(regs_5[18]), .Z(n_31885));
	notech_inv i_31920(.A(regs_5[19]), .Z(n_31886));
	notech_inv i_31921(.A(regs_5[20]), .Z(n_31887));
	notech_inv i_31922(.A(regs_5[21]), .Z(n_31888));
	notech_inv i_31923(.A(regs_5[22]), .Z(n_31889));
	notech_inv i_31924(.A(regs_5[23]), .Z(n_31890));
	notech_inv i_31925(.A(regs_5[24]), .Z(n_31891));
	notech_inv i_31926(.A(regs_5[25]), .Z(n_31892));
	notech_inv i_31927(.A(regs_5[26]), .Z(n_31893));
	notech_inv i_31928(.A(regs_5[27]), .Z(n_31894));
	notech_inv i_31929(.A(regs_5[28]), .Z(n_31895));
	notech_inv i_31930(.A(regs_5[29]), .Z(n_31896));
	notech_inv i_31931(.A(regs_5[30]), .Z(n_31897));
	notech_inv i_31932(.A(regs_5[31]), .Z(n_31898));
	notech_inv i_31933(.A(regs_7[0]), .Z(n_31899));
	notech_inv i_31934(.A(regs_7[1]), .Z(n_31900));
	notech_inv i_31935(.A(regs_7[2]), .Z(n_31901));
	notech_inv i_31936(.A(regs_7[3]), .Z(n_31902));
	notech_inv i_31937(.A(regs_7[4]), .Z(n_31903));
	notech_inv i_31938(.A(regs_7[5]), .Z(n_31904));
	notech_inv i_31939(.A(regs_7[6]), .Z(n_31905));
	notech_inv i_31940(.A(regs_7[7]), .Z(n_31906));
	notech_inv i_31941(.A(regs_7[8]), .Z(n_31907));
	notech_inv i_31942(.A(regs_7[9]), .Z(n_31908));
	notech_inv i_31943(.A(regs_7[10]), .Z(n_31909));
	notech_inv i_31944(.A(regs_7[11]), .Z(n_31910));
	notech_inv i_31945(.A(regs_7[12]), .Z(n_31911));
	notech_inv i_31946(.A(regs_7[13]), .Z(n_31912));
	notech_inv i_31947(.A(regs_7[14]), .Z(n_31913));
	notech_inv i_31948(.A(regs_7[15]), .Z(n_31914));
	notech_inv i_31949(.A(regs_7[16]), .Z(n_31915));
	notech_inv i_31950(.A(regs_7[17]), .Z(n_31916));
	notech_inv i_31951(.A(regs_7[18]), .Z(n_31917));
	notech_inv i_31952(.A(regs_7[19]), .Z(n_31918));
	notech_inv i_31953(.A(regs_7[20]), .Z(n_31919));
	notech_inv i_31954(.A(regs_7[21]), .Z(n_31920));
	notech_inv i_31955(.A(regs_7[22]), .Z(n_31921));
	notech_inv i_31956(.A(regs_7[23]), .Z(n_31922));
	notech_inv i_31957(.A(regs_7[24]), .Z(n_31923));
	notech_inv i_31958(.A(regs_7[25]), .Z(n_31924));
	notech_inv i_31959(.A(regs_7[26]), .Z(n_31925));
	notech_inv i_31960(.A(regs_7[27]), .Z(n_31926));
	notech_inv i_31961(.A(regs_7[28]), .Z(n_31927));
	notech_inv i_31962(.A(regs_7[29]), .Z(n_31928));
	notech_inv i_31963(.A(regs_7[30]), .Z(n_31929));
	notech_inv i_31964(.A(regs_7[31]), .Z(n_31930));
	notech_inv i_31965(.A(regs_4[0]), .Z(n_31931));
	notech_inv i_31966(.A(regs_4[1]), .Z(n_31932));
	notech_inv i_31967(.A(regs_4[2]), .Z(n_31933));
	notech_inv i_31968(.A(regs_4[3]), .Z(n_31934));
	notech_inv i_31969(.A(regs_4[4]), .Z(n_31935));
	notech_inv i_31970(.A(regs_4[5]), .Z(n_31936));
	notech_inv i_31971(.A(regs_4[6]), .Z(n_31937));
	notech_inv i_31972(.A(regs_4[7]), .Z(n_31938));
	notech_inv i_31973(.A(regs_4[8]), .Z(n_31939));
	notech_inv i_31974(.A(regs_4[9]), .Z(n_31940));
	notech_inv i_31975(.A(regs_4[10]), .Z(n_31941));
	notech_inv i_31976(.A(regs_4[11]), .Z(n_31943));
	notech_inv i_31977(.A(regs_4[12]), .Z(n_31944));
	notech_inv i_31978(.A(regs_4[13]), .Z(n_31945));
	notech_inv i_31979(.A(regs_4[14]), .Z(n_31946));
	notech_inv i_31980(.A(regs_4[15]), .Z(n_31947));
	notech_inv i_31981(.A(regs_4[16]), .Z(n_31948));
	notech_inv i_31982(.A(regs_4[17]), .Z(n_31949));
	notech_inv i_31983(.A(regs_4[18]), .Z(n_31950));
	notech_inv i_31984(.A(regs_4[19]), .Z(n_31951));
	notech_inv i_31985(.A(regs_4[20]), .Z(n_31952));
	notech_inv i_31986(.A(regs_4[21]), .Z(n_31953));
	notech_inv i_31987(.A(regs_4[22]), .Z(n_31954));
	notech_inv i_31988(.A(regs_4[23]), .Z(n_31955));
	notech_inv i_31989(.A(regs_4[24]), .Z(n_31956));
	notech_inv i_31990(.A(regs_4[25]), .Z(n_31957));
	notech_inv i_31991(.A(regs_4[26]), .Z(n_31958));
	notech_inv i_31992(.A(regs_4[27]), .Z(n_31959));
	notech_inv i_31993(.A(regs_4[28]), .Z(n_31960));
	notech_inv i_31994(.A(regs_4[29]), .Z(n_31961));
	notech_inv i_31995(.A(regs_4[30]), .Z(n_31962));
	notech_inv i_31996(.A(regs_4[31]), .Z(n_31963));
	notech_inv i_31997(.A(regs_0[0]), .Z(n_31964));
	notech_inv i_31998(.A(regs_0[1]), .Z(n_31965));
	notech_inv i_31999(.A(regs_0[2]), .Z(n_31966));
	notech_inv i_32000(.A(regs_0[3]), .Z(n_31967));
	notech_inv i_32001(.A(regs_0[4]), .Z(n_31968));
	notech_inv i_32002(.A(regs_0[5]), .Z(n_31969));
	notech_inv i_32003(.A(regs_0[6]), .Z(n_31970));
	notech_inv i_32004(.A(regs_0[7]), .Z(n_31971));
	notech_inv i_32005(.A(regs_0[8]), .Z(n_31972));
	notech_inv i_32006(.A(regs_0[9]), .Z(n_31973));
	notech_inv i_32007(.A(regs_0[10]), .Z(n_31974));
	notech_inv i_32008(.A(regs_0[11]), .Z(n_31975));
	notech_inv i_32009(.A(regs_0[12]), .Z(n_31976));
	notech_inv i_32010(.A(regs_0[13]), .Z(n_31977));
	notech_inv i_32011(.A(regs_0[14]), .Z(n_31978));
	notech_inv i_32012(.A(regs_0[15]), .Z(n_31979));
	notech_inv i_32013(.A(regs_0[16]), .Z(n_31980));
	notech_inv i_32014(.A(regs_0[17]), .Z(n_31981));
	notech_inv i_32015(.A(regs_0[18]), .Z(n_31982));
	notech_inv i_32016(.A(regs_0[19]), .Z(n_31983));
	notech_inv i_32017(.A(regs_0[20]), .Z(n_31984));
	notech_inv i_32018(.A(regs_0[21]), .Z(n_31985));
	notech_inv i_32019(.A(regs_0[22]), .Z(n_31986));
	notech_inv i_32020(.A(regs_0[23]), .Z(n_31987));
	notech_inv i_32021(.A(regs_0[24]), .Z(n_31988));
	notech_inv i_32022(.A(regs_0[25]), .Z(n_31989));
	notech_inv i_32023(.A(regs_0[26]), .Z(n_31990));
	notech_inv i_32024(.A(regs_0[27]), .Z(n_31991));
	notech_inv i_32025(.A(regs_0[28]), .Z(n_31992));
	notech_inv i_32026(.A(regs_0[29]), .Z(n_31993));
	notech_inv i_32028(.A(regs_0[30]), .Z(n_31994));
	notech_inv i_32029(.A(regs_0[31]), .Z(n_31995));
	notech_inv i_32030(.A(regs_2[0]), .Z(n_31996));
	notech_inv i_32031(.A(regs_2[1]), .Z(n_31997));
	notech_inv i_32032(.A(regs_2[2]), .Z(n_31998));
	notech_inv i_32033(.A(regs_2[3]), .Z(n_31999));
	notech_inv i_32034(.A(regs_2[4]), .Z(n_32000));
	notech_inv i_32035(.A(regs_2[5]), .Z(n_32001));
	notech_inv i_32036(.A(regs_2[6]), .Z(n_32002));
	notech_inv i_32037(.A(regs_2[7]), .Z(n_32003));
	notech_inv i_32038(.A(regs_2[8]), .Z(n_32004));
	notech_inv i_32039(.A(regs_2[9]), .Z(n_32005));
	notech_inv i_32040(.A(regs_2[10]), .Z(n_32006));
	notech_inv i_32041(.A(regs_2[11]), .Z(n_32007));
	notech_inv i_32042(.A(regs_2[12]), .Z(n_32008));
	notech_inv i_32043(.A(regs_2[13]), .Z(n_32009));
	notech_inv i_32044(.A(regs_2[14]), .Z(n_32010));
	notech_inv i_32045(.A(regs_2[15]), .Z(n_32011));
	notech_inv i_32046(.A(regs_2[16]), .Z(n_32012));
	notech_inv i_32047(.A(regs_2[17]), .Z(n_32013));
	notech_inv i_32048(.A(regs_2[18]), .Z(n_32014));
	notech_inv i_32049(.A(regs_2[19]), .Z(n_32015));
	notech_inv i_32050(.A(regs_2[20]), .Z(n_32016));
	notech_inv i_32051(.A(regs_2[21]), .Z(n_32017));
	notech_inv i_32052(.A(regs_2[22]), .Z(n_32018));
	notech_inv i_32053(.A(regs_2[23]), .Z(n_32019));
	notech_inv i_32054(.A(regs_2[24]), .Z(n_32020));
	notech_inv i_32055(.A(regs_2[25]), .Z(n_32021));
	notech_inv i_32056(.A(regs_2[26]), .Z(n_32022));
	notech_inv i_32057(.A(regs_2[27]), .Z(n_32023));
	notech_inv i_32058(.A(regs_2[28]), .Z(n_32024));
	notech_inv i_32059(.A(regs_2[29]), .Z(n_32025));
	notech_inv i_32060(.A(regs_2[30]), .Z(n_32026));
	notech_inv i_32061(.A(regs_2[31]), .Z(n_32027));
	notech_inv i_32062(.A(nbus_11291[0]), .Z(n_32028));
	notech_inv i_32063(.A(nbus_11291[1]), .Z(n_32029));
	notech_inv i_32064(.A(nbus_11291[2]), .Z(n_32030));
	notech_inv i_32065(.A(nbus_11291[3]), .Z(n_32031));
	notech_inv i_32066(.A(nbus_11291[4]), .Z(n_32032));
	notech_inv i_32067(.A(nbus_11291[5]), .Z(n_32033));
	notech_inv i_32068(.A(nbus_11291[6]), .Z(n_32034));
	notech_inv i_32069(.A(nbus_11291[7]), .Z(n_32035));
	notech_inv i_32070(.A(nbus_11291[8]), .Z(n_32036));
	notech_inv i_32071(.A(nbus_11291[9]), .Z(n_32037));
	notech_inv i_32072(.A(nbus_11291[10]), .Z(n_32038));
	notech_inv i_32073(.A(nbus_11291[11]), .Z(n_32039));
	notech_inv i_32074(.A(nbus_11291[12]), .Z(n_32040));
	notech_inv i_32075(.A(nbus_11291[13]), .Z(n_32041));
	notech_inv i_32076(.A(nbus_11291[14]), .Z(n_32042));
	notech_inv i_32077(.A(nbus_11291[15]), .Z(n_32043));
	notech_inv i_32078(.A(nbus_11291[16]), .Z(n_32044));
	notech_inv i_32079(.A(nbus_11291[17]), .Z(n_32045));
	notech_inv i_32080(.A(nbus_11291[18]), .Z(n_32046));
	notech_inv i_32081(.A(nbus_11291[19]), .Z(n_32047));
	notech_inv i_32082(.A(nbus_11291[20]), .Z(n_32048));
	notech_inv i_32083(.A(nbus_11291[21]), .Z(n_32049));
	notech_inv i_32084(.A(nbus_11291[22]), .Z(n_32050));
	notech_inv i_32085(.A(nbus_11291[23]), .Z(n_32051));
	notech_inv i_32086(.A(nbus_11291[24]), .Z(n_32052));
	notech_inv i_32087(.A(nbus_11291[25]), .Z(n_32053));
	notech_inv i_32088(.A(nbus_11291[26]), .Z(n_32054));
	notech_inv i_32089(.A(nbus_11291[27]), .Z(n_32055));
	notech_inv i_32090(.A(nbus_11291[28]), .Z(n_32056));
	notech_inv i_32091(.A(nbus_11291[29]), .Z(n_32057));
	notech_inv i_32092(.A(nbus_11291[30]), .Z(n_32058));
	notech_inv i_32093(.A(nbus_11291[31]), .Z(n_32059));
	notech_inv i_32094(.A(regs_4_2[1]), .Z(n_32060));
	notech_inv i_32095(.A(regs_4_2[2]), .Z(n_32061));
	notech_inv i_32096(.A(regs_4_2[3]), .Z(n_32062));
	notech_inv i_32097(.A(regs_4_2[4]), .Z(n_32063));
	notech_inv i_32098(.A(regs_4_2[5]), .Z(n_32064));
	notech_inv i_32099(.A(regs_4_2[6]), .Z(n_32065));
	notech_inv i_32100(.A(regs_4_2[7]), .Z(n_32066));
	notech_inv i_32101(.A(regs_4_2[8]), .Z(n_32067));
	notech_inv i_32102(.A(regs_4_2[9]), .Z(n_32068));
	notech_inv i_32103(.A(regs_4_2[10]), .Z(n_32069));
	notech_inv i_32104(.A(regs_4_2[11]), .Z(n_32070));
	notech_inv i_32105(.A(regs_4_2[12]), .Z(n_32071));
	notech_inv i_32106(.A(regs_4_2[13]), .Z(n_32072));
	notech_inv i_32107(.A(regs_4_2[14]), .Z(n_32073));
	notech_inv i_32108(.A(regs_4_2[15]), .Z(n_32074));
	notech_inv i_32109(.A(regs_4_2[16]), .Z(n_32075));
	notech_inv i_32110(.A(regs_4_2[17]), .Z(n_32076));
	notech_inv i_32111(.A(regs_4_2[18]), .Z(n_32077));
	notech_inv i_32112(.A(regs_4_2[19]), .Z(n_32078));
	notech_inv i_32113(.A(regs_4_2[20]), .Z(n_32079));
	notech_inv i_32114(.A(regs_4_2[21]), .Z(n_32080));
	notech_inv i_32115(.A(regs_4_2[22]), .Z(n_32081));
	notech_inv i_32116(.A(regs_4_2[23]), .Z(n_32082));
	notech_inv i_32117(.A(regs_4_2[24]), .Z(n_32083));
	notech_inv i_32118(.A(regs_4_2[25]), .Z(n_32084));
	notech_inv i_32119(.A(regs_4_2[26]), .Z(n_32085));
	notech_inv i_32120(.A(regs_4_2[27]), .Z(n_32086));
	notech_inv i_32121(.A(regs_4_2[28]), .Z(n_32087));
	notech_inv i_32122(.A(regs_4_2[29]), .Z(n_32088));
	notech_inv i_32123(.A(regs_4_2[30]), .Z(n_32089));
	notech_inv i_32124(.A(regs_4_2[31]), .Z(n_32090));
	notech_inv i_32125(.A(instrc[0]), .Z(n_32091));
	notech_inv i_32126(.A(instrc[1]), .Z(n_32092));
	notech_inv i_32127(.A(instrc[2]), .Z(n_32093));
	notech_inv i_32128(.A(instrc[3]), .Z(n_32094));
	notech_inv i_32129(.A(instrc[4]), .Z(n_32095));
	notech_inv i_32130(.A(instrc[5]), .Z(n_32096));
	notech_inv i_32131(.A(instrc[6]), .Z(n_32097));
	notech_inv i_32132(.A(instrc[7]), .Z(n_32098));
	notech_inv i_32133(.A(instrc[8]), .Z(n_32099));
	notech_inv i_32134(.A(instrc[9]), .Z(n_32100));
	notech_inv i_32135(.A(instrc[10]), .Z(n_32101));
	notech_inv i_32136(.A(instrc[11]), .Z(n_32102));
	notech_inv i_32137(.A(instrc[12]), .Z(n_32103));
	notech_inv i_32138(.A(instrc[13]), .Z(n_32104));
	notech_inv i_32139(.A(instrc[14]), .Z(n_32105));
	notech_inv i_32140(.A(instrc[15]), .Z(n_32106));
	notech_inv i_32141(.A(instrc[16]), .Z(n_32107));
	notech_inv i_32142(.A(instrc[17]), .Z(n_32108));
	notech_inv i_32143(.A(instrc[18]), .Z(n_32109));
	notech_inv i_32144(.A(instrc[19]), .Z(n_32110));
	notech_inv i_32145(.A(instrc[20]), .Z(n_32111));
	notech_inv i_32146(.A(instrc[21]), .Z(n_32112));
	notech_inv i_32147(.A(instrc[22]), .Z(n_32113));
	notech_inv i_32148(.A(instrc[23]), .Z(n_32114));
	notech_inv i_32149(.A(instrc[24]), .Z(n_32115));
	notech_inv i_32150(.A(instrc[25]), .Z(n_32116));
	notech_inv i_32151(.A(instrc[26]), .Z(n_32117));
	notech_inv i_32152(.A(instrc[27]), .Z(n_32118));
	notech_inv i_32153(.A(instrc[28]), .Z(n_32119));
	notech_inv i_32154(.A(instrc[29]), .Z(n_32120));
	notech_inv i_32155(.A(instrc[30]), .Z(n_32121));
	notech_inv i_32156(.A(instrc[31]), .Z(n_32122));
	notech_inv i_32157(.A(instrc[32]), .Z(n_32123));
	notech_inv i_32158(.A(instrc[33]), .Z(n_32124));
	notech_inv i_32159(.A(instrc[34]), .Z(n_32125));
	notech_inv i_32160(.A(instrc[35]), .Z(n_32126));
	notech_inv i_32161(.A(instrc[36]), .Z(n_32127));
	notech_inv i_32162(.A(instrc[37]), .Z(n_32128));
	notech_inv i_32163(.A(instrc[38]), .Z(n_32129));
	notech_inv i_32164(.A(instrc[39]), .Z(n_32130));
	notech_inv i_32165(.A(instrc[40]), .Z(n_32131));
	notech_inv i_32166(.A(instrc[41]), .Z(n_32132));
	notech_inv i_32167(.A(instrc[42]), .Z(n_32133));
	notech_inv i_32168(.A(instrc[43]), .Z(n_32134));
	notech_inv i_32169(.A(instrc[44]), .Z(n_32135));
	notech_inv i_32170(.A(instrc[45]), .Z(n_32136));
	notech_inv i_32171(.A(instrc[46]), .Z(n_32137));
	notech_inv i_32172(.A(instrc[47]), .Z(n_32138));
	notech_inv i_32173(.A(instrc[64]), .Z(n_32139));
	notech_inv i_32174(.A(instrc[65]), .Z(n_32140));
	notech_inv i_32175(.A(instrc[66]), .Z(n_32141));
	notech_inv i_32176(.A(instrc[67]), .Z(n_32142));
	notech_inv i_32177(.A(instrc[68]), .Z(n_32143));
	notech_inv i_32178(.A(instrc[69]), .Z(n_32144));
	notech_inv i_32179(.A(instrc[70]), .Z(n_32145));
	notech_inv i_32180(.A(instrc[71]), .Z(n_32146));
	notech_inv i_32181(.A(instrc[72]), .Z(n_32147));
	notech_inv i_32182(.A(instrc[73]), .Z(n_32148));
	notech_inv i_32183(.A(instrc[74]), .Z(n_32149));
	notech_inv i_32184(.A(instrc[75]), .Z(n_32150));
	notech_inv i_32185(.A(instrc[76]), .Z(n_32151));
	notech_inv i_32186(.A(instrc[77]), .Z(n_32152));
	notech_inv i_32187(.A(instrc[78]), .Z(n_32153));
	notech_inv i_32188(.A(instrc[79]), .Z(n_32154));
	notech_inv i_32189(.A(instrc[108]), .Z(n_32155));
	notech_inv i_32190(.A(instrc[109]), .Z(n_32156));
	notech_inv i_32191(.A(n_60431), .Z(n_32157));
	notech_inv i_32192(.A(instrc[115]), .Z(n_32158));
	notech_inv i_32193(.A(n_61786), .Z(n_32159));
	notech_inv i_32194(.A(n_61964), .Z(n_32160));
	notech_inv i_32195(.A(n_61944), .Z(n_32161));
	notech_inv i_32196(.A(resb_shiftbox[0]), .Z(n_32162));
	notech_inv i_32197(.A(resb_shiftbox[1]), .Z(n_32163));
	notech_inv i_32198(.A(resb_shiftbox[2]), .Z(n_32164));
	notech_inv i_32199(.A(resb_shiftbox[8]), .Z(n_32165));
	notech_inv i_32202(.A(resb_shiftbox[9]), .Z(n_32166));
	notech_inv i_32204(.A(resb_shiftbox[10]), .Z(n_32167));
	notech_inv i_32205(.A(resb_shiftbox[11]), .Z(n_32168));
	notech_inv i_32206(.A(resb_shiftbox[12]), .Z(n_32169));
	notech_inv i_32207(.A(resb_shiftbox[13]), .Z(n_32170));
	notech_inv i_32208(.A(resb_shiftbox[14]), .Z(n_32171));
	notech_inv i_32209(.A(resb_shiftbox[15]), .Z(n_32172));
	notech_inv i_32210(.A(resb_shiftbox[16]), .Z(n_32173));
	notech_inv i_32211(.A(resb_shiftbox[19]), .Z(n_32174));
	notech_inv i_32212(.A(resb_shiftbox[20]), .Z(n_32175));
	notech_inv i_32213(.A(resb_shiftbox[21]), .Z(n_32177));
	notech_inv i_32215(.A(resb_shiftbox[22]), .Z(n_32178));
	notech_inv i_32216(.A(resb_shiftbox[23]), .Z(n_32179));
	notech_inv i_32217(.A(resb_shiftbox[24]), .Z(n_32180));
	notech_inv i_32218(.A(resb_shiftbox[25]), .Z(n_32182));
	notech_inv i_32219(.A(resb_shiftbox[26]), .Z(n_32183));
	notech_inv i_32220(.A(resb_shiftbox[27]), .Z(n_32185));
	notech_inv i_32221(.A(resb_shiftbox[28]), .Z(n_32187));
	notech_inv i_32222(.A(resb_shiftbox[29]), .Z(n_32189));
	notech_inv i_32223(.A(resb_shiftbox[30]), .Z(n_32190));
	notech_inv i_32224(.A(resb_shiftbox[31]), .Z(n_32191));
	notech_inv i_32225(.A(resb_shift4box[0]), .Z(n_32197));
	notech_inv i_32226(.A(resb_shift4box[1]), .Z(n_32198));
	notech_inv i_32227(.A(resb_shift4box[2]), .Z(n_32200));
	notech_inv i_32228(.A(resb_shift4box[3]), .Z(n_32201));
	notech_inv i_32229(.A(resb_shift4box[4]), .Z(n_32202));
	notech_inv i_32230(.A(resb_shift4box[8]), .Z(n_32205));
	notech_inv i_32231(.A(resb_shift4box[9]), .Z(n_32206));
	notech_inv i_32232(.A(resb_shift4box[10]), .Z(n_32207));
	notech_inv i_32233(.A(resb_shift4box[11]), .Z(n_32209));
	notech_inv i_32234(.A(resb_shift4box[12]), .Z(n_32212));
	notech_inv i_32235(.A(resb_shift4box[13]), .Z(n_32213));
	notech_inv i_32236(.A(resb_shift4box[14]), .Z(n_32214));
	notech_inv i_32237(.A(resb_shift4box[15]), .Z(n_32218));
	notech_inv i_32238(.A(resb_shift4box[16]), .Z(n_32221));
	notech_inv i_32239(.A(resb_shift4box[17]), .Z(n_32222));
	notech_inv i_32240(.A(resb_shift4box[18]), .Z(n_32225));
	notech_inv i_32241(.A(resb_shift4box[19]), .Z(n_32226));
	notech_inv i_32242(.A(resb_shift4box[20]), .Z(n_32228));
	notech_inv i_32243(.A(resb_shift4box[21]), .Z(n_32229));
	notech_inv i_32244(.A(resb_shift4box[22]), .Z(n_32230));
	notech_inv i_32245(.A(resb_shift4box[23]), .Z(n_32231));
	notech_inv i_32246(.A(resb_shift4box[24]), .Z(n_32232));
	notech_inv i_32247(.A(resb_shift4box[25]), .Z(n_32233));
	notech_inv i_32248(.A(resb_shift4box[26]), .Z(n_32234));
	notech_inv i_32249(.A(resb_shift4box[27]), .Z(n_32236));
	notech_inv i_32250(.A(resb_shift4box[28]), .Z(n_32237));
	notech_inv i_32251(.A(resb_shift4box[29]), .Z(n_32238));
	notech_inv i_32252(.A(resb_shift4box[30]), .Z(n_32239));
	notech_inv i_32253(.A(resb_shift4box[31]), .Z(n_32240));
	notech_inv i_32254(.A(imm[42]), .Z(n_32242));
	notech_inv i_32255(.A(imm[10]), .Z(n_32245));
	notech_inv i_32256(.A(imm[47]), .Z(n_32246));
	notech_inv i_32257(.A(imm[44]), .Z(n_32248));
	notech_inv i_32258(.A(imm[43]), .Z(n_32251));
	notech_inv i_32259(.A(imm[11]), .Z(n_32253));
	notech_inv i_32260(.A(imm[12]), .Z(n_32255));
	notech_inv i_32261(.A(imm[31]), .Z(n_32256));
	notech_inv i_32262(.A(imm[45]), .Z(n_32257));
	notech_inv i_32263(.A(imm[35]), .Z(n_32258));
	notech_inv i_32264(.A(imm[3]), .Z(n_32260));
	notech_inv i_32265(.A(imm[13]), .Z(n_32262));
	notech_inv i_32266(.A(imm[29]), .Z(n_32264));
	notech_inv i_32267(.A(imm[7]), .Z(n_32265));
	notech_inv i_32268(.A(imm[0]), .Z(n_32267));
	notech_inv i_32269(.A(imm[1]), .Z(n_32270));
	notech_inv i_32270(.A(imm[2]), .Z(n_32271));
	notech_inv i_32271(.A(imm[5]), .Z(n_32274));
	notech_inv i_32272(.A(imm[6]), .Z(n_32276));
	notech_inv i_32273(.A(imm[14]), .Z(n_32277));
	notech_inv i_32274(.A(imm[41]), .Z(n_32279));
	notech_inv i_32275(.A(imm[9]), .Z(n_32280));
	notech_inv i_32276(.A(imm[46]), .Z(n_32281));
	notech_inv i_32277(.A(imm[16]), .Z(n_32282));
	notech_inv i_32278(.A(imm[17]), .Z(n_32283));
	notech_inv i_32279(.A(imm[18]), .Z(n_32284));
	notech_inv i_32280(.A(imm[19]), .Z(n_32285));
	notech_inv i_32281(.A(imm[20]), .Z(n_32286));
	notech_inv i_32282(.A(imm[21]), .Z(n_32287));
	notech_inv i_32283(.A(imm[22]), .Z(n_32289));
	notech_inv i_32284(.A(imm[23]), .Z(n_32291));
	notech_inv i_32285(.A(imm[24]), .Z(n_32293));
	notech_inv i_32286(.A(imm[25]), .Z(n_32294));
	notech_inv i_32287(.A(imm[26]), .Z(n_32295));
	notech_inv i_32288(.A(imm[27]), .Z(n_32296));
	notech_inv i_32289(.A(imm[28]), .Z(n_32297));
	notech_inv i_32290(.A(imm[30]), .Z(n_32298));
	notech_inv i_32291(.A(imm[4]), .Z(n_32300));
	notech_inv i_32292(.A(imm[36]), .Z(n_32301));
	notech_inv i_32293(.A(imm[37]), .Z(n_32303));
	notech_inv i_32294(.A(imm[38]), .Z(n_32306));
	notech_inv i_32295(.A(imm[39]), .Z(n_32307));
	notech_inv i_32296(.A(imm[40]), .Z(n_32309));
	notech_inv i_32297(.A(imm[8]), .Z(n_32312));
	notech_inv i_32298(.A(add_src[0]), .Z(n_32313));
	notech_inv i_32299(.A(add_src[1]), .Z(n_32316));
	notech_inv i_32300(.A(add_src[2]), .Z(n_32318));
	notech_inv i_32301(.A(add_src[3]), .Z(n_32320));
	notech_inv i_32302(.A(add_src[5]), .Z(n_32322));
	notech_inv i_32303(.A(add_src[6]), .Z(n_32324));
	notech_inv i_32305(.A(add_src[7]), .Z(n_32325));
	notech_inv i_32306(.A(add_src[15]), .Z(n_32326));
	notech_inv i_32307(.A(add_src[16]), .Z(n_32327));
	notech_inv i_32308(.A(add_src[17]), .Z(n_32328));
	notech_inv i_32309(.A(add_src[18]), .Z(n_32329));
	notech_inv i_32310(.A(add_src[19]), .Z(n_32330));
	notech_inv i_32311(.A(add_src[20]), .Z(n_32331));
	notech_inv i_32312(.A(add_src[21]), .Z(n_32332));
	notech_inv i_32313(.A(add_src[22]), .Z(n_32333));
	notech_inv i_32314(.A(add_src[23]), .Z(n_32336));
	notech_inv i_32315(.A(add_src[24]), .Z(n_32337));
	notech_inv i_32316(.A(add_src[25]), .Z(n_32338));
	notech_inv i_32317(.A(add_src[26]), .Z(n_32339));
	notech_inv i_32318(.A(add_src[27]), .Z(n_32340));
	notech_inv i_32319(.A(add_src[28]), .Z(n_32341));
	notech_inv i_32320(.A(add_src[29]), .Z(n_32343));
	notech_inv i_32321(.A(add_src[30]), .Z(n_32344));
	notech_inv i_32322(.A(add_src[31]), .Z(n_32345));
	notech_inv i_32323(.A(opa_0[2]), .Z(n_32346));
	notech_inv i_32324(.A(opa_0[7]), .Z(n_32347));
	notech_inv i_32325(.A(opa_0[8]), .Z(n_32348));
	notech_inv i_32326(.A(opa_0[9]), .Z(n_32349));
	notech_inv i_32327(.A(opa_0[10]), .Z(n_32350));
	notech_inv i_32328(.A(opa_0[11]), .Z(n_32351));
	notech_inv i_32329(.A(opa_0[12]), .Z(n_32352));
	notech_inv i_32330(.A(opa_0[13]), .Z(n_32354));
	notech_inv i_32331(.A(opa_0[14]), .Z(n_32355));
	notech_inv i_32332(.A(opa_0[15]), .Z(n_32356));
	notech_inv i_32333(.A(opa_0[16]), .Z(n_32357));
	notech_inv i_32334(.A(opa_0[17]), .Z(n_32358));
	notech_inv i_32335(.A(opa_0[18]), .Z(n_32359));
	notech_inv i_32336(.A(opa_0[19]), .Z(n_32360));
	notech_inv i_32337(.A(opa_0[20]), .Z(n_32362));
	notech_inv i_32338(.A(opa_0[21]), .Z(n_32363));
	notech_inv i_32339(.A(opa_0[22]), .Z(n_32364));
	notech_inv i_32340(.A(opa_0[23]), .Z(n_32365));
	notech_inv i_32341(.A(opa_0[24]), .Z(n_32366));
	notech_inv i_32342(.A(opa_0[25]), .Z(n_32367));
	notech_inv i_32343(.A(opa_0[26]), .Z(n_32369));
	notech_inv i_32344(.A(opa_0[27]), .Z(n_32370));
	notech_inv i_32345(.A(opa_0[29]), .Z(n_32371));
	notech_inv i_32346(.A(opa_0[30]), .Z(n_32373));
	notech_inv i_32347(.A(opa_0[31]), .Z(n_32374));
	notech_inv i_32348(.A(resa_shiftbox[0]), .Z(n_32376));
	notech_inv i_32349(.A(resa_shiftbox[1]), .Z(n_32377));
	notech_inv i_32350(.A(resa_shiftbox[2]), .Z(n_32378));
	notech_inv i_32351(.A(resa_shiftbox[3]), .Z(n_32380));
	notech_inv i_32352(.A(resa_shiftbox[4]), .Z(n_32381));
	notech_inv i_32353(.A(resa_shiftbox[6]), .Z(n_32382));
	notech_inv i_32354(.A(resa_shiftbox[7]), .Z(n_32384));
	notech_inv i_32355(.A(resa_shiftbox[8]), .Z(n_32385));
	notech_inv i_32356(.A(resa_shiftbox[9]), .Z(n_32387));
	notech_inv i_32357(.A(resa_shiftbox[10]), .Z(n_32389));
	notech_inv i_32358(.A(resa_shiftbox[11]), .Z(n_32392));
	notech_inv i_32359(.A(resa_shiftbox[12]), .Z(n_32395));
	notech_inv i_32360(.A(resa_shiftbox[13]), .Z(n_32398));
	notech_inv i_32361(.A(resa_shiftbox[14]), .Z(n_32399));
	notech_inv i_32362(.A(resa_shiftbox[15]), .Z(n_32403));
	notech_inv i_32363(.A(resa_shiftbox[16]), .Z(n_32405));
	notech_inv i_32364(.A(resa_shiftbox[17]), .Z(n_32406));
	notech_inv i_32365(.A(resa_shiftbox[18]), .Z(n_32408));
	notech_inv i_32366(.A(resa_shiftbox[19]), .Z(n_32409));
	notech_inv i_32367(.A(resa_shiftbox[20]), .Z(n_32410));
	notech_inv i_32368(.A(resa_shiftbox[21]), .Z(n_32411));
	notech_inv i_32369(.A(resa_shiftbox[22]), .Z(n_32412));
	notech_inv i_32370(.A(resa_shiftbox[23]), .Z(n_32413));
	notech_inv i_32371(.A(resa_shiftbox[24]), .Z(n_32414));
	notech_inv i_32372(.A(resa_shiftbox[25]), .Z(n_32415));
	notech_inv i_32373(.A(resa_shiftbox[26]), .Z(n_32416));
	notech_inv i_32374(.A(resa_shiftbox[27]), .Z(n_32417));
	notech_inv i_32375(.A(resa_shiftbox[28]), .Z(n_32418));
	notech_inv i_32376(.A(resa_shiftbox[29]), .Z(n_32419));
	notech_inv i_32377(.A(resa_shiftbox[30]), .Z(n_32420));
	notech_inv i_32378(.A(resa_shiftbox[31]), .Z(n_32421));
	notech_inv i_32379(.A(resa_arithbox[0]), .Z(n_32422));
	notech_inv i_32380(.A(resa_arithbox[1]), .Z(n_32423));
	notech_inv i_32381(.A(resa_arithbox[2]), .Z(n_32424));
	notech_inv i_32382(.A(resa_arithbox[3]), .Z(n_32425));
	notech_inv i_32383(.A(resa_arithbox[4]), .Z(n_32426));
	notech_inv i_32384(.A(resa_arithbox[6]), .Z(n_32427));
	notech_inv i_32385(.A(resa_arithbox[7]), .Z(n_32428));
	notech_inv i_32386(.A(resa_arithbox[8]), .Z(n_32429));
	notech_inv i_32387(.A(resa_arithbox[9]), .Z(n_32430));
	notech_inv i_32388(.A(resa_arithbox[10]), .Z(n_32431));
	notech_inv i_32389(.A(resa_arithbox[13]), .Z(n_32432));
	notech_inv i_32390(.A(resa_arithbox[14]), .Z(n_32433));
	notech_inv i_32391(.A(resa_arithbox[15]), .Z(n_32434));
	notech_inv i_32392(.A(resa_arithbox[16]), .Z(n_32435));
	notech_inv i_32393(.A(resa_arithbox[17]), .Z(n_32436));
	notech_inv i_32394(.A(resa_arithbox[18]), .Z(n_32437));
	notech_inv i_32395(.A(resa_arithbox[19]), .Z(n_32438));
	notech_inv i_32396(.A(resa_arithbox[20]), .Z(n_32439));
	notech_inv i_32397(.A(resa_arithbox[21]), .Z(n_32440));
	notech_inv i_32398(.A(resa_arithbox[22]), .Z(n_32441));
	notech_inv i_32399(.A(resa_arithbox[23]), .Z(n_32442));
	notech_inv i_32400(.A(resa_arithbox[24]), .Z(n_32443));
	notech_inv i_32401(.A(resa_arithbox[25]), .Z(n_32444));
	notech_inv i_32402(.A(resa_arithbox[26]), .Z(n_32445));
	notech_inv i_32403(.A(resa_arithbox[27]), .Z(n_32446));
	notech_inv i_32404(.A(resa_arithbox[28]), .Z(n_32447));
	notech_inv i_32405(.A(resa_arithbox[29]), .Z(n_32448));
	notech_inv i_32406(.A(resa_arithbox[30]), .Z(n_32449));
	notech_inv i_32407(.A(resa_arithbox[31]), .Z(n_32450));
	notech_inv i_32408(.A(n_61279), .Z(n_32451));
	notech_inv i_32409(.A(resa_shift4box[0]), .Z(n_32452));
	notech_inv i_32412(.A(resa_shift4box[1]), .Z(n_32453));
	notech_inv i_32413(.A(resa_shift4box[2]), .Z(n_32454));
	notech_inv i_32414(.A(resa_shift4box[3]), .Z(n_32455));
	notech_inv i_32415(.A(resa_shift4box[4]), .Z(n_32456));
	notech_inv i_32416(.A(resa_shift4box[6]), .Z(n_32457));
	notech_inv i_32417(.A(resa_shift4box[7]), .Z(n_32458));
	notech_inv i_32418(.A(resa_shift4box[8]), .Z(n_32459));
	notech_inv i_32419(.A(resa_shift4box[9]), .Z(n_32460));
	notech_inv i_32421(.A(resa_shift4box[10]), .Z(n_32461));
	notech_inv i_32422(.A(resa_shift4box[11]), .Z(n_32462));
	notech_inv i_32423(.A(resa_shift4box[12]), .Z(n_32463));
	notech_inv i_32424(.A(resa_shift4box[13]), .Z(n_32464));
	notech_inv i_32425(.A(resa_shift4box[14]), .Z(n_32465));
	notech_inv i_32426(.A(resa_shift4box[15]), .Z(n_32466));
	notech_inv i_32427(.A(resa_shift4box[16]), .Z(n_32467));
	notech_inv i_32428(.A(resa_shift4box[17]), .Z(n_32468));
	notech_inv i_32429(.A(resa_shift4box[18]), .Z(n_32469));
	notech_inv i_32430(.A(resa_shift4box[19]), .Z(n_32470));
	notech_inv i_32431(.A(resa_shift4box[20]), .Z(n_32471));
	notech_inv i_32432(.A(resa_shift4box[21]), .Z(n_32472));
	notech_inv i_32433(.A(resa_shift4box[22]), .Z(n_32473));
	notech_inv i_32434(.A(resa_shift4box[23]), .Z(n_32474));
	notech_inv i_32435(.A(resa_shift4box[24]), .Z(n_32475));
	notech_inv i_32436(.A(resa_shift4box[25]), .Z(n_32476));
	notech_inv i_32437(.A(resa_shift4box[26]), .Z(n_32478));
	notech_inv i_32438(.A(resa_shift4box[27]), .Z(n_32480));
	notech_inv i_32439(.A(resa_shift4box[28]), .Z(n_32482));
	notech_inv i_32440(.A(resa_shift4box[29]), .Z(n_32483));
	notech_inv i_32441(.A(resa_shift4box[30]), .Z(n_32488));
	notech_inv i_32442(.A(resa_shift4box[31]), .Z(n_32489));
	notech_inv i_32443(.A(readio_data[0]), .Z(n_32490));
	notech_inv i_32444(.A(readio_data[1]), .Z(n_32491));
	notech_inv i_32446(.A(readio_data[2]), .Z(n_32492));
	notech_inv i_32447(.A(readio_data[3]), .Z(n_32493));
	notech_inv i_32448(.A(readio_data[4]), .Z(n_32494));
	notech_inv i_32449(.A(readio_data[5]), .Z(n_32496));
	notech_inv i_32450(.A(readio_data[6]), .Z(n_32500));
	notech_inv i_32451(.A(readio_data[7]), .Z(n_32501));
	notech_inv i_32452(.A(readio_data[8]), .Z(n_32502));
	notech_inv i_32453(.A(readio_data[9]), .Z(n_32503));
	notech_inv i_32454(.A(readio_data[10]), .Z(n_32504));
	notech_inv i_32455(.A(readio_data[11]), .Z(n_32507));
	notech_inv i_32456(.A(readio_data[12]), .Z(n_32509));
	notech_inv i_32458(.A(readio_data[13]), .Z(n_32510));
	notech_inv i_32459(.A(readio_data[14]), .Z(n_32511));
	notech_inv i_32460(.A(readio_data[15]), .Z(n_32512));
	notech_inv i_32461(.A(readio_data[16]), .Z(n_32513));
	notech_inv i_32463(.A(readio_data[17]), .Z(n_32515));
	notech_inv i_32464(.A(readio_data[18]), .Z(n_32516));
	notech_inv i_32465(.A(readio_data[19]), .Z(n_32517));
	notech_inv i_32467(.A(readio_data[20]), .Z(n_32518));
	notech_inv i_32468(.A(readio_data[21]), .Z(n_32519));
	notech_inv i_32469(.A(readio_data[22]), .Z(n_32523));
	notech_inv i_32470(.A(readio_data[24]), .Z(n_32524));
	notech_inv i_32471(.A(readio_data[25]), .Z(n_32525));
	notech_inv i_32472(.A(readio_data[26]), .Z(n_32526));
	notech_inv i_32473(.A(readio_data[27]), .Z(n_32527));
	notech_inv i_32474(.A(readio_data[28]), .Z(n_32528));
	notech_inv i_32475(.A(tsc[0]), .Z(n_32529));
	notech_inv i_32476(.A(tsc[2]), .Z(n_32530));
	notech_inv i_32477(.A(tsc[3]), .Z(n_32531));
	notech_inv i_32478(.A(tsc[4]), .Z(n_32532));
	notech_inv i_32479(.A(tsc[5]), .Z(n_32533));
	notech_inv i_32480(.A(tsc[6]), .Z(n_32534));
	notech_inv i_32481(.A(tsc[7]), .Z(n_32535));
	notech_inv i_32482(.A(tsc[8]), .Z(n_32537));
	notech_inv i_32483(.A(tsc[9]), .Z(n_32538));
	notech_inv i_32484(.A(tsc[10]), .Z(n_32539));
	notech_inv i_32485(.A(tsc[11]), .Z(n_32540));
	notech_inv i_32486(.A(tsc[12]), .Z(n_32541));
	notech_inv i_32487(.A(tsc[13]), .Z(n_32542));
	notech_inv i_32488(.A(tsc[14]), .Z(n_32543));
	notech_inv i_32489(.A(tsc[15]), .Z(n_32545));
	notech_inv i_32490(.A(tsc[20]), .Z(n_32546));
	notech_inv i_32491(.A(tsc[21]), .Z(n_32549));
	notech_inv i_32492(.A(tsc[22]), .Z(n_32550));
	notech_inv i_32493(.A(tsc[23]), .Z(n_32551));
	notech_inv i_32494(.A(tsc[25]), .Z(n_32552));
	notech_inv i_32495(.A(tsc[33]), .Z(n_32553));
	notech_inv i_32496(.A(tsc[34]), .Z(n_32554));
	notech_inv i_32497(.A(tsc[35]), .Z(n_32555));
	notech_inv i_32498(.A(tsc[36]), .Z(n_32556));
	notech_inv i_32499(.A(tsc[37]), .Z(n_32557));
	notech_inv i_32500(.A(tsc[38]), .Z(n_32558));
	notech_inv i_32501(.A(tsc[39]), .Z(n_32559));
	notech_inv i_32502(.A(tsc[40]), .Z(n_32560));
	notech_inv i_32503(.A(tsc[41]), .Z(n_32561));
	notech_inv i_32504(.A(tsc[42]), .Z(n_32562));
	notech_inv i_32505(.A(tsc[43]), .Z(n_32563));
	notech_inv i_32506(.A(tsc[44]), .Z(n_32564));
	notech_inv i_32507(.A(tsc[45]), .Z(n_32565));
	notech_inv i_32508(.A(tsc[46]), .Z(n_32566));
	notech_inv i_32509(.A(tsc[47]), .Z(n_32567));
	notech_inv i_32510(.A(tsc[49]), .Z(n_32568));
	notech_inv i_32511(.A(tsc[51]), .Z(n_32569));
	notech_inv i_32512(.A(tsc[52]), .Z(n_32570));
	notech_inv i_32513(.A(tsc[55]), .Z(n_32571));
	notech_inv i_32514(.A(tsc[56]), .Z(n_32572));
	notech_inv i_32515(.A(tsc[57]), .Z(n_32577));
	notech_inv i_32516(.A(tsc[58]), .Z(n_32578));
	notech_inv i_32517(.A(tsc[60]), .Z(n_32579));
	notech_inv i_32518(.A(tsc[61]), .Z(n_32580));
	notech_inv i_32519(.A(tsc[62]), .Z(n_32581));
	notech_inv i_32520(.A(tsc[63]), .Z(n_32582));
	notech_inv i_32521(.A(mul64[0]), .Z(n_32584));
	notech_inv i_32522(.A(mul64[1]), .Z(n_32585));
	notech_inv i_32523(.A(mul64[3]), .Z(n_32587));
	notech_inv i_32524(.A(mul64[4]), .Z(n_32588));
	notech_inv i_32525(.A(mul64[6]), .Z(n_32591));
	notech_inv i_32526(.A(divr_1[0]), .Z(n_32592));
	notech_inv i_32527(.A(divr_1[1]), .Z(n_32593));
	notech_inv i_32528(.A(divr_1[2]), .Z(n_32594));
	notech_inv i_32529(.A(divr_1[3]), .Z(n_32595));
	notech_inv i_32530(.A(divr_1[4]), .Z(n_32596));
	notech_inv i_32531(.A(divr_1[5]), .Z(n_32597));
	notech_inv i_32532(.A(divr_1[6]), .Z(n_32598));
	notech_inv i_32533(.A(divr_1[7]), .Z(n_32599));
	notech_inv i_32534(.A(divr_1[8]), .Z(n_32600));
	notech_inv i_32535(.A(divr_1[9]), .Z(n_32601));
	notech_inv i_32536(.A(divr_1[10]), .Z(n_32602));
	notech_inv i_32537(.A(divr_1[11]), .Z(n_32603));
	notech_inv i_32538(.A(divr_1[12]), .Z(n_32604));
	notech_inv i_32539(.A(divr_1[13]), .Z(n_32605));
	notech_inv i_32540(.A(divr_1[14]), .Z(n_32606));
	notech_inv i_32541(.A(divr_1[15]), .Z(n_32607));
	notech_inv i_32542(.A(divr_1[16]), .Z(n_32608));
	notech_inv i_32543(.A(divr_1[17]), .Z(n_32609));
	notech_inv i_32544(.A(divr_1[18]), .Z(n_32610));
	notech_inv i_32545(.A(divr_1[19]), .Z(n_32611));
	notech_inv i_32546(.A(divr_1[20]), .Z(n_32612));
	notech_inv i_32547(.A(divr_1[21]), .Z(n_32613));
	notech_inv i_32548(.A(divr_1[22]), .Z(n_32615));
	notech_inv i_32549(.A(divr_1[23]), .Z(n_32616));
	notech_inv i_32550(.A(divr_1[24]), .Z(n_32617));
	notech_inv i_32551(.A(divr_1[25]), .Z(n_32619));
	notech_inv i_32552(.A(divr_1[26]), .Z(n_32620));
	notech_inv i_32553(.A(divr_1[27]), .Z(n_32621));
	notech_inv i_32554(.A(divr_1[28]), .Z(n_32622));
	notech_inv i_32555(.A(divr_1[29]), .Z(n_32623));
	notech_inv i_32556(.A(divr_1[30]), .Z(n_32624));
	notech_inv i_32557(.A(divr_1[31]), .Z(n_32625));
	notech_inv i_32558(.A(divr_1[32]), .Z(n_32626));
	notech_inv i_32559(.A(divr_1[33]), .Z(n_32630));
	notech_inv i_32560(.A(divr_1[34]), .Z(n_32631));
	notech_inv i_32561(.A(divr_1[35]), .Z(n_32632));
	notech_inv i_32562(.A(divr_1[36]), .Z(n_32634));
	notech_inv i_32563(.A(divr_1[37]), .Z(n_32635));
	notech_inv i_32564(.A(divr_1[38]), .Z(n_32636));
	notech_inv i_32565(.A(divr_1[39]), .Z(n_32637));
	notech_inv i_32566(.A(divr_1[40]), .Z(n_32638));
	notech_inv i_32567(.A(divr_1[41]), .Z(n_32639));
	notech_inv i_32568(.A(divr_1[42]), .Z(n_32640));
	notech_inv i_32569(.A(divr_1[43]), .Z(n_32641));
	notech_inv i_32570(.A(divr_1[46]), .Z(n_32642));
	notech_inv i_32571(.A(divr_1[53]), .Z(n_32643));
	notech_inv i_32572(.A(divr_1[62]), .Z(n_32644));
	notech_inv i_32573(.A(divr_1[63]), .Z(n_32645));
	notech_inv i_32574(.A(Daddrs_3[2]), .Z(n_32647));
	notech_inv i_32575(.A(Daddrs_3[3]), .Z(n_32648));
	notech_inv i_32576(.A(Daddrs_3[4]), .Z(n_32649));
	notech_inv i_32577(.A(Daddrs_3[5]), .Z(n_32651));
	notech_inv i_32578(.A(Daddrs_3[6]), .Z(n_32652));
	notech_inv i_32579(.A(Daddrs_3[7]), .Z(n_32653));
	notech_inv i_32580(.A(Daddrs_3[8]), .Z(n_32654));
	notech_inv i_32581(.A(Daddrs_3[9]), .Z(n_32655));
	notech_inv i_32582(.A(Daddrs_1[2]), .Z(n_32656));
	notech_inv i_32583(.A(Daddrs_1[3]), .Z(n_32657));
	notech_inv i_32584(.A(Daddrs_1[4]), .Z(n_32658));
	notech_inv i_32585(.A(Daddrs_1[5]), .Z(n_32659));
	notech_inv i_32586(.A(Daddrs_1[6]), .Z(n_32660));
	notech_inv i_32587(.A(Daddrs_1[7]), .Z(n_32661));
	notech_inv i_32588(.A(Daddrs_1[8]), .Z(n_32662));
	notech_inv i_32589(.A(Daddrs_1[9]), .Z(n_32664));
	notech_inv i_32590(.A(write_data_33[0]), .Z(n_32665));
	notech_inv i_32591(.A(write_data_33[1]), .Z(n_32666));
	notech_inv i_32592(.A(write_data_33[2]), .Z(n_32667));
	notech_inv i_32593(.A(write_data_33[3]), .Z(n_32668));
	notech_inv i_32594(.A(write_data_33[4]), .Z(n_32669));
	notech_inv i_32595(.A(write_data_33[5]), .Z(n_32670));
	notech_inv i_32596(.A(write_data_33[6]), .Z(n_32671));
	notech_inv i_32597(.A(write_data_33[7]), .Z(n_32672));
	notech_inv i_32598(.A(write_data_33[8]), .Z(n_32673));
	notech_inv i_32599(.A(write_data_33[9]), .Z(n_32674));
	notech_inv i_32600(.A(write_data_33[10]), .Z(n_32675));
	notech_inv i_32601(.A(write_data_33[11]), .Z(n_32676));
	notech_inv i_32602(.A(write_data_33[12]), .Z(n_32677));
	notech_inv i_32603(.A(write_data_33[13]), .Z(n_32678));
	notech_inv i_32604(.A(write_data_33[14]), .Z(n_32679));
	notech_inv i_32605(.A(write_data_33[15]), .Z(n_32680));
	notech_inv i_32606(.A(write_data_33[16]), .Z(n_32681));
	notech_inv i_32607(.A(write_data_33[17]), .Z(n_32682));
	notech_inv i_32608(.A(write_data_33[18]), .Z(n_32683));
	notech_inv i_32609(.A(write_data_33[19]), .Z(n_32685));
	notech_inv i_32610(.A(write_data_33[20]), .Z(n_32686));
	notech_inv i_32611(.A(write_data_33[21]), .Z(n_32687));
	notech_inv i_32612(.A(write_data_33[22]), .Z(n_32688));
	notech_inv i_32613(.A(write_data_33[23]), .Z(n_32690));
	notech_inv i_32614(.A(write_data_33[24]), .Z(n_32691));
	notech_inv i_32615(.A(write_data_33[25]), .Z(n_32692));
	notech_inv i_32616(.A(write_data_33[26]), .Z(n_32693));
	notech_inv i_32617(.A(write_data_33[27]), .Z(n_32694));
	notech_inv i_32618(.A(write_data_33[28]), .Z(n_32695));
	notech_inv i_32619(.A(write_data_33[29]), .Z(n_32696));
	notech_inv i_32620(.A(write_data_33[30]), .Z(n_32698));
	notech_inv i_32621(.A(write_data_33[31]), .Z(n_32699));
	notech_inv i_32622(.A(nbus_135[5]), .Z(n_32700));
	notech_inv i_32623(.A(nbus_135[7]), .Z(n_32701));
	notech_inv i_32624(.A(nbus_135[8]), .Z(n_32702));
	notech_inv i_32625(.A(nbus_136[0]), .Z(n_32703));
	notech_inv i_32626(.A(nbus_136[1]), .Z(n_32704));
	notech_inv i_32627(.A(nbus_136[2]), .Z(n_32705));
	notech_inv i_32628(.A(nbus_136[3]), .Z(n_32706));
	notech_inv i_32629(.A(nbus_136[4]), .Z(n_32707));
	notech_inv i_32630(.A(nbus_136[5]), .Z(n_32708));
	notech_inv i_32631(.A(nbus_136[6]), .Z(n_32709));
	notech_inv i_32632(.A(nbus_136[7]), .Z(n_32710));
	notech_inv i_32633(.A(nbus_136[8]), .Z(n_32711));
	notech_inv i_32634(.A(nbus_136[9]), .Z(n_32712));
	notech_inv i_32635(.A(nbus_136[10]), .Z(n_32713));
	notech_inv i_32636(.A(nbus_136[11]), .Z(n_32714));
	notech_inv i_32637(.A(nbus_136[12]), .Z(n_32715));
	notech_inv i_32638(.A(nbus_136[13]), .Z(n_32716));
	notech_inv i_32639(.A(nbus_136[14]), .Z(n_32717));
	notech_inv i_32640(.A(nbus_136[16]), .Z(n_32718));
	notech_inv i_32641(.A(nbus_136[17]), .Z(n_32719));
	notech_inv i_32642(.A(nbus_136[18]), .Z(n_32720));
	notech_inv i_32643(.A(nbus_136[19]), .Z(n_32722));
	notech_inv i_32644(.A(nbus_136[20]), .Z(n_32723));
	notech_inv i_32645(.A(nbus_136[21]), .Z(n_32724));
	notech_inv i_32646(.A(nbus_136[22]), .Z(n_32725));
	notech_inv i_32647(.A(nbus_136[23]), .Z(n_32726));
	notech_inv i_32648(.A(nbus_136[24]), .Z(n_32727));
	notech_inv i_32649(.A(nbus_136[25]), .Z(n_32728));
	notech_inv i_32650(.A(nbus_136[26]), .Z(n_32729));
	notech_inv i_32651(.A(nbus_136[27]), .Z(n_32730));
	notech_inv i_32652(.A(nbus_136[28]), .Z(n_32731));
	notech_inv i_32653(.A(nbus_136[29]), .Z(n_32732));
	notech_inv i_32654(.A(nbus_136[30]), .Z(n_32733));
	notech_inv i_32655(.A(nbus_136[31]), .Z(n_32734));
	notech_inv i_32656(.A(nbus_136[32]), .Z(n_32735));
	notech_inv i_32657(.A(nbus_140[0]), .Z(n_32736));
	notech_inv i_32658(.A(nbus_140[1]), .Z(n_32737));
	notech_inv i_32659(.A(nbus_140[2]), .Z(n_32738));
	notech_inv i_32660(.A(nbus_140[3]), .Z(n_32739));
	notech_inv i_32661(.A(nbus_140[4]), .Z(n_32740));
	notech_inv i_32662(.A(nbus_140[6]), .Z(n_32741));
	notech_inv i_32663(.A(nbus_140[7]), .Z(n_32742));
	notech_inv i_32664(.A(nbus_140[8]), .Z(n_32743));
	notech_inv i_32665(.A(nbus_140[9]), .Z(n_32744));
	notech_inv i_32666(.A(nbus_140[10]), .Z(n_32745));
	notech_inv i_32667(.A(nbus_140[11]), .Z(n_32746));
	notech_inv i_32668(.A(nbus_140[12]), .Z(n_32747));
	notech_inv i_32669(.A(nbus_140[13]), .Z(n_32748));
	notech_inv i_32670(.A(nbus_140[14]), .Z(n_32749));
	notech_inv i_32671(.A(nbus_140[15]), .Z(n_32750));
	notech_inv i_32672(.A(nbus_140[28]), .Z(n_32751));
	notech_inv i_32673(.A(nbus_140[32]), .Z(n_32752));
	notech_inv i_32674(.A(nbus_138[0]), .Z(n_32753));
	notech_inv i_32675(.A(nbus_138[1]), .Z(n_32754));
	notech_inv i_32676(.A(nbus_138[2]), .Z(n_32755));
	notech_inv i_32677(.A(nbus_138[3]), .Z(n_32757));
	notech_inv i_32678(.A(nbus_138[4]), .Z(n_32758));
	notech_inv i_32679(.A(nbus_138[6]), .Z(n_32759));
	notech_inv i_32680(.A(nbus_138[8]), .Z(n_32760));
	notech_inv i_32681(.A(nbus_138[9]), .Z(n_32761));
	notech_inv i_32682(.A(nbus_138[10]), .Z(n_32762));
	notech_inv i_32683(.A(nbus_138[11]), .Z(n_32763));
	notech_inv i_32684(.A(nbus_138[12]), .Z(n_32764));
	notech_inv i_32685(.A(nbus_138[13]), .Z(n_32765));
	notech_inv i_32686(.A(nbus_138[14]), .Z(n_32766));
	notech_inv i_32687(.A(nbus_138[15]), .Z(n_32767));
	notech_inv i_32688(.A(nbus_138[32]), .Z(n_32768));
	notech_inv i_32689(.A(nbus_133[0]), .Z(n_32769));
	notech_inv i_32690(.A(nbus_133[1]), .Z(n_32770));
	notech_inv i_32691(.A(nbus_133[2]), .Z(n_32771));
	notech_inv i_32692(.A(nbus_133[3]), .Z(n_32772));
	notech_inv i_32693(.A(nbus_133[4]), .Z(n_32773));
	notech_inv i_32694(.A(nbus_133[5]), .Z(n_32774));
	notech_inv i_32695(.A(nbus_133[6]), .Z(n_32775));
	notech_inv i_32696(.A(nbus_133[7]), .Z(n_32776));
	notech_inv i_32697(.A(nbus_133[8]), .Z(n_32777));
	notech_inv i_32698(.A(nbus_133[9]), .Z(n_32778));
	notech_inv i_32699(.A(nbus_133[10]), .Z(n_32780));
	notech_inv i_32700(.A(nbus_133[11]), .Z(n_32781));
	notech_inv i_32701(.A(nbus_133[12]), .Z(n_32782));
	notech_inv i_32702(.A(nbus_133[13]), .Z(n_32783));
	notech_inv i_32703(.A(nbus_133[14]), .Z(n_32784));
	notech_inv i_32704(.A(nbus_133[15]), .Z(n_32786));
	notech_inv i_32705(.A(nbus_133[16]), .Z(n_32787));
	notech_inv i_32706(.A(nbus_133[17]), .Z(n_32788));
	notech_inv i_32707(.A(nbus_133[18]), .Z(n_32790));
	notech_inv i_32708(.A(nbus_133[19]), .Z(n_32791));
	notech_inv i_32709(.A(nbus_133[20]), .Z(n_32792));
	notech_inv i_32710(.A(nbus_133[21]), .Z(n_32793));
	notech_inv i_32711(.A(nbus_133[22]), .Z(n_32794));
	notech_inv i_32712(.A(nbus_133[23]), .Z(n_32795));
	notech_inv i_32713(.A(nbus_133[24]), .Z(n_32796));
	notech_inv i_32714(.A(nbus_133[25]), .Z(n_32797));
	notech_inv i_32715(.A(nbus_133[26]), .Z(n_32798));
	notech_inv i_32716(.A(nbus_133[27]), .Z(n_32799));
	notech_inv i_32717(.A(nbus_133[28]), .Z(n_32800));
	notech_inv i_32718(.A(nbus_133[29]), .Z(n_32801));
	notech_inv i_32719(.A(nbus_133[30]), .Z(n_32802));
	notech_inv i_32720(.A(nbus_133[31]), .Z(n_32803));
	notech_inv i_32721(.A(nbus_141[0]), .Z(n_32804));
	notech_inv i_32722(.A(nbus_141[1]), .Z(n_32805));
	notech_inv i_3272398760(.A(nbus_141[2]), .Z(n_32806));
	notech_inv i_32724(.A(nbus_141[3]), .Z(n_32807));
	notech_inv i_32725(.A(nbus_141[4]), .Z(n_32808));
	notech_inv i_32726(.A(nbus_141[5]), .Z(n_32809));
	notech_inv i_32727(.A(nbus_141[6]), .Z(n_32810));
	notech_inv i_3272898759(.A(nbus_141[7]), .Z(n_32811));
	notech_inv i_32729(.A(nbus_141[8]), .Z(n_32812));
	notech_inv i_32730(.A(nbus_141[9]), .Z(n_32813));
	notech_inv i_32731(.A(nbus_141[10]), .Z(n_32814));
	notech_inv i_32732(.A(nbus_141[11]), .Z(n_32815));
	notech_inv i_3273398758(.A(nbus_141[12]), .Z(n_32816));
	notech_inv i_32734(.A(nbus_141[13]), .Z(n_32817));
	notech_inv i_32737(.A(nbus_141[14]), .Z(n_32818));
	notech_inv i_3273898757(.A(nbus_141[15]), .Z(n_32819));
	notech_inv i_32739(.A(nbus_141[16]), .Z(n_32820));
	notech_inv i_32740(.A(nbus_139[0]), .Z(n_32821));
	notech_inv i_32741(.A(nbus_139[1]), .Z(n_32822));
	notech_inv i_32742(.A(nbus_139[2]), .Z(n_32823));
	notech_inv i_3274398756(.A(nbus_139[3]), .Z(n_32824));
	notech_inv i_32744(.A(nbus_139[4]), .Z(n_32825));
	notech_inv i_32745(.A(nbus_139[5]), .Z(n_32826));
	notech_inv i_32746(.A(nbus_139[6]), .Z(n_32827));
	notech_inv i_32747(.A(nbus_139[7]), .Z(n_32828));
	notech_inv i_3274898755(.A(nbus_139[8]), .Z(n_32829));
	notech_inv i_32749(.A(nbus_139[9]), .Z(n_32830));
	notech_inv i_32750(.A(nbus_139[10]), .Z(n_32831));
	notech_inv i_32751(.A(nbus_139[11]), .Z(n_32832));
	notech_inv i_32752(.A(nbus_139[12]), .Z(n_32833));
	notech_inv i_32753(.A(nbus_139[13]), .Z(n_32834));
	notech_inv i_32754(.A(nbus_139[14]), .Z(n_32835));
	notech_inv i_32755(.A(nbus_139[15]), .Z(n_32836));
	notech_inv i_32756(.A(nbus_139[16]), .Z(n_32837));
	notech_inv i_32757(.A(nbus_134[0]), .Z(n_32838));
	notech_inv i_32758(.A(nbus_134[1]), .Z(n_32839));
	notech_inv i_32759(.A(nbus_134[2]), .Z(n_32840));
	notech_inv i_32760(.A(nbus_134[3]), .Z(n_32841));
	notech_inv i_32761(.A(nbus_134[4]), .Z(n_32842));
	notech_inv i_32762(.A(nbus_134[6]), .Z(n_32843));
	notech_inv i_32763(.A(nbus_134[7]), .Z(n_32844));
	notech_inv i_32764(.A(nbus_134[8]), .Z(n_32845));
	notech_inv i_32765(.A(nbus_134[9]), .Z(n_32846));
	notech_inv i_32766(.A(nbus_134[10]), .Z(n_32847));
	notech_inv i_32768(.A(nbus_134[11]), .Z(n_32848));
	notech_inv i_32769(.A(nbus_134[12]), .Z(n_32849));
	notech_inv i_32770(.A(nbus_134[13]), .Z(n_32850));
	notech_inv i_32772(.A(nbus_134[14]), .Z(n_32851));
	notech_inv i_32773(.A(nbus_134[15]), .Z(n_32852));
	notech_inv i_32774(.A(nbus_143[0]), .Z(n_32853));
	notech_inv i_32775(.A(nbus_143[1]), .Z(n_32854));
	notech_inv i_32776(.A(nbus_143[2]), .Z(n_32855));
	notech_inv i_32777(.A(nbus_143[3]), .Z(n_32856));
	notech_inv i_32778(.A(nbus_143[5]), .Z(n_32857));
	notech_inv i_32779(.A(nbus_143[6]), .Z(n_32858));
	notech_inv i_32780(.A(nbus_143[7]), .Z(n_32859));
	notech_inv i_32781(.A(nbus_143[8]), .Z(n_32860));
	notech_inv i_32782(.A(nbus_143[9]), .Z(n_32861));
	notech_inv i_32783(.A(nbus_143[10]), .Z(n_32862));
	notech_inv i_32784(.A(nbus_143[11]), .Z(n_32863));
	notech_inv i_32785(.A(nbus_143[12]), .Z(n_32864));
	notech_inv i_32786(.A(nbus_143[13]), .Z(n_32865));
	notech_inv i_32787(.A(nbus_143[14]), .Z(n_32866));
	notech_inv i_32788(.A(nbus_143[15]), .Z(n_32867));
	notech_inv i_32789(.A(nbus_137[3]), .Z(n_32868));
	notech_inv i_32790(.A(nbus_137[4]), .Z(n_32869));
	notech_inv i_32791(.A(nbus_137[5]), .Z(n_32870));
	notech_inv i_32792(.A(nbus_137[6]), .Z(n_32871));
	notech_inv i_32793(.A(nbus_137[7]), .Z(n_32872));
	notech_inv i_32794(.A(nbus_137[8]), .Z(n_32873));
	notech_inv i_32795(.A(nbus_137[9]), .Z(n_32874));
	notech_inv i_32796(.A(nbus_137[10]), .Z(n_32875));
	notech_inv i_32797(.A(nbus_137[11]), .Z(n_32876));
	notech_inv i_32799(.A(nbus_137[12]), .Z(n_32877));
	notech_inv i_32800(.A(nbus_137[13]), .Z(n_32878));
	notech_inv i_32801(.A(nbus_137[14]), .Z(n_32879));
	notech_inv i_32802(.A(nbus_137[15]), .Z(n_32880));
	notech_inv i_32803(.A(nbus_142[0]), .Z(n_32881));
	notech_inv i_32804(.A(nbus_142[1]), .Z(n_32882));
	notech_inv i_32805(.A(nbus_142[2]), .Z(n_32883));
	notech_inv i_32806(.A(nbus_142[3]), .Z(n_32884));
	notech_inv i_32807(.A(nbus_142[4]), .Z(n_32885));
	notech_inv i_32808(.A(nbus_142[5]), .Z(n_32886));
	notech_inv i_32809(.A(nbus_142[6]), .Z(n_32887));
	notech_inv i_32810(.A(nbus_142[7]), .Z(n_32888));
	notech_inv i_32811(.A(nbus_142[8]), .Z(n_32889));
	notech_inv i_32812(.A(nbus_142[9]), .Z(n_32890));
	notech_inv i_32813(.A(nbus_142[10]), .Z(n_32891));
	notech_inv i_32814(.A(nbus_142[11]), .Z(n_32892));
	notech_inv i_32815(.A(nbus_142[12]), .Z(n_32893));
	notech_inv i_32816(.A(nbus_142[13]), .Z(n_32894));
	notech_inv i_32817(.A(nbus_142[14]), .Z(n_32895));
	notech_inv i_32818(.A(nbus_142[15]), .Z(n_32896));
	notech_inv i_32819(.A(nbus_142[16]), .Z(n_32897));
	notech_inv i_32820(.A(nbus_142[17]), .Z(n_32898));
	notech_inv i_32821(.A(nbus_142[18]), .Z(n_32899));
	notech_inv i_32822(.A(nbus_142[19]), .Z(n_32900));
	notech_inv i_32823(.A(nbus_142[20]), .Z(n_32901));
	notech_inv i_32824(.A(nbus_142[21]), .Z(n_32902));
	notech_inv i_32825(.A(nbus_142[22]), .Z(n_32903));
	notech_inv i_32826(.A(nbus_142[23]), .Z(n_32904));
	notech_inv i_32827(.A(nbus_142[24]), .Z(n_32905));
	notech_inv i_32828(.A(nbus_142[25]), .Z(n_32906));
	notech_inv i_32829(.A(nbus_142[26]), .Z(n_32907));
	notech_inv i_32830(.A(nbus_142[27]), .Z(n_32908));
	notech_inv i_32831(.A(nbus_142[28]), .Z(n_32909));
	notech_inv i_32832(.A(nbus_142[29]), .Z(n_32910));
	notech_inv i_32833(.A(nbus_142[30]), .Z(n_32911));
	notech_inv i_32834(.A(nbus_142[31]), .Z(n_32912));
	notech_inv i_32835(.A(nbus_142[32]), .Z(n_32913));
	notech_inv i_32836(.A(opc_14[0]), .Z(n_32914));
	notech_inv i_32837(.A(opc_14[1]), .Z(n_32915));
	notech_inv i_32838(.A(opc_14[2]), .Z(n_32916));
	notech_inv i_32839(.A(opc_14[3]), .Z(n_32917));
	notech_inv i_32840(.A(opc_14[4]), .Z(n_32918));
	notech_inv i_32841(.A(opc_14[5]), .Z(n_32919));
	notech_inv i_32842(.A(opc_14[6]), .Z(n_32920));
	notech_inv i_32843(.A(opc_14[7]), .Z(n_32921));
	notech_inv i_32844(.A(opc_14[8]), .Z(n_32922));
	notech_inv i_32845(.A(opc_14[9]), .Z(n_32923));
	notech_inv i_32846(.A(opc_14[10]), .Z(n_32924));
	notech_inv i_32847(.A(opc_14[11]), .Z(n_32925));
	notech_inv i_32848(.A(opc_14[12]), .Z(n_32926));
	notech_inv i_32849(.A(opc_14[13]), .Z(n_32927));
	notech_inv i_32850(.A(opc_14[14]), .Z(n_32928));
	notech_inv i_32851(.A(opc_14[15]), .Z(n_32929));
	notech_inv i_32852(.A(opc_14[16]), .Z(n_32930));
	notech_inv i_32853(.A(opc_14[31]), .Z(n_32931));
	notech_inv i_32854(.A(from_acu[0]), .Z(n_32932));
	notech_inv i_32855(.A(from_acu[1]), .Z(n_32933));
	notech_inv i_32856(.A(from_acu[2]), .Z(n_32934));
	notech_inv i_32857(.A(from_acu[3]), .Z(n_32935));
	notech_inv i_32858(.A(from_acu[4]), .Z(n_32936));
	notech_inv i_32859(.A(from_acu[5]), .Z(n_32937));
	notech_inv i_32860(.A(from_acu[6]), .Z(n_32938));
	notech_inv i_32861(.A(from_acu[7]), .Z(n_32939));
	notech_inv i_32862(.A(divq[0]), .Z(n_32940));
	notech_inv i_32863(.A(divq[1]), .Z(n_32941));
	notech_inv i_32864(.A(divq[2]), .Z(n_32942));
	notech_inv i_32865(.A(divq[3]), .Z(n_32943));
	notech_inv i_32866(.A(divq[4]), .Z(n_32944));
	notech_inv i_32867(.A(divq[5]), .Z(n_32945));
	notech_inv i_32868(.A(divq[6]), .Z(n_32946));
	notech_inv i_32869(.A(divq[7]), .Z(n_32947));
	notech_inv i_32870(.A(divq[8]), .Z(n_32948));
	notech_inv i_32871(.A(divq[9]), .Z(n_32949));
	notech_inv i_32872(.A(divq[10]), .Z(n_32950));
	notech_inv i_32873(.A(divq[11]), .Z(n_32951));
	notech_inv i_32874(.A(divq[12]), .Z(n_32952));
	notech_inv i_32875(.A(divq[13]), .Z(n_32953));
	notech_inv i_32876(.A(divq[14]), .Z(n_32954));
	notech_inv i_32877(.A(divq[15]), .Z(n_32955));
	notech_inv i_32878(.A(divq[16]), .Z(n_32956));
	notech_inv i_32879(.A(divq[17]), .Z(n_32957));
	notech_inv i_32880(.A(divq[18]), .Z(n_32958));
	notech_inv i_32881(.A(divq[19]), .Z(n_32959));
	notech_inv i_32882(.A(divq[20]), .Z(n_32960));
	notech_inv i_32883(.A(divq[21]), .Z(n_32961));
	notech_inv i_32884(.A(divq[22]), .Z(n_32962));
	notech_inv i_32885(.A(divq[23]), .Z(n_32963));
	notech_inv i_32886(.A(divq[24]), .Z(n_32964));
	notech_inv i_32887(.A(divq[25]), .Z(n_32965));
	notech_inv i_32888(.A(divq[26]), .Z(n_32966));
	notech_inv i_32889(.A(divq[27]), .Z(n_32967));
	notech_inv i_32890(.A(divq[28]), .Z(n_32968));
	notech_inv i_32891(.A(divq[29]), .Z(n_32969));
	notech_inv i_32892(.A(divq[30]), .Z(n_32970));
	notech_inv i_32893(.A(divq[31]), .Z(n_32971));
	notech_inv i_32894(.A(divq[32]), .Z(n_32972));
	notech_inv i_32895(.A(divq[33]), .Z(n_32973));
	notech_inv i_32896(.A(divq[34]), .Z(n_32974));
	notech_inv i_32897(.A(divq[35]), .Z(n_32975));
	notech_inv i_32898(.A(divq[36]), .Z(n_32976));
	notech_inv i_32899(.A(divq[37]), .Z(n_32977));
	notech_inv i_32900(.A(divq[38]), .Z(n_32978));
	notech_inv i_32901(.A(divq[39]), .Z(n_32979));
	notech_inv i_32902(.A(divq[40]), .Z(n_32980));
	notech_inv i_32903(.A(divq[41]), .Z(n_32981));
	notech_inv i_32904(.A(divq[42]), .Z(n_32982));
	notech_inv i_32905(.A(divq[43]), .Z(n_32983));
	notech_inv i_32906(.A(divq[44]), .Z(n_32984));
	notech_inv i_32907(.A(divq[45]), .Z(n_32985));
	notech_inv i_32908(.A(divq[46]), .Z(n_32986));
	notech_inv i_32909(.A(divq[47]), .Z(n_32987));
	notech_inv i_32910(.A(divq[48]), .Z(n_32988));
	notech_inv i_32911(.A(divq[49]), .Z(n_32989));
	notech_inv i_32912(.A(divq[50]), .Z(n_32990));
	notech_inv i_32913(.A(divq[51]), .Z(n_32991));
	notech_inv i_32914(.A(divq[52]), .Z(n_32992));
	notech_inv i_32915(.A(divq[53]), .Z(n_32993));
	notech_inv i_32916(.A(divq[54]), .Z(n_32994));
	notech_inv i_32917(.A(divq[55]), .Z(n_32995));
	notech_inv i_32918(.A(divq[56]), .Z(n_32996));
	notech_inv i_32919(.A(divq[57]), .Z(n_32997));
	notech_inv i_32920(.A(divq[58]), .Z(n_32998));
	notech_inv i_32921(.A(divq[59]), .Z(n_32999));
	notech_inv i_32922(.A(divq[60]), .Z(n_33000));
	notech_inv i_32923(.A(divq[61]), .Z(n_33001));
	notech_inv i_32924(.A(divq[62]), .Z(n_33002));
	notech_inv i_32925(.A(divq[63]), .Z(n_33003));
	notech_inv i_32926(.A(to_acu101153[0]), .Z(to_acu[0]));
	notech_inv i_32927(.A(to_acu101153[1]), .Z(to_acu[1]));
	notech_inv i_32928(.A(to_acu101153[2]), .Z(to_acu[2]));
	notech_inv i_32929(.A(to_acu101153[3]), .Z(to_acu[3]));
	notech_inv i_32930(.A(to_acu101153[4]), .Z(to_acu[4]));
	notech_inv i_32931(.A(to_acu101153[5]), .Z(to_acu[5]));
	notech_inv i_32932(.A(to_acu101153[6]), .Z(to_acu[6]));
	notech_inv i_32933(.A(to_acu101153[7]), .Z(to_acu[7]));
	notech_inv i_32934(.A(to_acu101153[8]), .Z(to_acu[8]));
	notech_inv i_32935(.A(to_acu101153[9]), .Z(to_acu[9]));
	notech_inv i_32936(.A(to_acu101153[10]), .Z(to_acu[10]));
	notech_inv i_32937(.A(to_acu101153[11]), .Z(to_acu[11]));
	notech_inv i_32938(.A(to_acu101153[12]), .Z(to_acu[12]));
	notech_inv i_32939(.A(to_acu101153[13]), .Z(to_acu[13]));
	notech_inv i_32940(.A(to_acu101153[14]), .Z(to_acu[14]));
	notech_inv i_32941(.A(to_acu101153[15]), .Z(to_acu[15]));
	notech_inv i_32942(.A(to_acu101153[16]), .Z(to_acu[16]));
	notech_inv i_32943(.A(to_acu101153[17]), .Z(to_acu[17]));
	notech_inv i_32944(.A(to_acu101153[18]), .Z(to_acu[18]));
	notech_inv i_32945(.A(to_acu101153[19]), .Z(to_acu[19]));
	notech_inv i_32946(.A(to_acu101153[20]), .Z(to_acu[20]));
	notech_inv i_32947(.A(to_acu101153[21]), .Z(to_acu[21]));
	notech_inv i_32948(.A(to_acu101153[22]), .Z(to_acu[22]));
	notech_inv i_32949(.A(to_acu101153[23]), .Z(to_acu[23]));
	notech_inv i_32950(.A(to_acu101153[24]), .Z(to_acu[24]));
	notech_inv i_32951(.A(to_acu101153[25]), .Z(to_acu[25]));
	notech_inv i_32952(.A(to_acu101153[26]), .Z(to_acu[26]));
	notech_inv i_32953(.A(to_acu101153[27]), .Z(to_acu[27]));
	notech_inv i_32954(.A(to_acu101153[28]), .Z(to_acu[28]));
	notech_inv i_32955(.A(to_acu101153[29]), .Z(to_acu[29]));
	notech_inv i_32956(.A(to_acu101153[30]), .Z(to_acu[30]));
	notech_inv i_32957(.A(to_acu101153[31]), .Z(to_acu[31]));
	notech_inv i_32958(.A(to_acu101153[32]), .Z(to_acu[32]));
	notech_inv i_32959(.A(to_acu101153[33]), .Z(to_acu[33]));
	notech_inv i_32960(.A(to_acu101153[34]), .Z(to_acu[34]));
	notech_inv i_32961(.A(to_acu101153[35]), .Z(to_acu[35]));
	notech_inv i_32962(.A(to_acu101153[36]), .Z(to_acu[36]));
	notech_inv i_32963(.A(to_acu101153[37]), .Z(to_acu[37]));
	notech_inv i_32964(.A(to_acu101153[38]), .Z(to_acu[38]));
	notech_inv i_32965(.A(to_acu101153[39]), .Z(to_acu[39]));
	notech_inv i_32966(.A(to_acu101153[40]), .Z(to_acu[40]));
	notech_inv i_32967(.A(to_acu101153[41]), .Z(to_acu[41]));
	notech_inv i_32968(.A(to_acu101153[42]), .Z(to_acu[42]));
	notech_inv i_32969(.A(to_acu101153[43]), .Z(to_acu[43]));
	notech_inv i_32970(.A(to_acu101153[44]), .Z(to_acu[44]));
	notech_inv i_32971(.A(to_acu101153[45]), .Z(to_acu[45]));
	notech_inv i_32972(.A(to_acu101153[46]), .Z(to_acu[46]));
	notech_inv i_32973(.A(to_acu101153[47]), .Z(to_acu[47]));
	notech_inv i_32974(.A(to_acu101153[48]), .Z(to_acu[48]));
	notech_inv i_32975(.A(to_acu101153[49]), .Z(to_acu[49]));
	notech_inv i_32976(.A(to_acu101153[50]), .Z(to_acu[50]));
	notech_inv i_32977(.A(to_acu101153[51]), .Z(to_acu[51]));
	notech_inv i_32978(.A(to_acu101153[52]), .Z(to_acu[52]));
	notech_inv i_32979(.A(to_acu101153[53]), .Z(to_acu[53]));
	notech_inv i_32980(.A(to_acu101153[54]), .Z(to_acu[54]));
	notech_inv i_32981(.A(to_acu101153[55]), .Z(to_acu[55]));
	notech_inv i_32982(.A(to_acu101153[56]), .Z(to_acu[56]));
	notech_inv i_32983(.A(to_acu101153[57]), .Z(to_acu[57]));
	notech_inv i_32984(.A(to_acu101153[58]), .Z(to_acu[58]));
	notech_inv i_32985(.A(to_acu101153[59]), .Z(to_acu[59]));
	notech_inv i_32986(.A(to_acu101153[60]), .Z(to_acu[60]));
	notech_inv i_32987(.A(to_acu101153[61]), .Z(to_acu[61]));
	notech_inv i_32988(.A(to_acu101153[62]), .Z(to_acu[62]));
	notech_inv i_32989(.A(to_acu101153[63]), .Z(to_acu[63]));
	notech_inv i_32990(.A(divr[0]), .Z(nbus_11270[0]));
	notech_inv i_32991(.A(divr[1]), .Z(nbus_11270[1]));
	notech_inv i_32992(.A(divr[2]), .Z(nbus_11270[2]));
	notech_inv i_32993(.A(divr[3]), .Z(nbus_11270[3]));
	notech_inv i_32994(.A(divr[4]), .Z(nbus_11270[4]));
	notech_inv i_32995(.A(divr[5]), .Z(nbus_11270[5]));
	notech_inv i_32996(.A(divr[6]), .Z(nbus_11270[6]));
	notech_inv i_32997(.A(divr[7]), .Z(nbus_11270[7]));
	notech_inv i_32998(.A(divr[8]), .Z(nbus_11270[8]));
	notech_inv i_32999(.A(divr[9]), .Z(nbus_11270[9]));
	notech_inv i_33000(.A(divr[10]), .Z(nbus_11270[10]));
	notech_inv i_33003(.A(divr[11]), .Z(nbus_11270[11]));
	notech_inv i_33006(.A(divr[12]), .Z(nbus_11270[12]));
	notech_inv i_33007(.A(divr[13]), .Z(nbus_11270[13]));
	notech_inv i_33008(.A(divr[14]), .Z(nbus_11270[14]));
	notech_inv i_33009(.A(divr[15]), .Z(nbus_11270[15]));
	notech_inv i_33010(.A(divr[16]), .Z(nbus_11270[16]));
	notech_inv i_33011(.A(divr[17]), .Z(nbus_11270[17]));
	notech_inv i_33012(.A(divr[18]), .Z(nbus_11270[18]));
	notech_inv i_33013(.A(divr[19]), .Z(nbus_11270[19]));
	notech_inv i_33015(.A(divr[20]), .Z(nbus_11270[20]));
	notech_inv i_33016(.A(divr[21]), .Z(nbus_11270[21]));
	notech_inv i_33017(.A(divr[22]), .Z(nbus_11270[22]));
	notech_inv i_33018(.A(divr[23]), .Z(nbus_11270[23]));
	notech_inv i_33019(.A(divr[24]), .Z(nbus_11270[24]));
	notech_inv i_33020(.A(divr[25]), .Z(nbus_11270[25]));
	notech_inv i_33021(.A(divr[26]), .Z(nbus_11270[26]));
	notech_inv i_33022(.A(divr[27]), .Z(nbus_11270[27]));
	notech_inv i_33023(.A(divr[28]), .Z(nbus_11270[28]));
	notech_inv i_33024(.A(divr[29]), .Z(nbus_11270[29]));
	notech_inv i_33025(.A(divr[30]), .Z(nbus_11270[30]));
	notech_inv i_33026(.A(divr[31]), .Z(nbus_11270[31]));
	notech_inv i_33027(.A(\regs_1[5] ), .Z(n_33100));
	notech_inv i_33028(.A(n_3477), .Z(n_33101));
	notech_inv i_33029(.A(\regs_1[4] ), .Z(n_33102));
	notech_inv i_33030(.A(\opa_12[1] ), .Z(n_33103));
	notech_inv i_33031(.A(\opa_12[4] ), .Z(n_33104));
	notech_inv i_33032(.A(n_1753), .Z(n_33105));
	notech_inv i_33033(.A(n_1754), .Z(n_33106));
	notech_inv i_33034(.A(n_2687), .Z(n_33107));
	notech_inv i_33035(.A(\eflags[10] ), .Z(n_33108));
	notech_inv i_33036(.A(n_2688), .Z(n_33109));
	notech_inv i_33037(.A(n_2732), .Z(n_33110));
	notech_inv i_33038(.A(\nbus_14543[23] ), .Z(n_33111));
	notech_inv i_33039(.A(\eflags[23] ), .Z(n_33112));
	notech_inv i_33040(.A(\nbus_14543[24] ), .Z(n_33113));
	notech_inv i_33041(.A(\eflags[24] ), .Z(n_33114));
	notech_inv i_33042(.A(\nbus_14543[25] ), .Z(n_33115));
	notech_inv i_33043(.A(\eflags[25] ), .Z(n_33116));
	notech_inv i_33044(.A(n_2710), .Z(n_33117));
	notech_inv i_33045(.A(\opa_12[3] ), .Z(n_33118));
	notech_inv i_33046(.A(\eflags[3] ), .Z(n_33119));
	notech_inv i_33047(.A(\nbus_14543[3] ), .Z(n_33120));
	notech_inv i_33048(.A(\eflags[7] ), .Z(n_33121));
	notech_inv i_33049(.A(\nbus_14543[7] ), .Z(n_33122));
	notech_inv i_33050(.A(\eflags[6] ), .Z(n_33123));
	notech_inv i_33051(.A(\nbus_14543[6] ), .Z(n_33124));
	notech_inv i_33052(.A(\eflags[5] ), .Z(n_33125));
	notech_inv i_33053(.A(\nbus_14543[5] ), .Z(n_33126));
	notech_inv i_33054(.A(\eflags[4] ), .Z(n_33127));
	notech_inv i_33055(.A(\nbus_14543[4] ), .Z(n_33128));
	notech_inv i_33056(.A(\eflags[2] ), .Z(n_33129));
	notech_inv i_33057(.A(\nbus_14543[2] ), .Z(n_33130));
	notech_inv i_33058(.A(ie), .Z(n_33131));
	notech_inv i_33059(.A(\nbus_14543[9] ), .Z(n_33132));
	notech_inv i_33060(.A(\eflags[1] ), .Z(n_33133));
	notech_inv i_33061(.A(\eflags[0] ), .Z(n_33134));
	notech_inv i_33062(.A(\opa_12[5] ), .Z(n_33135));
	notech_inv i_33063(.A(\opa_1[5] ), .Z(n_33136));
	notech_inv i_33064(.A(n_6264), .Z(n_33137));
	notech_inv i_33065(.A(instrc[91]), .Z(n_33138));
	notech_inv i_33066(.A(instrc[99]), .Z(n_33139));
	notech_inv i_33067(.A(instrc[96]), .Z(n_33140));
	notech_inv i_33068(.A(instrc[95]), .Z(n_33141));
	notech_inv i_33069(.A(instrc[103]), .Z(n_33142));
	notech_inv i_33070(.A(instrc[100]), .Z(n_33143));
	notech_inv i_33071(.A(instrc[80]), .Z(n_33144));
	notech_inv i_33072(.A(instrc[83]), .Z(n_33145));
	notech_inv i_33073(.A(instrc[87]), .Z(n_33146));
	notech_inv i_33074(.A(instrc[85]), .Z(n_33147));
	notech_inv i_33075(.A(instrc[86]), .Z(n_33148));
	notech_inv i_33076(.A(instrc[84]), .Z(n_33149));
	notech_inv i_33077(.A(instrc[81]), .Z(n_33150));
	notech_inv i_33078(.A(instrc[82]), .Z(n_33151));
	notech_inv i_33079(.A(instrc[116]), .Z(n_33152));
	notech_inv i_33080(.A(instrc[127]), .Z(n_33153));
	notech_inv i_33081(.A(instrc[89]), .Z(n_33154));
	notech_inv i_33082(.A(instrc[93]), .Z(n_33155));
	notech_inv i_33083(.A(instrc[105]), .Z(n_33156));
	notech_inv i_33084(.A(instrc[107]), .Z(n_33157));
	notech_inv i_33085(.A(n_61864), .Z(n_33158));
	notech_inv i_33086(.A(instrc[97]), .Z(n_33159));
	notech_inv i_33087(.A(instrc[88]), .Z(n_33160));
	notech_inv i_33088(.A(instrc[101]), .Z(n_33161));
	notech_inv i_33089(.A(instrc[124]), .Z(n_33162));
	notech_inv i_33090(.A(instrc[92]), .Z(n_33163));
	notech_inv i_33091(.A(instrc[106]), .Z(n_33164));
	notech_inv i_33092(.A(\opa_12[7] ), .Z(n_33165));
	notech_inv i_33093(.A(\opa_12[6] ), .Z(n_33166));
	notech_inv i_33094(.A(\opa_12[2] ), .Z(n_33167));
	notech_inv i_33095(.A(\opa_12[9] ), .Z(n_33168));
	notech_inv i_33096(.A(\opa_12[0] ), .Z(n_33169));
	notech_inv i_33097(.A(\regs_13_14[23] ), .Z(n_33170));
	notech_inv i_33098(.A(\regs_13_14[24] ), .Z(n_33171));
	notech_inv i_33099(.A(\regs_13_14[25] ), .Z(n_33172));
	notech_inv i_33100(.A(n_57696), .Z(n_33173));
	notech_inv i_33101(.A(instrc[104]), .Z(n_33174));
	notech_inv i_33102(.A(instrc[126]), .Z(n_33175));
	notech_inv i_33103(.A(instrc[102]), .Z(n_33176));
	notech_inv i_33104(.A(instrc[94]), .Z(n_33177));
	notech_inv i_33105(.A(instrc[98]), .Z(n_33178));
	notech_inv i_33106(.A(instrc[90]), .Z(n_33179));
	notech_inv i_33107(.A(n_1734), .Z(n_33180));
	notech_inv i_33108(.A(n_1733), .Z(n_33181));
	notech_inv i_33109(.A(n_1728), .Z(n_33182));
	notech_inv i_33110(.A(n_1727), .Z(n_33183));
	notech_inv i_33111(.A(n_2665), .Z(n_33184));
	notech_inv i_33112(.A(n_2666), .Z(n_33185));
	notech_inv i_33113(.A(n_2659), .Z(n_33186));
	notech_inv i_33114(.A(n_2660), .Z(n_33187));
	notech_inv i_33115(.A(n_2717), .Z(n_33188));
	notech_inv i_33116(.A(\regs_1[13] ), .Z(n_33189));
	notech_inv i_33117(.A(n_3485), .Z(n_33190));
	notech_inv i_33118(.A(\regs_1[10] ), .Z(n_33191));
	notech_inv i_33119(.A(n_3482), .Z(n_33192));
	notech_inv i_33120(.A(\regs_1[7] ), .Z(n_33193));
	notech_inv i_33124(.A(\regs_13_14[30] ), .Z(n_33194));
	notech_inv i_33125(.A(\regs_13_14[27] ), .Z(n_33195));
	notech_inv i_33128(.A(\regs_13_14[28] ), .Z(n_33196));
	notech_inv i_33129(.A(\regs_13_14[29] ), .Z(n_33197));
	notech_inv i_33131(.A(\regs_13_14[26] ), .Z(n_33198));
	notech_inv i_33132(.A(\regs_13_14[16] ), .Z(n_33199));
	notech_inv i_33133(.A(\regs_13_14[17] ), .Z(n_33200));
	notech_inv i_33134(.A(\regs_13_14[18] ), .Z(n_33201));
	notech_inv i_33135(.A(\regs_13_14[19] ), .Z(n_33202));
	notech_inv i_33136(.A(n_6774), .Z(n_33203));
	notech_inv i_33137(.A(\opa_12[10] ), .Z(n_33204));
	notech_inv i_33138(.A(n_6771), .Z(n_33205));
	notech_inv i_33139(.A(\regs_13_14[31] ), .Z(n_33206));
	notech_inv i_33140(.A(\eflags[14] ), .Z(n_33207));
	notech_inv i_33141(.A(\nbus_14543[14] ), .Z(n_33208));
	notech_inv i_33142(.A(\nbus_14543[10] ), .Z(n_33209));
	notech_inv i_33143(.A(n_2720), .Z(n_33210));
	notech_inv i_33144(.A(\nbus_14543[13] ), .Z(n_33211));
	notech_inv i_33145(.A(\eflags[13] ), .Z(n_33212));
	notech_inv i_33146(.A(\opa_12[13] ), .Z(n_33213));
	notech_inv i_33147(.A(n_1568), .Z(n_33214));
	notech_inv i_33148(.A(\opa_12[14] ), .Z(n_33215));
	notech_inv i_33149(.A(n_1738), .Z(n_33216));
	notech_inv i_33150(.A(n_1737), .Z(n_33217));
	notech_inv i_33151(.A(n_1732), .Z(n_33218));
	notech_inv i_33152(.A(n_1731), .Z(n_33219));
	notech_inv i_33153(.A(n_1730), .Z(n_33220));
	notech_inv i_33154(.A(n_1729), .Z(n_33221));
	notech_inv i_33155(.A(n_1712), .Z(n_33222));
	notech_inv i_33156(.A(n_1711), .Z(n_33223));
	notech_inv i_33157(.A(n_2669), .Z(n_33224));
	notech_inv i_33158(.A(n_2670), .Z(n_33225));
	notech_inv i_33159(.A(n_2663), .Z(n_33226));
	notech_inv i_33160(.A(n_2664), .Z(n_33227));
	notech_inv i_33161(.A(n_2661), .Z(n_33228));
	notech_inv i_33162(.A(n_2662), .Z(n_33229));
	notech_inv i_33163(.A(n_2722), .Z(n_33230));
	notech_inv i_33164(.A(n_2719), .Z(n_33231));
	notech_inv i_33165(.A(n_2718), .Z(n_33232));
	notech_inv i_33166(.A(n_2709), .Z(n_33233));
	notech_inv i_33167(.A(\regs_1[12] ), .Z(n_33234));
	notech_inv i_33168(.A(n_3484), .Z(n_33235));
	notech_inv i_33169(.A(\regs_1[11] ), .Z(n_33236));
	notech_inv i_33170(.A(n_3483), .Z(n_33237));
	notech_inv i_33171(.A(\regs_1[2] ), .Z(n_33238));
	notech_inv i_33172(.A(n_3474), .Z(n_33239));
	notech_inv i_33173(.A(\regs_1[15] ), .Z(n_33240));
	notech_inv i_33174(.A(n_3487), .Z(n_33241));
	notech_inv i_33175(.A(read_ack), .Z(n_33242));
	notech_inv i_33176(.A(n_1757), .Z(n_33243));
	notech_inv i_33177(.A(n_1758), .Z(n_33244));
	notech_inv i_33178(.A(n_1755), .Z(n_33245));
	notech_inv i_33179(.A(n_1756), .Z(n_33246));
	notech_inv i_33180(.A(n_2731), .Z(n_33247));
	notech_inv i_33181(.A(\opa_12[15] ), .Z(n_33248));
	notech_inv i_33182(.A(n_6776), .Z(n_33249));
	notech_inv i_33183(.A(\opa_12[12] ), .Z(n_33250));
	notech_inv i_33184(.A(n_6773), .Z(n_33251));
	notech_inv i_33185(.A(n_6772), .Z(n_33252));
	notech_inv i_33186(.A(\opa_12[8] ), .Z(n_33253));
	notech_inv i_33187(.A(\nbus_14543[15] ), .Z(n_33254));
	notech_inv i_33188(.A(\eflags[15] ), .Z(n_33255));
	notech_inv i_33189(.A(\nbus_14543[12] ), .Z(n_33256));
	notech_inv i_33190(.A(\eflags[12] ), .Z(n_33257));
	notech_inv i_33191(.A(\opa_12[11] ), .Z(n_33258));
	notech_inv i_33192(.A(\nbus_14543[11] ), .Z(n_33259));
	notech_inv i_33193(.A(\eflags[11] ), .Z(n_33260));
	notech_inv i_33194(.A(n_2713), .Z(n_33261));
	notech_inv i_33195(.A(n_2652), .Z(n_33262));
	notech_inv i_33196(.A(n_2651), .Z(n_33263));
	notech_inv i_33197(.A(n_1720), .Z(n_33264));
	notech_inv i_33198(.A(n_1719), .Z(n_33265));
	notech_inv i_33199(.A(\regs_1[1] ), .Z(n_33266));
	notech_inv i_33200(.A(n_3473), .Z(n_33267));
	notech_inv i_33201(.A(\regs_1[6] ), .Z(n_33268));
	notech_inv i_33202(.A(n_3478), .Z(n_33269));
	notech_inv i_33203(.A(\regs_1[14] ), .Z(n_33270));
	notech_inv i_33204(.A(\regs_1_0[30] ), .Z(n_33271));
	notech_inv i_33205(.A(\regs_1_0[26] ), .Z(n_33272));
	notech_inv i_33206(.A(\regs_1_0[27] ), .Z(n_33273));
	notech_inv i_33207(.A(\regs_1_0[29] ), .Z(n_33274));
	notech_inv i_33208(.A(\nbus_14543[26] ), .Z(n_33275));
	notech_inv i_33209(.A(\eflags[26] ), .Z(n_33276));
	notech_inv i_33210(.A(\nbus_14543[27] ), .Z(n_33277));
	notech_inv i_33211(.A(\eflags[27] ), .Z(n_33278));
	notech_inv i_33212(.A(n_6786), .Z(n_33279));
	notech_inv i_33213(.A(n_6785), .Z(n_33280));
	notech_inv i_33214(.A(n_6784), .Z(n_33281));
	notech_inv i_33215(.A(\nbus_14543[22] ), .Z(n_33282));
	notech_inv i_33216(.A(\eflags[22] ), .Z(n_33283));
	notech_inv i_33217(.A(\regs_13_14[22] ), .Z(n_33284));
	notech_inv i_33218(.A(n_6783), .Z(n_33285));
	notech_inv i_33219(.A(\nbus_14543[21] ), .Z(n_33286));
	notech_inv i_33220(.A(\eflags[21] ), .Z(n_33287));
	notech_inv i_33221(.A(\regs_13_14[21] ), .Z(n_33288));
	notech_inv i_33222(.A(n_6782), .Z(n_33289));
	notech_inv i_33223(.A(\nbus_14543[20] ), .Z(n_33290));
	notech_inv i_33224(.A(\eflags[20] ), .Z(n_33291));
	notech_inv i_33225(.A(\regs_13_14[20] ), .Z(n_33292));
	notech_inv i_33226(.A(n_6781), .Z(n_33293));
	notech_inv i_33227(.A(\regs_1[3] ), .Z(n_33294));
	notech_inv i_33228(.A(n_3475), .Z(n_33295));
	notech_inv i_33229(.A(\regs_1_0[16] ), .Z(n_33296));
	notech_inv i_33230(.A(\regs_1_0[18] ), .Z(n_33297));
	notech_inv i_33231(.A(n_6767), .Z(n_33298));
	notech_inv i_33232(.A(\add_len_pc[6] ), .Z(n_33299));
	notech_inv i_33233(.A(n_6768), .Z(n_33300));
	notech_inv i_33234(.A(\add_len_pc[7] ), .Z(n_33301));
	notech_inv i_33235(.A(\nbus_14543[16] ), .Z(n_33302));
	notech_inv i_33236(.A(\eflags[16] ), .Z(n_33303));
	notech_inv i_33237(.A(\nbus_14543[17] ), .Z(n_33304));
	notech_inv i_33238(.A(\eflags[17] ), .Z(n_33305));
	notech_inv i_33239(.A(\nbus_14543[18] ), .Z(n_33306));
	notech_inv i_33240(.A(\eflags[18] ), .Z(n_33307));
	notech_inv i_33241(.A(\nbus_14543[19] ), .Z(n_33308));
	notech_inv i_33242(.A(\eflags[19] ), .Z(n_33309));
	notech_inv i_33243(.A(n_6761), .Z(n_33310));
	notech_inv i_33244(.A(n_6762), .Z(n_33311));
	notech_inv i_33245(.A(n_6769), .Z(n_33312));
	notech_inv i_33246(.A(\add_len_pc[8] ), .Z(n_33313));
	notech_inv i_33247(.A(\nbus_14543[8] ), .Z(n_33314));
	notech_inv i_33248(.A(\eflags[8] ), .Z(n_33315));
	notech_inv i_33249(.A(n_6775), .Z(n_33316));
	notech_inv i_33250(.A(\nbus_14543[31] ), .Z(n_33317));
	notech_inv i_33251(.A(\eflags[31] ), .Z(n_33318));
	notech_inv i_33252(.A(\eflags[30] ), .Z(n_33319));
	notech_inv i_33253(.A(\nbus_14543[30] ), .Z(n_33320));
	notech_inv i_33254(.A(start_up), .Z(n_33321));
	notech_inv i_33255(.A(\add_len_pc[30] ), .Z(n_33322));
	notech_inv i_33256(.A(n_6791), .Z(n_33323));
	notech_inv i_33257(.A(n_1445), .Z(n_33324));
	notech_inv i_33258(.A(n_1443), .Z(n_33325));
	notech_inv i_33259(.A(n_2711), .Z(n_33326));
	notech_inv i_33260(.A(n_2712), .Z(n_33327));
	notech_inv i_33261(.A(n_1751), .Z(n_33328));
	notech_inv i_33262(.A(n_1752), .Z(n_33329));
	notech_inv i_33263(.A(n_1749), .Z(n_33330));
	notech_inv i_33264(.A(n_1750), .Z(n_33331));
	notech_inv i_33266(.A(n_1747), .Z(n_33332));
	notech_inv i_33267(.A(n_1748), .Z(n_33333));
	notech_inv i_33268(.A(n_2689), .Z(n_33334));
	notech_inv i_33269(.A(n_2690), .Z(n_33335));
	notech_inv i_33270(.A(n_2685), .Z(n_33336));
	notech_inv i_33271(.A(n_2686), .Z(n_33337));
	notech_inv i_33272(.A(n_2683), .Z(n_33338));
	notech_inv i_33273(.A(n_2684), .Z(n_33339));
	notech_inv i_33274(.A(n_2681), .Z(n_33340));
	notech_inv i_33275(.A(n_2682), .Z(n_33341));
	notech_inv i_33276(.A(n_2679), .Z(n_33342));
	notech_inv i_33277(.A(n_2680), .Z(n_33343));
	notech_inv i_33278(.A(n_2730), .Z(n_33344));
	notech_inv i_33279(.A(n_2729), .Z(n_33345));
	notech_inv i_33280(.A(n_2728), .Z(n_33346));
	notech_inv i_33281(.A(n_2727), .Z(n_33347));
	notech_inv i_33282(.A(\opa_1[0] ), .Z(n_33348));
	notech_inv i_33283(.A(\opa_1[1] ), .Z(n_33349));
	notech_inv i_33284(.A(n_6260), .Z(n_33350));
	notech_inv i_33285(.A(\opa_1[3] ), .Z(n_33351));
	notech_inv i_33286(.A(n_6262), .Z(n_33352));
	notech_inv i_33287(.A(\opa_1[4] ), .Z(n_33353));
	notech_inv i_33288(.A(n_6263), .Z(n_33354));
	notech_inv i_33289(.A(\opa_1[6] ), .Z(n_33355));
	notech_inv i_33290(.A(n_6265), .Z(n_33356));
	notech_inv i_33291(.A(n_6266), .Z(n_33357));
	notech_inv i_33292(.A(\opa_1[7] ), .Z(n_33358));
	notech_inv i_33293(.A(\opa_1[8] ), .Z(n_33359));
	notech_inv i_33294(.A(mul64[8]), .Z(n_33360));
	notech_inv i_33295(.A(n_6267), .Z(n_33361));
	notech_inv i_33296(.A(\opa_1[9] ), .Z(n_33362));
	notech_inv i_33297(.A(mul64[9]), .Z(n_33363));
	notech_inv i_33298(.A(n_6268), .Z(n_33364));
	notech_inv i_33299(.A(\opa_1[10] ), .Z(n_33365));
	notech_inv i_33300(.A(mul64[10]), .Z(n_33366));
	notech_inv i_33301(.A(n_6269), .Z(n_33367));
	notech_inv i_33302(.A(\opa_1[11] ), .Z(n_33368));
	notech_inv i_33303(.A(mul64[11]), .Z(n_33369));
	notech_inv i_33304(.A(n_6270), .Z(n_33370));
	notech_inv i_33305(.A(\opa_1[12] ), .Z(n_33371));
	notech_inv i_33306(.A(mul64[12]), .Z(n_33372));
	notech_inv i_33307(.A(n_6271), .Z(n_33373));
	notech_inv i_33308(.A(\opa_1[13] ), .Z(n_33374));
	notech_inv i_33309(.A(mul64[13]), .Z(n_33375));
	notech_inv i_33310(.A(n_6272), .Z(n_33376));
	notech_inv i_33311(.A(\opa_1[14] ), .Z(n_33377));
	notech_inv i_33313(.A(mul64[14]), .Z(n_33378));
	notech_inv i_33314(.A(n_6273), .Z(n_33379));
	notech_inv i_33315(.A(\opa_1[15] ), .Z(n_33380));
	notech_inv i_33316(.A(mul64[15]), .Z(n_33381));
	notech_inv i_33317(.A(n_6274), .Z(n_33382));
	notech_inv i_33318(.A(n_6275), .Z(n_33383));
	notech_inv i_33319(.A(mul64[16]), .Z(n_33384));
	notech_inv i_33320(.A(n_6276), .Z(n_33385));
	notech_inv i_33321(.A(mul64[17]), .Z(n_33386));
	notech_inv i_33322(.A(n_6277), .Z(n_33387));
	notech_inv i_33323(.A(mul64[18]), .Z(n_33388));
	notech_inv i_33324(.A(n_6278), .Z(n_33389));
	notech_inv i_33325(.A(mul64[19]), .Z(n_33390));
	notech_inv i_33326(.A(n_6279), .Z(n_33391));
	notech_inv i_33327(.A(mul64[20]), .Z(n_33392));
	notech_inv i_33328(.A(n_6280), .Z(n_33393));
	notech_inv i_33329(.A(mul64[21]), .Z(n_33394));
	notech_inv i_33330(.A(n_6281), .Z(n_33395));
	notech_inv i_33331(.A(mul64[22]), .Z(n_33396));
	notech_inv i_33332(.A(n_6282), .Z(n_33397));
	notech_inv i_33333(.A(mul64[23]), .Z(n_33398));
	notech_inv i_33334(.A(n_6283), .Z(n_33399));
	notech_inv i_33335(.A(mul64[24]), .Z(n_33400));
	notech_inv i_33336(.A(n_6284), .Z(n_33401));
	notech_inv i_33337(.A(mul64[25]), .Z(n_33402));
	notech_inv i_33338(.A(n_6285), .Z(n_33403));
	notech_inv i_33341(.A(mul64[26]), .Z(n_33404));
	notech_inv i_33342(.A(n_6286), .Z(n_33405));
	notech_inv i_33343(.A(mul64[27]), .Z(n_33406));
	notech_inv i_33346(.A(n_6287), .Z(n_33407));
	notech_inv i_33347(.A(mul64[28]), .Z(n_33408));
	notech_inv i_33348(.A(n_6288), .Z(n_33409));
	notech_inv i_33349(.A(mul64[29]), .Z(n_33410));
	notech_inv i_33353(.A(n_6289), .Z(n_33411));
	notech_inv i_33354(.A(mul64[30]), .Z(n_33412));
	notech_inv i_33358(.A(n_6290), .Z(n_33413));
	notech_inv i_33359(.A(mul64[31]), .Z(n_33414));
	notech_inv i_33361(.A(n_2639), .Z(n_33415));
	notech_inv i_33362(.A(n_2641), .Z(n_33416));
	notech_inv i_33363(.A(n_2642), .Z(n_33417));
	notech_inv i_33364(.A(n_2644), .Z(n_33418));
	notech_inv i_33365(.A(n_2643), .Z(n_33419));
	notech_inv i_33366(.A(n_2648), .Z(n_33420));
	notech_inv i_33367(.A(n_2647), .Z(n_33421));
	notech_inv i_33368(.A(n_2650), .Z(n_33422));
	notech_inv i_33369(.A(n_2649), .Z(n_33423));
	notech_inv i_33370(.A(n_2654), .Z(n_33424));
	notech_inv i_33371(.A(n_2653), .Z(n_33425));
	notech_inv i_33372(.A(n_2657), .Z(n_33426));
	notech_inv i_33373(.A(n_2658), .Z(n_33427));
	notech_inv i_33374(.A(n_2699), .Z(n_33428));
	notech_inv i_33375(.A(n_2700), .Z(n_33429));
	notech_inv i_33376(.A(n_1716), .Z(n_33430));
	notech_inv i_33377(.A(n_1715), .Z(n_33431));
	notech_inv i_33378(.A(n_1718), .Z(n_33432));
	notech_inv i_33379(.A(n_1717), .Z(n_33433));
	notech_inv i_33380(.A(n_1722), .Z(n_33434));
	notech_inv i_33381(.A(n_1721), .Z(n_33435));
	notech_inv i_33382(.A(\regs_1[0] ), .Z(n_33436));
	notech_inv i_33383(.A(n_3472), .Z(n_33437));
	notech_inv i_33384(.A(n_2714), .Z(n_33438));
	notech_inv i_33385(.A(n_2668), .Z(n_33439));
	notech_inv i_33386(.A(n_2667), .Z(n_33440));
	notech_inv i_33387(.A(\regs_1_0[28] ), .Z(n_33441));
	notech_inv i_33388(.A(n_2692), .Z(n_33442));
	notech_inv i_33389(.A(n_2694), .Z(n_33443));
	notech_inv i_33390(.A(n_2696), .Z(n_33444));
	notech_inv i_33391(.A(n_2698), .Z(n_33445));
	notech_inv i_33392(.A(\regs_1_0[25] ), .Z(n_33446));
	notech_inv i_33393(.A(\regs_1_0[24] ), .Z(n_33447));
	notech_inv i_33394(.A(\regs_1_0[23] ), .Z(n_33448));
	notech_inv i_33395(.A(\regs_1_0[20] ), .Z(n_33449));
	notech_inv i_33396(.A(\regs_1_0[17] ), .Z(n_33450));
	notech_inv i_33397(.A(\regs_1_0[19] ), .Z(n_33451));
	notech_inv i_33398(.A(n_2646), .Z(n_33452));
	notech_inv i_33399(.A(n_2672), .Z(n_33453));
	notech_inv i_33400(.A(n_2674), .Z(n_33454));
	notech_inv i_33401(.A(n_2676), .Z(n_33455));
	notech_inv i_33402(.A(n_2678), .Z(n_33456));
	notech_inv i_33403(.A(n_6766), .Z(n_33457));
	notech_inv i_33404(.A(\add_len_pc[5] ), .Z(n_33458));
	notech_inv i_33405(.A(\regs_1_0[31] ), .Z(n_33459));
	notech_inv i_33406(.A(n_2656), .Z(n_33460));
	notech_inv i_33407(.A(n_2702), .Z(n_33461));
	notech_inv i_33408(.A(n_4727), .Z(n_33462));
	notech_inv i_33409(.A(n_4729), .Z(n_33463));
	notech_inv i_33410(.A(n_4730), .Z(n_33464));
	notech_inv i_33411(.A(n_1726), .Z(n_33465));
	notech_inv i_33412(.A(n_1725), .Z(n_33466));
	notech_inv i_33413(.A(n_2737), .Z(n_33467));
	notech_inv i_33414(.A(n_2716), .Z(n_33468));
	notech_inv i_33415(.A(\regs_1[9] ), .Z(n_33469));
	notech_inv i_33416(.A(n_3481), .Z(n_33470));
	notech_inv i_33417(.A(n_1766), .Z(n_33471));
	notech_inv i_33418(.A(n_2736), .Z(n_33472));
	notech_inv i_33419(.A(n_2735), .Z(n_33473));
	notech_inv i_33420(.A(n_2734), .Z(n_33474));
	notech_inv i_33421(.A(n_2733), .Z(n_33475));
	notech_inv i_33422(.A(n_6765), .Z(n_33476));
	notech_inv i_33423(.A(n_6764), .Z(n_33477));
	notech_inv i_33424(.A(n_6763), .Z(n_33478));
	notech_inv i_33425(.A(n_1714), .Z(n_33479));
	notech_inv i_33426(.A(n_2726), .Z(n_33480));
	notech_inv i_33427(.A(n_2725), .Z(n_33481));
	notech_inv i_33428(.A(n_2724), .Z(n_33482));
	notech_inv i_33429(.A(n_2723), .Z(n_33483));
	notech_inv i_33430(.A(n_6770), .Z(n_33484));
	notech_inv i_33431(.A(n_2738), .Z(n_33485));
	notech_inv i_33432(.A(\nbus_14543[28] ), .Z(n_33486));
	notech_inv i_33433(.A(\eflags[28] ), .Z(n_33487));
	notech_inv i_33434(.A(\nbus_14543[29] ), .Z(n_33488));
	notech_inv i_33435(.A(\eflags[29] ), .Z(n_33489));
	notech_inv i_33436(.A(n_3653), .Z(n_33490));
	notech_inv i_33437(.A(\opc_1[4] ), .Z(n_33491));
	notech_inv i_33438(.A(n_3686), .Z(n_33492));
	notech_inv i_33439(.A(mul64[36]), .Z(n_33493));
	notech_inv i_33440(.A(n_577), .Z(n_33494));
	notech_inv i_33441(.A(n_579), .Z(n_33495));
	notech_inv i_33442(.A(n_62397), .Z(n_33496));
	notech_inv i_33443(.A(n_4642), .Z(n_33497));
	notech_inv i_33444(.A(n_4643), .Z(n_33498));
	notech_inv i_33445(.A(n_4644), .Z(n_33499));
	notech_inv i_33446(.A(n_4637), .Z(n_33500));
	notech_inv i_33447(.A(n_4638), .Z(n_33501));
	notech_inv i_33448(.A(n_4639), .Z(n_33502));
	notech_inv i_33449(.A(n_4632), .Z(n_33503));
	notech_inv i_33450(.A(n_4633), .Z(n_33504));
	notech_inv i_33451(.A(n_4634), .Z(n_33505));
	notech_inv i_33452(.A(n_4627), .Z(n_33506));
	notech_inv i_33453(.A(n_4628), .Z(n_33507));
	notech_inv i_33454(.A(n_4629), .Z(n_33508));
	notech_inv i_33455(.A(n_4607), .Z(n_33509));
	notech_inv i_33456(.A(n_4608), .Z(n_33510));
	notech_inv i_33457(.A(n_4609), .Z(n_33511));
	notech_inv i_33458(.A(n_4602), .Z(n_33512));
	notech_inv i_33459(.A(n_4603), .Z(n_33513));
	notech_inv i_33460(.A(n_4604), .Z(n_33514));
	notech_inv i_33461(.A(n_4597), .Z(n_33515));
	notech_inv i_33462(.A(n_4598), .Z(n_33516));
	notech_inv i_33463(.A(n_4599), .Z(n_33517));
	notech_inv i_33464(.A(n_350885916), .Z(n_33518));
	notech_inv i_33465(.A(n_4587), .Z(n_33519));
	notech_inv i_33466(.A(n_4588), .Z(n_33520));
	notech_inv i_33467(.A(n_4589), .Z(n_33521));
	notech_inv i_33468(.A(n_350785915101152), .Z(n_350785915));
	notech_inv i_33469(.A(n_4582), .Z(n_33523));
	notech_inv i_33470(.A(n_4583), .Z(n_33524));
	notech_inv i_33471(.A(n_4584), .Z(n_33525));
	notech_inv i_33472(.A(n_350685914101151), .Z(n_350685914));
	notech_inv i_33473(.A(n_4577), .Z(n_33527));
	notech_inv i_33474(.A(n_4578), .Z(n_33528));
	notech_inv i_33475(.A(n_4579), .Z(n_33529));
	notech_inv i_33476(.A(n_350585913101150), .Z(n_350585913));
	notech_inv i_33477(.A(n_4572), .Z(n_33531));
	notech_inv i_33478(.A(n_4573), .Z(n_33532));
	notech_inv i_33479(.A(n_4574), .Z(n_33533));
	notech_inv i_33480(.A(n_2708), .Z(n_33534));
	notech_inv i_33485(.A(n_2721), .Z(n_33535));
	notech_inv i_33486(.A(n_1709), .Z(n_33536));
	notech_inv i_33487(.A(n_1710), .Z(n_33537));
	notech_inv i_33488(.A(n_1735), .Z(n_33538));
	notech_inv i_33489(.A(n_1768), .Z(n_33539));
	notech_inv i_33490(.A(n_1707), .Z(n_33540));
	notech_inv i_33491(.A(n_1760), .Z(n_33541));
	notech_inv i_33492(.A(n_1762), .Z(n_33542));
	notech_inv i_33493(.A(n_1764), .Z(n_33543));
	notech_inv i_33494(.A(n_1740), .Z(n_33544));
	notech_inv i_33495(.A(n_1742), .Z(n_33545));
	notech_inv i_33496(.A(n_1744), .Z(n_33546));
	notech_inv i_33497(.A(n_1746), .Z(n_33547));
	notech_inv i_33498(.A(\regs_1[8] ), .Z(n_33548));
	notech_inv i_33499(.A(n_2715), .Z(n_33549));
	notech_inv i_33500(.A(n_1724), .Z(n_33550));
	notech_inv i_33501(.A(n_1770), .Z(n_33551));
	notech_inv i_33503(.A(n_4593), .Z(n_33552));
	notech_inv i_33504(.A(\nbus_11309[4] ), .Z(n_33553));
	notech_inv i_33505(.A(n_3538), .Z(n_33554));
	notech_inv i_33506(.A(n_4707), .Z(n_33555));
	notech_inv i_33507(.A(n_4708), .Z(n_33556));
	notech_inv i_33508(.A(n_4709), .Z(n_33557));
	notech_inv i_33509(.A(n_4697), .Z(n_33558));
	notech_inv i_33510(.A(n_4698), .Z(n_33559));
	notech_inv i_33511(.A(n_4699), .Z(n_33560));
	notech_inv i_33512(.A(n_4677), .Z(n_33561));
	notech_inv i_33513(.A(n_4678), .Z(n_33562));
	notech_inv i_33514(.A(n_4679), .Z(n_33563));
	notech_inv i_33515(.A(n_4672), .Z(n_33564));
	notech_inv i_33516(.A(n_4673), .Z(n_33565));
	notech_inv i_33517(.A(n_4674), .Z(n_33566));
	notech_inv i_33518(.A(n_4667), .Z(n_33567));
	notech_inv i_33519(.A(n_4668), .Z(n_33568));
	notech_inv i_33520(.A(n_4669), .Z(n_33569));
	notech_inv i_33521(.A(n_4662), .Z(n_33570));
	notech_inv i_33522(.A(n_4663), .Z(n_33571));
	notech_inv i_33523(.A(n_4664), .Z(n_33572));
	notech_inv i_33524(.A(n_4657), .Z(n_33573));
	notech_inv i_33525(.A(n_4658), .Z(n_33574));
	notech_inv i_33526(.A(n_4659), .Z(n_33575));
	notech_inv i_33527(.A(n_4652), .Z(n_33576));
	notech_inv i_33528(.A(n_4653), .Z(n_33577));
	notech_inv i_33529(.A(n_4654), .Z(n_33578));
	notech_inv i_33530(.A(n_4712), .Z(n_33579));
	notech_inv i_33531(.A(n_4713), .Z(n_33580));
	notech_inv i_33532(.A(n_4714), .Z(n_33581));
	notech_inv i_33533(.A(n_4702), .Z(n_33582));
	notech_inv i_33534(.A(n_4703), .Z(n_33583));
	notech_inv i_33535(.A(n_4704), .Z(n_33584));
	notech_inv i_33536(.A(n_4692), .Z(n_33585));
	notech_inv i_33537(.A(n_4693), .Z(n_33586));
	notech_inv i_33538(.A(n_4694), .Z(n_33587));
	notech_inv i_33539(.A(n_4687), .Z(n_33588));
	notech_inv i_33540(.A(n_4688), .Z(n_33589));
	notech_inv i_33541(.A(n_4689), .Z(n_33590));
	notech_inv i_33542(.A(n_4682), .Z(n_33591));
	notech_inv i_33543(.A(n_4683), .Z(n_33592));
	notech_inv i_33544(.A(n_4684), .Z(n_33593));
	notech_inv i_33545(.A(n_6614), .Z(n_33594));
	notech_inv i_33546(.A(n_5280), .Z(n_33595));
	notech_inv i_33547(.A(n_6613), .Z(n_33596));
	notech_inv i_33548(.A(n_6618), .Z(n_33597));
	notech_inv i_33549(.A(n_6617), .Z(n_33598));
	notech_inv i_33550(.A(n_5282), .Z(n_33599));
	notech_inv i_33551(.A(n_6620), .Z(n_33600));
	notech_inv i_33552(.A(n_6619), .Z(n_33601));
	notech_inv i_33553(.A(n_5283), .Z(n_33602));
	notech_inv i_33554(.A(n_6622), .Z(n_33603));
	notech_inv i_33555(.A(n_6621), .Z(n_33604));
	notech_inv i_33556(.A(n_5284), .Z(n_33605));
	notech_inv i_33557(.A(n_6624), .Z(n_33606));
	notech_inv i_33558(.A(n_6623), .Z(n_33607));
	notech_inv i_33559(.A(n_5285), .Z(n_33608));
	notech_inv i_33560(.A(n_6626), .Z(n_33609));
	notech_inv i_33561(.A(n_6625), .Z(n_33610));
	notech_inv i_33562(.A(n_5286), .Z(n_33611));
	notech_inv i_33563(.A(n_6628), .Z(n_33612));
	notech_inv i_33564(.A(n_6627), .Z(n_33613));
	notech_inv i_33565(.A(n_5287), .Z(n_33614));
	notech_inv i_33566(.A(n_6630), .Z(n_33615));
	notech_inv i_33567(.A(n_6629), .Z(n_33616));
	notech_inv i_33568(.A(n_5288), .Z(n_33617));
	notech_inv i_33571(.A(n_6632), .Z(n_33618));
	notech_inv i_33572(.A(n_6631), .Z(n_33619));
	notech_inv i_33573(.A(n_5289), .Z(n_33620));
	notech_inv i_33574(.A(n_6634), .Z(n_33621));
	notech_inv i_33575(.A(n_5290), .Z(n_33622));
	notech_inv i_33576(.A(n_6633), .Z(n_33623));
	notech_inv i_33577(.A(n_6636), .Z(n_33624));
	notech_inv i_33578(.A(n_5291), .Z(n_33625));
	notech_inv i_33579(.A(n_6635), .Z(n_33626));
	notech_inv i_33580(.A(n_6638), .Z(n_33627));
	notech_inv i_33581(.A(n_5292), .Z(n_33628));
	notech_inv i_33582(.A(n_6637), .Z(n_33629));
	notech_inv i_33583(.A(n_6640), .Z(n_33630));
	notech_inv i_33584(.A(n_5293), .Z(n_33631));
	notech_inv i_33585(.A(n_6639), .Z(n_33632));
	notech_inv i_33586(.A(n_6642), .Z(n_33633));
	notech_inv i_33587(.A(n_5294), .Z(n_33634));
	notech_inv i_33588(.A(n_6641), .Z(n_33635));
	notech_inv i_33589(.A(n_6644), .Z(n_33636));
	notech_inv i_33590(.A(n_5295), .Z(n_33637));
	notech_inv i_33591(.A(n_6643), .Z(n_33638));
	notech_inv i_33592(.A(n_6646), .Z(n_33639));
	notech_inv i_33593(.A(n_5296), .Z(n_33640));
	notech_inv i_33594(.A(n_6645), .Z(n_33641));
	notech_inv i_33595(.A(n_6648), .Z(n_33642));
	notech_inv i_33596(.A(n_5297), .Z(n_33643));
	notech_inv i_33597(.A(n_6647), .Z(n_33644));
	notech_inv i_33598(.A(n_6650), .Z(n_33645));
	notech_inv i_33599(.A(n_5298), .Z(n_33646));
	notech_inv i_33600(.A(n_6649), .Z(n_33647));
	notech_inv i_33601(.A(n_6652), .Z(n_33648));
	notech_inv i_33602(.A(n_5299), .Z(n_33649));
	notech_inv i_33603(.A(n_6651), .Z(n_33650));
	notech_inv i_33604(.A(n_6654), .Z(n_33651));
	notech_inv i_33605(.A(n_5300), .Z(n_33652));
	notech_inv i_33606(.A(n_6653), .Z(n_33653));
	notech_inv i_33607(.A(n_6656), .Z(n_33654));
	notech_inv i_33608(.A(n_5301), .Z(n_33655));
	notech_inv i_33609(.A(n_6655), .Z(n_33656));
	notech_inv i_33610(.A(n_6658), .Z(n_33657));
	notech_inv i_33611(.A(n_5302), .Z(n_33658));
	notech_inv i_33612(.A(n_6657), .Z(n_33659));
	notech_inv i_33613(.A(n_6660), .Z(n_33660));
	notech_inv i_33614(.A(n_5303), .Z(n_33661));
	notech_inv i_33615(.A(n_6659), .Z(n_33662));
	notech_inv i_33616(.A(n_6662), .Z(n_33663));
	notech_inv i_33617(.A(n_5304), .Z(n_33664));
	notech_inv i_33618(.A(n_6661), .Z(n_33665));
	notech_inv i_33619(.A(n_6664), .Z(n_33666));
	notech_inv i_33620(.A(n_5305), .Z(n_33667));
	notech_inv i_33621(.A(n_6663), .Z(n_33668));
	notech_inv i_33622(.A(n_6666), .Z(n_33669));
	notech_inv i_33623(.A(n_5306), .Z(n_33670));
	notech_inv i_33624(.A(n_6665), .Z(n_33671));
	notech_inv i_33625(.A(n_6668), .Z(n_33672));
	notech_inv i_33626(.A(n_5307), .Z(n_33673));
	notech_inv i_33627(.A(n_6667), .Z(n_33674));
	notech_inv i_33628(.A(n_6670), .Z(n_33675));
	notech_inv i_33629(.A(n_5308), .Z(n_33676));
	notech_inv i_33630(.A(n_6669), .Z(n_33677));
	notech_inv i_33631(.A(n_6672), .Z(n_33678));
	notech_inv i_33632(.A(n_5309), .Z(n_33679));
	notech_inv i_33633(.A(n_6671), .Z(n_33680));
	notech_inv i_33634(.A(n_6674), .Z(n_33681));
	notech_inv i_33635(.A(n_5310), .Z(n_33682));
	notech_inv i_33636(.A(n_6673), .Z(n_33683));
	notech_inv i_33637(.A(n_6676), .Z(n_33684));
	notech_inv i_33638(.A(n_5311), .Z(n_33685));
	notech_inv i_33639(.A(n_6675), .Z(n_33686));
	notech_inv i_33640(.A(\opa_1[2] ), .Z(n_33687));
	notech_inv i_33641(.A(n_6261), .Z(n_33688));
	notech_inv i_33642(.A(mul64[63]), .Z(n_33689));
	notech_inv i_33643(.A(mul64[62]), .Z(n_33690));
	notech_inv i_33644(.A(mul64[61]), .Z(n_33691));
	notech_inv i_33645(.A(mul64[59]), .Z(n_33692));
	notech_inv i_33646(.A(mul64[58]), .Z(n_33693));
	notech_inv i_33647(.A(mul64[57]), .Z(n_33694));
	notech_inv i_33648(.A(mul64[56]), .Z(n_33695));
	notech_inv i_33649(.A(mul64[55]), .Z(n_33696));
	notech_inv i_33650(.A(mul64[54]), .Z(n_33697));
	notech_inv i_33651(.A(mul64[53]), .Z(n_33698));
	notech_inv i_33652(.A(mul64[52]), .Z(n_33699));
	notech_inv i_33653(.A(mul64[51]), .Z(n_33700));
	notech_inv i_33654(.A(mul64[50]), .Z(n_33701));
	notech_inv i_33655(.A(mul64[49]), .Z(n_33702));
	notech_inv i_33656(.A(mul64[48]), .Z(n_33703));
	notech_inv i_33657(.A(mul64[46]), .Z(n_33704));
	notech_inv i_33658(.A(mul64[45]), .Z(n_33705));
	notech_inv i_33659(.A(mul64[44]), .Z(n_33706));
	notech_inv i_33660(.A(mul64[43]), .Z(n_33707));
	notech_inv i_33661(.A(mul64[42]), .Z(n_33708));
	notech_inv i_33662(.A(mul64[41]), .Z(n_33709));
	notech_inv i_33663(.A(mul64[40]), .Z(n_33710));
	notech_inv i_33664(.A(mul64[35]), .Z(n_33711));
	notech_inv i_33665(.A(mul64[34]), .Z(n_33712));
	notech_inv i_33666(.A(mul64[33]), .Z(n_33713));
	notech_inv i_33667(.A(mul64[32]), .Z(n_33714));
	notech_inv i_33668(.A(mul64[60]), .Z(n_33715));
	notech_inv i_33669(.A(mul64[47]), .Z(n_33716));
	notech_inv i_33670(.A(n_538), .Z(n_33717));
	notech_inv i_33671(.A(n_3582), .Z(n_33718));
	notech_inv i_33672(.A(n_3569), .Z(n_33719));
	notech_inv i_33673(.A(n_3566), .Z(n_33720));
	notech_inv i_33674(.A(n_3562), .Z(n_33721));
	notech_inv i_33675(.A(n_3561), .Z(n_33722));
	notech_inv i_33676(.A(n_3560), .Z(n_33723));
	notech_inv i_33677(.A(n_3559), .Z(n_33724));
	notech_inv i_33678(.A(n_3558), .Z(n_33725));
	notech_inv i_33679(.A(n_3553), .Z(n_33726));
	notech_inv i_33680(.A(n_3549), .Z(n_33727));
	notech_inv i_33681(.A(n_3548), .Z(n_33728));
	notech_inv i_33682(.A(n_3547), .Z(n_33729));
	notech_inv i_33683(.A(n_3546), .Z(n_33730));
	notech_inv i_33684(.A(n_3545), .Z(n_33731));
	notech_inv i_33686(.A(n_3544), .Z(n_33732));
	notech_inv i_33687(.A(n_3543), .Z(n_33733));
	notech_inv i_33688(.A(n_3542), .Z(n_33734));
	notech_inv i_33689(.A(n_3540), .Z(n_33735));
	notech_inv i_33690(.A(n_3539), .Z(n_33736));
	notech_inv i_33691(.A(n_3537), .Z(n_33737));
	notech_inv i_33692(.A(n_3536), .Z(n_33738));
	notech_inv i_33693(.A(n_3535), .Z(n_33739));
	notech_inv i_33694(.A(n_3533), .Z(n_33740));
	notech_inv i_33695(.A(n_3532), .Z(n_33741));
	notech_inv i_33696(.A(n_4647), .Z(n_33742));
	notech_inv i_33697(.A(n_4648), .Z(n_33743));
	notech_inv i_33698(.A(n_4649), .Z(n_33744));
	notech_inv i_33699(.A(n_4622), .Z(n_33745));
	notech_inv i_33700(.A(n_4623), .Z(n_33746));
	notech_inv i_33701(.A(n_4624), .Z(n_33747));
	notech_inv i_33702(.A(n_4617), .Z(n_33748));
	notech_inv i_33703(.A(n_4618), .Z(n_33749));
	notech_inv i_33704(.A(n_4619), .Z(n_33750));
	notech_inv i_33705(.A(n_4612), .Z(n_33751));
	notech_inv i_33706(.A(n_4613), .Z(n_33752));
	notech_inv i_33707(.A(n_4614), .Z(n_33753));
	notech_inv i_33708(.A(n_543), .Z(n_33754));
	notech_inv i_33710(.A(n_4717), .Z(n_33755));
	notech_inv i_33711(.A(n_4718), .Z(n_33756));
	notech_inv i_33712(.A(n_4719), .Z(n_33757));
	notech_inv i_33713(.A(n_2707), .Z(n_33758));
	notech_inv i_33714(.A(n_6616), .Z(n_33759));
	notech_inv i_33715(.A(n_5281), .Z(n_33760));
	notech_inv i_33716(.A(n_6615), .Z(n_33761));
	notech_inv i_33717(.A(nCF_arithbox), .Z(n_33762));
	notech_inv i_33718(.A(nCF_shiftbox), .Z(n_33763));
	notech_inv i_33719(.A(\opc_1[0] ), .Z(n_33764));
	notech_inv i_33720(.A(n_3682), .Z(n_33765));
	notech_inv i_33721(.A(n_3649), .Z(n_33766));
	notech_inv i_33722(.A(\opc_1[1] ), .Z(n_33767));
	notech_inv i_33723(.A(n_3650), .Z(n_33768));
	notech_inv i_33724(.A(\opc_1[2] ), .Z(n_33769));
	notech_inv i_33725(.A(n_3684), .Z(n_33770));
	notech_inv i_33726(.A(n_3651), .Z(n_33771));
	notech_inv i_33727(.A(\opc_1[3] ), .Z(n_33772));
	notech_inv i_33729(.A(n_3685), .Z(n_33773));
	notech_inv i_33730(.A(n_3652), .Z(n_33774));
	notech_inv i_33731(.A(\opc_5[8] ), .Z(n_33775));
	notech_inv i_33732(.A(\opc_5[9] ), .Z(n_33776));
	notech_inv i_33733(.A(\opc_5[10] ), .Z(n_33777));
	notech_inv i_33734(.A(\opc_5[11] ), .Z(n_33778));
	notech_inv i_33735(.A(\opc_5[12] ), .Z(n_33779));
	notech_inv i_33736(.A(\opc_5[13] ), .Z(n_33780));
	notech_inv i_33737(.A(\opc_5[14] ), .Z(n_33781));
	notech_inv i_33738(.A(n_3665), .Z(n_33782));
	notech_inv i_33739(.A(n_3666), .Z(n_33783));
	notech_inv i_33740(.A(\opc_5[17] ), .Z(n_33784));
	notech_inv i_33741(.A(n_3667), .Z(n_33785));
	notech_inv i_33742(.A(\opc_5[18] ), .Z(n_33786));
	notech_inv i_33743(.A(n_3668), .Z(n_33787));
	notech_inv i_33744(.A(\opc_5[19] ), .Z(n_33788));
	notech_inv i_33745(.A(n_3669), .Z(n_33789));
	notech_inv i_33746(.A(\opc_5[20] ), .Z(n_33790));
	notech_inv i_33747(.A(n_3670), .Z(n_33791));
	notech_inv i_33748(.A(\opc_5[21] ), .Z(n_33792));
	notech_inv i_33750(.A(n_3671), .Z(n_33793));
	notech_inv i_33751(.A(\opc_5[22] ), .Z(n_33794));
	notech_inv i_33752(.A(n_3672), .Z(n_33795));
	notech_inv i_33753(.A(\opc_5[23] ), .Z(n_33796));
	notech_inv i_33754(.A(n_3673), .Z(n_33797));
	notech_inv i_33755(.A(\opc_5[24] ), .Z(n_33798));
	notech_inv i_33756(.A(n_3674), .Z(n_33799));
	notech_inv i_33757(.A(\opc_5[25] ), .Z(n_33800));
	notech_inv i_33758(.A(n_3675), .Z(n_33801));
	notech_inv i_33759(.A(\opc_5[26] ), .Z(n_33802));
	notech_inv i_33760(.A(n_3676), .Z(n_33803));
	notech_inv i_33761(.A(\opc_5[27] ), .Z(n_33804));
	notech_inv i_33762(.A(n_3678), .Z(n_33805));
	notech_inv i_33763(.A(\opc_5[29] ), .Z(n_33806));
	notech_inv i_33764(.A(n_3679), .Z(n_33807));
	notech_inv i_33765(.A(\opc_5[30] ), .Z(n_33808));
	notech_inv i_33766(.A(n_3680), .Z(n_33809));
	notech_inv i_33767(.A(\opc_5[31] ), .Z(n_33810));
	notech_inv i_33768(.A(n_4724), .Z(n_33811));
	notech_inv i_33769(.A(\nbus_11309[30] ), .Z(n_33812));
	notech_inv i_33770(.A(n_4722), .Z(n_33813));
	notech_inv i_33771(.A(n_4723), .Z(n_33814));
	notech_inv i_33772(.A(n_585), .Z(n_33815));
	notech_inv i_33773(.A(n_3654), .Z(n_33816));
	notech_inv i_33774(.A(\opc_1[5] ), .Z(n_33817));
	notech_inv i_33775(.A(\opc_5[5] ), .Z(n_33818));
	notech_inv i_33776(.A(n_3655), .Z(n_33819));
	notech_inv i_33777(.A(\opc_1[6] ), .Z(n_33820));
	notech_inv i_33778(.A(\opc_5[6] ), .Z(n_33821));
	notech_inv i_33779(.A(n_3656), .Z(n_33822));
	notech_inv i_33780(.A(\opc_1[7] ), .Z(n_33823));
	notech_inv i_33781(.A(\opc_5[7] ), .Z(n_33824));
	notech_inv i_33782(.A(\opc_5[15] ), .Z(n_33825));
	notech_inv i_33783(.A(n_3664), .Z(n_33826));
	notech_inv i_33784(.A(\opc_5[28] ), .Z(n_33827));
	notech_inv i_33785(.A(n_3563), .Z(n_33828));
	notech_inv i_33786(.A(n_61451), .Z(n_33829));
	notech_inv i_33787(.A(n_6578), .Z(n_33830));
	notech_inv i_33788(.A(n_6577), .Z(n_33831));
	notech_inv i_33789(.A(n_6576), .Z(n_33832));
	notech_inv i_33790(.A(n_6575), .Z(n_33833));
	notech_inv i_33791(.A(n_6574), .Z(n_33834));
	notech_inv i_33792(.A(n_6573), .Z(n_33835));
	notech_inv i_33793(.A(n_6572), .Z(n_33836));
	notech_inv i_33794(.A(n_6571), .Z(n_33837));
	notech_inv i_33795(.A(n_6570), .Z(n_33838));
	notech_inv i_33796(.A(n_6569), .Z(n_33839));
	notech_inv i_33797(.A(n_6568), .Z(n_33840));
	notech_inv i_33798(.A(n_6567), .Z(n_33841));
	notech_inv i_33799(.A(n_6566), .Z(n_33842));
	notech_inv i_33800(.A(n_6565), .Z(n_33843));
	notech_inv i_33801(.A(n_6564), .Z(n_33844));
	notech_inv i_33802(.A(n_6563), .Z(n_33845));
	notech_inv i_33803(.A(n_6562), .Z(n_33846));
	notech_inv i_33804(.A(n_6561), .Z(n_33847));
	notech_inv i_33805(.A(n_6560), .Z(n_33848));
	notech_inv i_33806(.A(n_6559), .Z(n_33849));
	notech_inv i_33807(.A(n_6558), .Z(n_33850));
	notech_inv i_33808(.A(n_6557), .Z(n_33851));
	notech_inv i_33809(.A(n_6556), .Z(n_33852));
	notech_inv i_33810(.A(n_6555), .Z(n_33853));
	notech_inv i_33811(.A(n_6554), .Z(n_33854));
	notech_inv i_33812(.A(n_6553), .Z(n_33855));
	notech_inv i_33813(.A(n_6552), .Z(n_33856));
	notech_inv i_33814(.A(n_6551), .Z(n_33857));
	notech_inv i_33815(.A(n_6550), .Z(n_33858));
	notech_inv i_33816(.A(n_6549), .Z(n_33859));
	notech_inv i_33817(.A(n_6548), .Z(n_33860));
	notech_inv i_33818(.A(n_6547), .Z(n_33861));
	notech_inv i_33819(.A(n_6546), .Z(n_33862));
	notech_inv i_33820(.A(n_6545), .Z(n_33863));
	notech_inv i_33821(.A(n_6544), .Z(n_33864));
	notech_inv i_33822(.A(n_6543), .Z(n_33865));
	notech_inv i_33823(.A(n_6542), .Z(n_33866));
	notech_inv i_33824(.A(n_6541), .Z(n_33867));
	notech_inv i_33825(.A(n_6540), .Z(n_33868));
	notech_inv i_33826(.A(n_6539), .Z(n_33869));
	notech_inv i_33827(.A(n_6538), .Z(n_33870));
	notech_inv i_33828(.A(n_6537), .Z(n_33871));
	notech_inv i_33829(.A(n_6536), .Z(n_33872));
	notech_inv i_33830(.A(n_6535), .Z(n_33873));
	notech_inv i_33831(.A(n_6534), .Z(n_33874));
	notech_inv i_33832(.A(n_6533), .Z(n_33875));
	notech_inv i_33833(.A(n_6532), .Z(n_33876));
	notech_inv i_33834(.A(n_6531), .Z(n_33877));
	notech_inv i_33835(.A(n_6530), .Z(n_33878));
	notech_inv i_33836(.A(n_6529), .Z(n_33879));
	notech_inv i_33837(.A(n_6528), .Z(n_33880));
	notech_inv i_33838(.A(n_6527), .Z(n_33881));
	notech_inv i_33839(.A(n_6526), .Z(n_33882));
	notech_inv i_33840(.A(n_6525), .Z(n_33883));
	notech_inv i_33841(.A(n_6524), .Z(n_33884));
	notech_inv i_33842(.A(n_6523), .Z(n_33885));
	notech_inv i_33843(.A(n_6522), .Z(n_33886));
	notech_inv i_33844(.A(n_6521), .Z(n_33887));
	notech_inv i_33845(.A(n_6520), .Z(n_33888));
	notech_inv i_33846(.A(n_6519), .Z(n_33889));
	notech_inv i_33847(.A(n_6518), .Z(n_33890));
	notech_inv i_33848(.A(n_6517), .Z(n_33891));
	notech_inv i_33849(.A(n_6516), .Z(n_33892));
	notech_inv i_33850(.A(n_6515), .Z(n_33893));
	notech_inv i_33851(.A(n_6450), .Z(n_33894));
	notech_inv i_33852(.A(n_6449), .Z(n_33895));
	notech_inv i_33853(.A(n_6448), .Z(n_33896));
	notech_inv i_33854(.A(n_6447), .Z(n_33897));
	notech_inv i_33855(.A(n_6446), .Z(n_33898));
	notech_inv i_33856(.A(n_6445), .Z(n_33899));
	notech_inv i_33857(.A(n_6444), .Z(n_33900));
	notech_inv i_33858(.A(n_6443), .Z(n_33901));
	notech_inv i_33859(.A(n_6442), .Z(n_33902));
	notech_inv i_33860(.A(n_6441), .Z(n_33903));
	notech_inv i_33861(.A(n_6440), .Z(n_33904));
	notech_inv i_33862(.A(n_6439), .Z(n_33905));
	notech_inv i_33863(.A(n_6438), .Z(n_33906));
	notech_inv i_33864(.A(n_6437), .Z(n_33907));
	notech_inv i_33865(.A(n_6436), .Z(n_33908));
	notech_inv i_33866(.A(n_6435), .Z(n_33909));
	notech_inv i_33867(.A(n_6434), .Z(n_33910));
	notech_inv i_33868(.A(n_6433), .Z(n_33911));
	notech_inv i_33869(.A(n_6432), .Z(n_33912));
	notech_inv i_33870(.A(n_6431), .Z(n_33913));
	notech_inv i_33871(.A(n_6430), .Z(n_33914));
	notech_inv i_33872(.A(n_6429), .Z(n_33915));
	notech_inv i_33873(.A(n_6428), .Z(n_33916));
	notech_inv i_33874(.A(n_6427), .Z(n_33917));
	notech_inv i_33875(.A(n_6426), .Z(n_33918));
	notech_inv i_33876(.A(n_6425), .Z(n_33919));
	notech_inv i_33877(.A(n_6424), .Z(n_33920));
	notech_inv i_33878(.A(n_6423), .Z(n_33921));
	notech_inv i_33879(.A(n_6422), .Z(n_33922));
	notech_inv i_33880(.A(n_6421), .Z(n_33923));
	notech_inv i_33881(.A(n_6420), .Z(n_33924));
	notech_inv i_33882(.A(n_6419), .Z(n_33925));
	notech_inv i_33883(.A(n_6514), .Z(n_33926));
	notech_inv i_33884(.A(n_6513), .Z(n_33927));
	notech_inv i_33885(.A(n_6512), .Z(n_33928));
	notech_inv i_33886(.A(n_6511), .Z(n_33929));
	notech_inv i_33887(.A(n_6510), .Z(n_33930));
	notech_inv i_33888(.A(n_6509), .Z(n_33931));
	notech_inv i_33889(.A(n_6508), .Z(n_33932));
	notech_inv i_33890(.A(n_6507), .Z(n_33933));
	notech_inv i_33891(.A(n_6506), .Z(n_33934));
	notech_inv i_33892(.A(n_6505), .Z(n_33935));
	notech_inv i_33893(.A(n_6504), .Z(n_33936));
	notech_inv i_33894(.A(n_6503), .Z(n_33937));
	notech_inv i_33895(.A(n_6502), .Z(n_33938));
	notech_inv i_33896(.A(n_6501), .Z(n_33939));
	notech_inv i_33897(.A(n_6500), .Z(n_33940));
	notech_inv i_33898(.A(n_6499), .Z(n_33941));
	notech_inv i_33899(.A(n_6498), .Z(n_33942));
	notech_inv i_33900(.A(n_6497), .Z(n_33943));
	notech_inv i_33901(.A(n_6496), .Z(n_33944));
	notech_inv i_33902(.A(n_6495), .Z(n_33945));
	notech_inv i_33903(.A(n_6494), .Z(n_33946));
	notech_inv i_33904(.A(n_6493), .Z(n_33947));
	notech_inv i_33905(.A(n_6492), .Z(n_33948));
	notech_inv i_33906(.A(n_6491), .Z(n_33949));
	notech_inv i_33907(.A(n_6490), .Z(n_33950));
	notech_inv i_33908(.A(n_6489), .Z(n_33951));
	notech_inv i_33909(.A(n_6488), .Z(n_33952));
	notech_inv i_33910(.A(n_6487), .Z(n_33953));
	notech_inv i_33911(.A(n_6486), .Z(n_33954));
	notech_inv i_33912(.A(n_6485), .Z(n_33955));
	notech_inv i_33913(.A(n_6484), .Z(n_33956));
	notech_inv i_33914(.A(n_6483), .Z(n_33957));
	notech_inv i_33916(.A(n_6482), .Z(n_33958));
	notech_inv i_33917(.A(n_6481), .Z(n_33959));
	notech_inv i_33918(.A(n_6480), .Z(n_33960));
	notech_inv i_33919(.A(n_6479), .Z(n_33961));
	notech_inv i_33920(.A(n_6478), .Z(n_33962));
	notech_inv i_33921(.A(n_6477), .Z(n_33963));
	notech_inv i_33922(.A(n_6476), .Z(n_33964));
	notech_inv i_33923(.A(n_6475), .Z(n_33965));
	notech_inv i_33924(.A(n_6474), .Z(n_33966));
	notech_inv i_33925(.A(n_6473), .Z(n_33967));
	notech_inv i_33926(.A(n_6472), .Z(n_33968));
	notech_inv i_33927(.A(n_6471), .Z(n_33969));
	notech_inv i_33928(.A(n_6470), .Z(n_33970));
	notech_inv i_33929(.A(n_6469), .Z(n_33971));
	notech_inv i_33930(.A(n_6468), .Z(n_33972));
	notech_inv i_33931(.A(n_6467), .Z(n_33973));
	notech_inv i_33932(.A(n_6466), .Z(n_33974));
	notech_inv i_33933(.A(n_6465), .Z(n_33975));
	notech_inv i_33934(.A(n_6464), .Z(n_33976));
	notech_inv i_33935(.A(n_6463), .Z(n_33977));
	notech_inv i_33936(.A(n_6462), .Z(n_33978));
	notech_inv i_33937(.A(n_6461), .Z(n_33979));
	notech_inv i_33938(.A(n_6460), .Z(n_33980));
	notech_inv i_33939(.A(n_6459), .Z(n_33981));
	notech_inv i_33940(.A(n_6458), .Z(n_33982));
	notech_inv i_33941(.A(n_6457), .Z(n_33983));
	notech_inv i_33942(.A(n_6456), .Z(n_33984));
	notech_inv i_33943(.A(n_6455), .Z(n_33985));
	notech_inv i_33944(.A(n_6454), .Z(n_33986));
	notech_inv i_33945(.A(n_6453), .Z(n_33987));
	notech_inv i_33946(.A(n_6452), .Z(n_33988));
	notech_inv i_33947(.A(n_6451), .Z(n_33989));
	AWMUX_16_32_7 i_32723(.I0(regs_0), .I1(ecx), .I2(regs_2), .I3(regs_3), .I4
		(regs_4), .I5(regs_5), .I6(regs_6), .I7(regs_7), .I8(regs_8), .I9
		({\nbus_14543[31] , \nbus_14543[30] , \nbus_14543[29] , \nbus_14543[28] 
		, \nbus_14543[27] , \nbus_14543[26] , \nbus_14543[25] , \nbus_14543[24] 
		, \nbus_14543[23] , \nbus_14543[22] , \nbus_14543[21] , \nbus_14543[20] 
		, \nbus_14543[19] , \nbus_14543[18] , \nbus_14543[17] , \nbus_14543[16] 
		, \nbus_14543[15] , \nbus_14543[14] , \nbus_14543[13] , \nbus_14543[12] 
		, \nbus_14543[11] , \nbus_14543[10] , \nbus_14543[9] , \nbus_14543[8] 
		, \nbus_14543[7] , \nbus_14543[6] , \nbus_14543[5] , \nbus_14543[4] 
		, \nbus_14543[3] , \nbus_14543[2] , cs[1], cs[0]}), .I10(regs_10
		), .I11(regs_11), .I12(regs_12), .I13({gs[31], gs[30], gs[29], gs
		[28], gs[27], gs[26], gs[25], gs[24], gs[23], gs[22], gs[21], gs
		[20], gs[19], gs[18], gs[17], gs[16], gs[15], gs[14], gs[13], gs
		[12], gs[11], gs[10], gs[9], gs[8], gs[7], gs[6], gs[5], gs[4], gs
		[3], n_56947, gs[1], gs[0]}), .I14(regs_14), .I15({\eflags[31] ,
		 \eflags[30] , \eflags[29] , \eflags[28] , \eflags[27] , \eflags[26] 
		, \eflags[25] , \eflags[24] , \eflags[23] , \eflags[22] , \eflags[21] 
		, \eflags[20] , \eflags[19] , \eflags[18] , \eflags[17] , \eflags[16] 
		, \eflags[15] , \eflags[14] , \eflags[13] , \eflags[12] , \eflags[11] 
		, \eflags[10] , ie, \eflags[8] , \eflags[7] , \eflags[6] , \eflags[5] 
		, \eflags[4] , \eflags[3] , \eflags[2] , \eflags[1] , \eflags[0] 
		}), .S({instrc[107], n_58201, instrc[105], instrc[104]}), .O0({n_6450
		, n_6449, n_6448, n_6447, n_6446, n_6445, n_6444, n_6443, n_6442
		, n_6441, n_6440, n_6439, n_6438, n_6437, n_6436, n_6435, n_6434
		, n_6433, n_6432, n_6431, n_6430, n_6429, n_6428, n_6427, n_6426
		, n_6425, n_6424, n_6423, n_6422, n_6421, n_6420, n_6419}));
	AWMUX_16_32_6 i_32728(.I0(regs_0), .I1(ecx), .I2(regs_2), .I3(regs_3), .I4
		(regs_4), .I5(regs_5), .I6(regs_6), .I7(regs_7), .I8(regs_8), .I9
		({\nbus_14543[31] , \nbus_14543[30] , \nbus_14543[29] , \nbus_14543[28] 
		, \nbus_14543[27] , \nbus_14543[26] , \nbus_14543[25] , \nbus_14543[24] 
		, \nbus_14543[23] , \nbus_14543[22] , \nbus_14543[21] , \nbus_14543[20] 
		, \nbus_14543[19] , \nbus_14543[18] , \nbus_14543[17] , \nbus_14543[16] 
		, \nbus_14543[15] , \nbus_14543[14] , \nbus_14543[13] , \nbus_14543[12] 
		, \nbus_14543[11] , \nbus_14543[10] , \nbus_14543[9] , \nbus_14543[8] 
		, \nbus_14543[7] , \nbus_14543[6] , \nbus_14543[5] , \nbus_14543[4] 
		, \nbus_14543[3] , \nbus_14543[2] , cs[1], cs[0]}), .I10(regs_10
		), .I11(regs_11), .I12(regs_12), .I13({gs[31], gs[30], gs[29], gs
		[28], gs[27], gs[26], gs[25], gs[24], gs[23], gs[22], gs[21], gs
		[20], gs[19], gs[18], gs[17], gs[16], gs[15], gs[14], gs[13], gs
		[12], gs[11], gs[10], gs[9], gs[8], gs[7], gs[6], gs[5], gs[4], gs
		[3], n_56947, gs[1], gs[0]}), .I14(regs_14), .I15({\eflags[31] ,
		 \eflags[30] , \eflags[29] , \eflags[28] , \eflags[27] , \eflags[26] 
		, \eflags[25] , \eflags[24] , \eflags[23] , \eflags[22] , \eflags[21] 
		, \eflags[20] , \eflags[19] , \eflags[18] , \eflags[17] , \eflags[16] 
		, \eflags[15] , \eflags[14] , \eflags[13] , \eflags[12] , \eflags[11] 
		, \eflags[10] , ie, \eflags[8] , \eflags[7] , \eflags[6] , \eflags[5] 
		, \eflags[4] , \eflags[3] , \eflags[2] , \eflags[1] , \eflags[0] 
		}), .S({instrc[103], instrc[102], instrc[101], instrc[100]}), .O0
		({n_6482, n_6481, n_6480, n_6479, n_6478, n_6477, n_6476, n_6475
		, n_6474, n_6473, n_6472, n_6471, n_6470, n_6469, n_6468, n_6467
		, n_6466, n_6465, n_6464, n_6463, n_6462, n_6461, n_6460, n_6459
		, n_6458, n_6457, n_6456, n_6455, n_6454, n_6453, n_6452, n_6451
		}));
	AWMUX_16_32_5 i_32733(.I0(regs_0), .I1(ecx), .I2(regs_2), .I3(regs_3), .I4
		(regs_4), .I5(regs_5), .I6(regs_6), .I7(regs_7), .I8(regs_8), .I9
		({\nbus_14543[31] , \nbus_14543[30] , \nbus_14543[29] , \nbus_14543[28] 
		, \nbus_14543[27] , \nbus_14543[26] , \nbus_14543[25] , \nbus_14543[24] 
		, \nbus_14543[23] , \nbus_14543[22] , \nbus_14543[21] , \nbus_14543[20] 
		, \nbus_14543[19] , \nbus_14543[18] , \nbus_14543[17] , \nbus_14543[16] 
		, \nbus_14543[15] , \nbus_14543[14] , \nbus_14543[13] , \nbus_14543[12] 
		, \nbus_14543[11] , \nbus_14543[10] , \nbus_14543[9] , \nbus_14543[8] 
		, \nbus_14543[7] , \nbus_14543[6] , \nbus_14543[5] , \nbus_14543[4] 
		, \nbus_14543[3] , \nbus_14543[2] , cs[1], cs[0]}), .I10(regs_10
		), .I11(regs_11), .I12(regs_12), .I13({gs[31], gs[30], gs[29], gs
		[28], gs[27], gs[26], gs[25], gs[24], gs[23], gs[22], gs[21], gs
		[20], gs[19], gs[18], gs[17], gs[16], gs[15], gs[14], gs[13], gs
		[12], gs[11], gs[10], gs[9], gs[8], gs[7], gs[6], gs[5], gs[4], gs
		[3], n_56947, gs[1], gs[0]}), .I14(regs_14), .I15({\eflags[31] ,
		 \eflags[30] , \eflags[29] , \eflags[28] , \eflags[27] , \eflags[26] 
		, \eflags[25] , \eflags[24] , \eflags[23] , \eflags[22] , \eflags[21] 
		, \eflags[20] , \eflags[19] , \eflags[18] , \eflags[17] , \eflags[16] 
		, \eflags[15] , \eflags[14] , \eflags[13] , \eflags[12] , \eflags[11] 
		, \eflags[10] , ie, \eflags[8] , \eflags[7] , \eflags[6] , \eflags[5] 
		, \eflags[4] , \eflags[3] , \eflags[2] , \eflags[1] , \eflags[0] 
		}), .S({instrc[99], instrc[98], instrc[97], instrc[96]}), .O0({n_6514
		, n_6513, n_6512, n_6511, n_6510, n_6509, n_6508, n_6507, n_6506
		, n_6505, n_6504, n_6503, n_6502, n_6501, n_6500, n_6499, n_6498
		, n_6497, n_6496, n_6495, n_6494, n_6493, n_6492, n_6491, n_6490
		, n_6489, n_6488, n_6487, n_6486, n_6485, n_6484, n_6483}));
	AWMUX_16_32_4 i_32738(.I0(regs_0), .I1(ecx), .I2(regs_2), .I3(regs_3), .I4
		(regs_4), .I5(regs_5), .I6(regs_6), .I7(regs_7), .I8(regs_8), .I9
		({\nbus_14543[31] , \nbus_14543[30] , \nbus_14543[29] , \nbus_14543[28] 
		, \nbus_14543[27] , \nbus_14543[26] , \nbus_14543[25] , \nbus_14543[24] 
		, \nbus_14543[23] , \nbus_14543[22] , \nbus_14543[21] , \nbus_14543[20] 
		, \nbus_14543[19] , \nbus_14543[18] , \nbus_14543[17] , \nbus_14543[16] 
		, \nbus_14543[15] , \nbus_14543[14] , \nbus_14543[13] , \nbus_14543[12] 
		, \nbus_14543[11] , \nbus_14543[10] , \nbus_14543[9] , \nbus_14543[8] 
		, \nbus_14543[7] , \nbus_14543[6] , \nbus_14543[5] , \nbus_14543[4] 
		, \nbus_14543[3] , \nbus_14543[2] , cs[1], cs[0]}), .I10(regs_10
		), .I11(regs_11), .I12(regs_12), .I13({gs[31], gs[30], gs[29], gs
		[28], gs[27], gs[26], gs[25], gs[24], gs[23], gs[22], gs[21], gs
		[20], gs[19], gs[18], gs[17], gs[16], gs[15], gs[14], gs[13], gs
		[12], gs[11], gs[10], gs[9], gs[8], gs[7], gs[6], gs[5], gs[4], gs
		[3], n_56947, gs[1], gs[0]}), .I14(regs_14), .I15({\eflags[31] ,
		 \eflags[30] , \eflags[29] , \eflags[28] , \eflags[27] , \eflags[26] 
		, \eflags[25] , \eflags[24] , \eflags[23] , \eflags[22] , \eflags[21] 
		, \eflags[20] , \eflags[19] , \eflags[18] , \eflags[17] , \eflags[16] 
		, \eflags[15] , \eflags[14] , \eflags[13] , \eflags[12] , \eflags[11] 
		, \eflags[10] , ie, \eflags[8] , \eflags[7] , \eflags[6] , \eflags[5] 
		, \eflags[4] , \eflags[3] , \eflags[2] , \eflags[1] , \eflags[0] 
		}), .S({instrc[95], instrc[94], instrc[93], instrc[92]}), .O0({n_6546
		, n_6545, n_6544, n_6543, n_6542, n_6541, n_6540, n_6539, n_6538
		, n_6537, n_6536, n_6535, n_6534, n_6533, n_6532, n_6531, n_6530
		, n_6529, n_6528, n_6527, n_6526, n_6525, n_6524, n_6523, n_6522
		, n_6521, n_6520, n_6519, n_6518, n_6517, n_6516, n_6515}));
	AWMUX_16_32_3 i_32743(.I0(regs_0), .I1(ecx), .I2(regs_2), .I3(regs_3), .I4
		(regs_4), .I5(regs_5), .I6(regs_6), .I7(regs_7), .I8(regs_8), .I9
		({\nbus_14543[31] , \nbus_14543[30] , \nbus_14543[29] , \nbus_14543[28] 
		, \nbus_14543[27] , \nbus_14543[26] , \nbus_14543[25] , \nbus_14543[24] 
		, \nbus_14543[23] , \nbus_14543[22] , \nbus_14543[21] , \nbus_14543[20] 
		, \nbus_14543[19] , \nbus_14543[18] , \nbus_14543[17] , \nbus_14543[16] 
		, \nbus_14543[15] , \nbus_14543[14] , \nbus_14543[13] , \nbus_14543[12] 
		, \nbus_14543[11] , \nbus_14543[10] , \nbus_14543[9] , \nbus_14543[8] 
		, \nbus_14543[7] , \nbus_14543[6] , \nbus_14543[5] , \nbus_14543[4] 
		, \nbus_14543[3] , \nbus_14543[2] , cs[1], cs[0]}), .I10(regs_10
		), .I11(regs_11), .I12(regs_12), .I13({gs[31], gs[30], gs[29], gs
		[28], gs[27], gs[26], gs[25], gs[24], gs[23], gs[22], gs[21], gs
		[20], gs[19], gs[18], gs[17], gs[16], gs[15], gs[14], gs[13], gs
		[12], gs[11], gs[10], gs[9], gs[8], gs[7], gs[6], gs[5], gs[4], gs
		[3], n_56947, gs[1], gs[0]}), .I14(regs_14), .I15({\eflags[31] ,
		 \eflags[30] , \eflags[29] , \eflags[28] , \eflags[27] , \eflags[26] 
		, \eflags[25] , \eflags[24] , \eflags[23] , \eflags[22] , \eflags[21] 
		, \eflags[20] , \eflags[19] , \eflags[18] , \eflags[17] , \eflags[16] 
		, \eflags[15] , \eflags[14] , \eflags[13] , \eflags[12] , \eflags[11] 
		, \eflags[10] , ie, \eflags[8] , \eflags[7] , \eflags[6] , \eflags[5] 
		, \eflags[4] , \eflags[3] , \eflags[2] , \eflags[1] , \eflags[0] 
		}), .S({instrc[91], instrc[90], instrc[89], instrc[88]}), .O0({n_6578
		, n_6577, n_6576, n_6575, n_6574, n_6573, n_6572, n_6571, n_6570
		, n_6569, n_6568, n_6567, n_6566, n_6565, n_6564, n_6563, n_6562
		, n_6561, n_6560, n_6559, n_6558, n_6557, n_6556, n_6555, n_6554
		, n_6553, n_6552, n_6551, n_6550, n_6549, n_6548, n_6547}));
	AWMUX_16_32_2 i_32748(.I0(write_data_25), .I1(write_data_26), .I2(write_data_27
		), .I3(write_data_28), .I4(write_data_29), .I5(write_data_30), .I6
		(write_data_31), .I7(write_data_32), .S(all_cnt), .O0(write_data_33
		));
	AWMUX_16_32_1 i_55513(.I0(regs_0), .I1(ecx), .I2(regs_2), .I3(regs_3), .I4
		(regs_4), .I5(regs_5), .I6(regs_6), .I7(regs_7), .I8(regs_8), .I9
		({\nbus_14543[31] , \nbus_14543[30] , \nbus_14543[29] , \nbus_14543[28] 
		, \nbus_14543[27] , \nbus_14543[26] , \nbus_14543[25] , \nbus_14543[24] 
		, \nbus_14543[23] , \nbus_14543[22] , \nbus_14543[21] , \nbus_14543[20] 
		, \nbus_14543[19] , \nbus_14543[18] , \nbus_14543[17] , \nbus_14543[16] 
		, \nbus_14543[15] , \nbus_14543[14] , \nbus_14543[13] , \nbus_14543[12] 
		, \nbus_14543[11] , \nbus_14543[10] , \nbus_14543[9] , \nbus_14543[8] 
		, \nbus_14543[7] , \nbus_14543[6] , \nbus_14543[5] , \nbus_14543[4] 
		, \nbus_14543[3] , \nbus_14543[2] , cs[1], cs[0]}), .I10(regs_10
		), .I11(regs_11), .I12(regs_12), .I13({gs[31], gs[30], gs[29], gs
		[28], gs[27], gs[26], gs[25], gs[24], gs[23], gs[22], gs[21], gs
		[20], gs[19], gs[18], gs[17], gs[16], gs[15], gs[14], gs[13], gs
		[12], gs[11], gs[10], gs[9], gs[8], gs[7], gs[6], gs[5], gs[4], gs
		[3], n_56947, gs[1], gs[0]}), .I14(regs_14), .I15({\eflags[31] ,
		 \eflags[30] , \eflags[29] , \eflags[28] , \eflags[27] , \eflags[26] 
		, \eflags[25] , \eflags[24] , \eflags[23] , \eflags[22] , \eflags[21] 
		, \eflags[20] , \eflags[19] , \eflags[18] , \eflags[17] , \eflags[16] 
		, \eflags[15] , \eflags[14] , \eflags[13] , \eflags[12] , \eflags[11] 
		, \eflags[10] , ie, \eflags[8] , \eflags[7] , \eflags[6] , \eflags[5] 
		, \eflags[4] , \eflags[3] , \eflags[2] , \eflags[1] , \eflags[0] 
		}), .S({instrc[127], instrc[126], instrc[125], instrc[124]}), .O0
		({\regs_13_14[31] , \regs_13_14[30] , \regs_13_14[29] , \regs_13_14[28] 
		, \regs_13_14[27] , \regs_13_14[26] , \regs_13_14[25] , \regs_13_14[24] 
		, \regs_13_14[23] , \regs_13_14[22] , \regs_13_14[21] , \regs_13_14[20] 
		, \regs_13_14[19] , \regs_13_14[18] , \regs_13_14[17] , \regs_13_14[16] 
		, \opa_12[15] , \opa_12[14] , \opa_12[13] , \opa_12[12] , \opa_12[11] 
		, \opa_12[10] , \opa_12[9] , \opa_12[8] , \opa_12[7] , \opa_12[6] 
		, \opa_12[5] , \opa_12[4] , \opa_12[3] , \opa_12[2] , \opa_12[1] 
		, \opa_12[0] }));
	AWMUX_16_32_0 i_55867(.I0(regs_0), .I1(ecx), .I2(regs_2), .I3(regs_3), .I4
		(regs_4), .I5(regs_5), .I6(regs_6), .I7(regs_7), .I8(regs_8), .I9
		({\nbus_14543[31] , \nbus_14543[30] , \nbus_14543[29] , \nbus_14543[28] 
		, \nbus_14543[27] , \nbus_14543[26] , \nbus_14543[25] , \nbus_14543[24] 
		, \nbus_14543[23] , \nbus_14543[22] , \nbus_14543[21] , \nbus_14543[20] 
		, \nbus_14543[19] , \nbus_14543[18] , \nbus_14543[17] , \nbus_14543[16] 
		, \nbus_14543[15] , \nbus_14543[14] , \nbus_14543[13] , \nbus_14543[12] 
		, \nbus_14543[11] , \nbus_14543[10] , \nbus_14543[9] , \nbus_14543[8] 
		, \nbus_14543[7] , \nbus_14543[6] , \nbus_14543[5] , \nbus_14543[4] 
		, \nbus_14543[3] , \nbus_14543[2] , cs[1], cs[0]}), .I10(regs_10
		), .I11(regs_11), .I12(regs_12), .I13({gs[31], gs[30], gs[29], gs
		[28], gs[27], gs[26], gs[25], gs[24], gs[23], gs[22], gs[21], gs
		[20], gs[19], gs[18], gs[17], gs[16], gs[15], gs[14], gs[13], gs
		[12], gs[11], gs[10], gs[9], gs[8], gs[7], gs[6], gs[5], gs[4], gs
		[3], n_56947, gs[1], gs[0]}), .I14(regs_14), .I15({\eflags[31] ,
		 \eflags[30] , \eflags[29] , \eflags[28] , \eflags[27] , \eflags[26] 
		, \eflags[25] , \eflags[24] , \eflags[23] , \eflags[22] , \eflags[21] 
		, \eflags[20] , \eflags[19] , \eflags[18] , \eflags[17] , \eflags[16] 
		, \eflags[15] , \eflags[14] , \eflags[13] , \eflags[12] , \eflags[11] 
		, \eflags[10] , ie, \eflags[8] , \eflags[7] , \eflags[6] , \eflags[5] 
		, \eflags[4] , \eflags[3] , \eflags[2] , \eflags[1] , \eflags[0] 
		}), .S({n_57714, n_57705, n_57696, instrc[116]}), .O0(opc_10));
	AWDP_INC_0 i_1014(.O0({n_454, n_452, n_450, n_448, n_446, n_444, n_442, n_440
		, n_438, n_436, n_434, n_432, n_430, n_428, n_426, n_424, n_422,
		 n_420, n_418, n_416, n_414, n_412, n_410, n_408, n_406, n_404, n_402
		, n_400, n_398, n_396, n_394, n_392, n_390, n_388, n_386, n_384,
		 n_382, n_380, n_378, n_376, n_374, n_372, n_370, n_368, n_366, n_364
		, n_362, n_360, n_358, n_356, n_354, n_352, n_350, n_348, n_346,
		 n_344, n_342, n_340, n_338, n_336, n_334, n_332, n_330, n_328})
		, .tsc(tsc));
	AWDP_SUB_37 i_968(.O0(regs_4_2), .regs_4(regs_4), .calc_sz({calc_sz[2], calc_sz
		[1], calc_sz[0]}));
	AWDP_ADD_110 i_967(.O0({n_2738, n_2737, n_2736, n_2735, n_2734, n_2733, n_2732
		, n_2731, n_2730, n_2729, n_2728, n_2727, n_2726, n_2725, n_2724
		, n_2723, n_2722, n_2721, n_2720, n_2719, n_2718, n_2717, n_2716
		, n_2715, n_2714, n_2713, n_2712, n_2711, n_2710, n_2709, n_2708
		, n_2707}), .regs_4(regs_4), .calc_sz({calc_sz[2], calc_sz[1], calc_sz
		[0]}));
	AWDP_ADD_52 i_964(.O0({n_1769, n_1767, n_1765, n_1763, n_1761, n_1759, n_1757
		, n_1755, n_1753, n_1751, n_1749, n_1747, n_1745, n_1743, n_1741
		, n_1739, n_1737, n_1735, n_1733, n_1731, n_1729, n_1727, n_1725
		, n_1723, n_1721, n_1719, n_1717, n_1715, n_1713, n_1711, n_1709
		, n_1707}), .regs_7(regs_7), .opd({n_58018, opd[30], n_57937, n_57946
		, n_57956, n_57965, opd[25], opd[24], opd[23], opd[22], opd[21],
		 opd[20], opd[19], opd[18], opd[17], opd[16], opd[15], opd[14], opd
		[13], opd[12], opd[11], opd[10], opd[9], opd[8], opd[7], opd[6],
		 n_56982, opd[4], n_58783, opd[2], n_56955, n_56964}));
	AWDP_SUB_129 i_963(.O0({n_1770, n_1768, n_1766, n_1764, n_1762, n_1760, n_1758
		, n_1756, n_1754, n_1752, n_1750, n_1748, n_1746, n_1744, n_1742
		, n_1740, n_1738, n_1736, n_1734, n_1732, n_1730, n_1728, n_1726
		, n_1724, n_1722, n_1720, n_1718, n_1716, n_1714, n_1712, n_1710
		, n_1708}), .regs_7(regs_7), .opd({n_58018, opd[30], n_57937, n_57946
		, n_57956, n_57965, opd[25], opd[24], opd[23], opd[22], opd[21],
		 opd[20], opd[19], opd[18], opd[17], opd[16], opd[15], opd[14], opd
		[13], opd[12], opd[11], opd[10], opd[9], opd[8], opd[7], opd[6],
		 n_56982, n_56973, n_58783, n_58801, n_56955, n_56964}));
	shiftbox shiftbox(.shiftop({\opcode[3] , \opcode[2] , \opcode[1] , \opcode[0] 
		}), .calc_sz(calc_sz), .ci(\eflags[0] ), .co(nCF_shiftbox), .co4
		(nCF_shift4box), .opa({opa[31], opa[30], opa[29], opa[28], opa[
		27], opa[26], opa[25], opa[24], opa[23], opa[22], opa[21], opa[
		20], opa[19], opa[18], opa[17], opa[16], n_61034, opa[14], n_61025
		, n_61016, opa[11], opa[10], n_61007, opa[8], n_60998, n_60989, n_60980
		, opa[4], n_60971, n_60962, opa[1], opa[0]}), .opb({n_60629, opb
		[30], opb[29], opb[28], opb[27], opb[26], opb[25], opb[24], opb[
		23], opb[22], opb[21], opb[20], opb[19], opb[18], opb[17], opb[
		16], opb[15], opb[14], opb[13], opb[12], opb[11], opb[10], opb[9
		], opb[8], opb[7], opb[6], opb[5], opb[4], opb[3], opb[2], opb[1
		], opb[0]}), .resa(resa_shiftbox), .resb(resb_shiftbox), .resa4(resa_shift4box
		), .resb4(resb_shift4box));
	AWMUX_16_1 i_947(.I0(\eflags[11] ), .I2(\eflags[0] ), .I4(\eflags[6] ), 
		.I6(\cond[6] ), .I8(\eflags[7] ), .I10(\eflags[2] ), .I12(\cond[12] 
		), .I14(\cond[14] ), .S({n_63800, n_63728, n_63716, n_63818}), .O0
		(cond_1));
	AWDP_ADD_33 i_945(.add_len_pc32(add_len_pc32), .regs_14(regs_14), .lenpc
		(lenpc));
	AWDP_ADD_222 i_944(.add_len_pc16({n_533, n_532, n_531, n_530, n_529, n_528
		, n_527, n_526, n_525, n_524, n_523, n_522, n_521, n_520, n_519,
		 n_518}), .regs_14({regs_14[15], regs_14[14], regs_14[13], regs_14
		[12], regs_14[11], regs_14[10], regs_14[9], regs_14[8], regs_14[
		7], regs_14[6], regs_14[5], regs_14[4], regs_14[3], regs_14[2], regs_14
		[1], regs_14[0]}), .lenpc({lenpc[15], lenpc[14], lenpc[13], lenpc
		[12], lenpc[11], lenpc[10], lenpc[9], lenpc[8], lenpc[7], lenpc[
		6], lenpc[5], lenpc[4], lenpc[3], lenpc[2], lenpc[1], lenpc[0]})
		);
	AWDP_ADD_43 i_939(.O0({n_6792, n_6791, n_6790, n_6789, n_6788, n_6787, n_6786
		, n_6785, n_6784, n_6783, n_6782, n_6781, n_6780, n_6779, n_6778
		, n_6777, n_6776, n_6775, n_6774, n_6773, n_6772, n_6771, n_6770
		, n_6769, n_6768, n_6767, n_6766, n_6765, n_6764, n_6763, n_6762
		, n_6761}), .I0({\nbus_11309[31] , \nbus_11309[30] , \nbus_11309[29] 
		, \nbus_11309[28] , n_348189363, \nbus_11309[26] , n_348089362, \nbus_11309[24] 
		, \nbus_11309[23] , \nbus_11309[22] , n_347989361, n_347889360, n_347789359
		, \nbus_11309[18] , n_347689358, n_347589357, \nbus_11309[15] , n_351585923
		, n_351485922, n_351385921, n_351285920, \nbus_11309[10] , \nbus_11309[9] 
		, \nbus_11309[8] , n_351185919, n_351085918, n_350985917, \nbus_11309[4] 
		, n_350885916, n_350785915, n_350685914, n_350585913}), .add_len_pc
		({\add_len_pc[31] , \add_len_pc[30] , \add_len_pc[29] , \add_len_pc[28] 
		, \add_len_pc[27] , \add_len_pc[26] , n_3463, n_3462, n_3461, n_3460
		, n_3459, n_3458, \add_len_pc[19] , \add_len_pc[18] , \add_len_pc[17] 
		, \add_len_pc[16] , \add_len_pc[15] , \add_len_pc[14] , \add_len_pc[13] 
		, \add_len_pc[12] , \add_len_pc[11] , \add_len_pc[10] , \add_len_pc[9] 
		, \add_len_pc[8] , \add_len_pc[7] , \add_len_pc[6] , \add_len_pc[5] 
		, \add_len_pc[4] , \add_len_pc[3] , \add_len_pc[2] , \add_len_pc[1] 
		, \add_len_pc[0] }));
	AWDP_EQ_85 i_915(.O0({n_537}), .mul64({mul64[63], mul64[62], mul64[61], mul64
		[60], mul64[59], mul64[58], mul64[57], mul64[56], mul64[55], mul64
		[54], mul64[53], mul64[52], mul64[51], mul64[50], mul64[49], mul64
		[48], mul64[47], mul64[46], mul64[45], mul64[44], mul64[43], mul64
		[42], mul64[41], mul64[40], mul64[39], mul64[38], mul64[37], mul64
		[36], mul64[35], mul64[34], mul64[33], mul64[32], mul64[31], mul64
		[30], mul64[29], mul64[28], mul64[27], mul64[26], mul64[25], mul64
		[24], mul64[23], mul64[22], mul64[21], mul64[20], mul64[19], mul64
		[18], mul64[17], mul64[16], mul64[15], mul64[14], mul64[13], mul64
		[12], mul64[11], mul64[10], mul64[9], mul64[8]}));
	AWDP_EQ_174 i_914(.O0({n_538}), .mul64({mul64[63], mul64[62], mul64[61],
		 mul64[60], mul64[59], mul64[58], mul64[57], mul64[56], mul64[55
		], mul64[54], mul64[53], mul64[52], mul64[51], mul64[50], mul64[
		49], mul64[48], mul64[47], mul64[46], mul64[45], mul64[44], mul64
		[43], mul64[42], mul64[41], mul64[40], mul64[39], mul64[38], mul64
		[37], mul64[36], mul64[35], mul64[34], mul64[33], mul64[32], mul64
		[31], mul64[30], mul64[29], mul64[28], mul64[27], mul64[26], mul64
		[25], mul64[24], mul64[23], mul64[22], mul64[21], mul64[20], mul64
		[19], mul64[18], mul64[17], mul64[16]}));
	AWDP_EQ_91 i_911(.O0({n_541}), .mul64({mul64[63], mul64[62], mul64[61], mul64
		[60], mul64[59], mul64[58], mul64[57], mul64[56], mul64[55], mul64
		[54], mul64[53], mul64[52], mul64[51], mul64[50], mul64[49], mul64
		[48], mul64[47], mul64[46], mul64[45], mul64[44], mul64[43], mul64
		[42], mul64[41], mul64[40], mul64[39], mul64[38], mul64[37], mul64
		[36], mul64[35], mul64[34], mul64[33], mul64[32], mul64[31], mul64
		[30], mul64[29], mul64[28], mul64[27], mul64[26], mul64[25], mul64
		[24], mul64[23], mul64[22], mul64[21], mul64[20], mul64[19], mul64
		[18], mul64[17], mul64[16], mul64[15], mul64[14], mul64[13], mul64
		[12], mul64[11], mul64[10], mul64[9], mul64[8]}));
	AWDP_EQ_24111880 i_909(.O0({n_543}), .mul64({mul64[63], mul64[62], mul64
		[61], mul64[60], mul64[59], mul64[58], mul64[57], mul64[56], mul64
		[55], mul64[54], mul64[53], mul64[52], mul64[51], mul64[50], mul64
		[49], mul64[48], mul64[47], mul64[46], mul64[45], mul64[44], mul64
		[43], mul64[42], mul64[41], mul64[40], mul64[39], mul64[38], mul64
		[37], mul64[36], mul64[35], mul64[34], mul64[33], mul64[32], mul64
		[31], mul64[30], mul64[29], mul64[28], mul64[27], mul64[26], mul64
		[25], mul64[24], mul64[23], mul64[22], mul64[21], mul64[20], mul64
		[19], mul64[18], mul64[17], mul64[16]}));
	AWDP_EQ_205 i_907(.O0({n_545}), .mul64({mul64[63], mul64[62], mul64[61],
		 mul64[60], mul64[59], mul64[58], mul64[57], mul64[56], mul64[55
		], mul64[54], mul64[53], mul64[52], mul64[51], mul64[50], mul64[
		49], mul64[48], mul64[47], mul64[46], mul64[45], mul64[44], mul64
		[43], mul64[42], mul64[41], mul64[40], mul64[39], mul64[38], mul64
		[37], mul64[36], mul64[35], mul64[34], mul64[33], mul64[32]}));
	AWDP_ADD_6 i_901(.O0(nbus_133), .opa({opa[31], opa[30], opa[29], opa[28]
		, opa[27], opa[26], opa[25], opa[24], opa[23], opa[22], opa[21],
		 opa[20], opa[19], opa[18], opa[17], opa[16], n_61034, opa[14], n_61025
		, n_61016, opa[11], opa[10], n_61007, opa[8], n_60998, n_60989, n_60980
		, opa[4], n_60971, n_60962, opa[1], n_60953}), .opd({n_58018, opd
		[30], n_57937, n_57946, n_57956, n_57965, opd[25], opd[24], opd[
		23], opd[22], opd[21], opd[20], opd[19], opd[18], opd[17], opd[
		16], opd[15], opd[14], opd[13], opd[12], opd[11], opd[10], opd[9
		], opd[8], opd[7], opd[6], n_56982, n_56973, n_58783, n_58801, n_56955
		, n_56964}));
	AWDP_ADD_103 i_899(.O0(nbus_134), .opa({n_61034, opa[14], n_61025, n_61016
		, opa[11], opa[10], n_61007, opa[8], n_60998, n_60989, n_60980, opa
		[4], n_60971, n_60962, opa[1], n_60953}), .opd({opd[15], opd[14]
		, opd[13], opd[12], opd[11], opd[10], opd[9], opd[8], opd[7], opd
		[6], n_56982, n_56973, n_58783, n_58801, n_56955, n_56964}));
	AWDP_ADD_101 i_898(.O0(nbus_135), .opa({n_60998, n_60989, n_60980, opa[4
		], n_60971, n_60962, opa[1], n_60953}), .opd({opd[7], opd[6], n_56982
		, n_56973, n_58783, n_58801, n_56955, n_56964}));
	AWDP_ADD_123 i_897(.O0(nbus_136), .opb({n_60629, opb[30], opb[29], opb[
		28], opb[27], opb[26], opb[25], opb[24], opb[23], opb[22], opb[
		21], opb[20], opb[19], opb[18], opb[17], opb[16], opb[15], opb[
		14], opb[13], opb[12], opb[11], opb[10], opb[9], opb[8], opb[7],
		 opb[6], opb[5], opb[4], opb[3], opb[2], opb[1], opb[0]}), .I0({
		UNCONNECTED_000, UNCONNECTED_001, UNCONNECTED_002, 
		UNCONNECTED_003, UNCONNECTED_004, UNCONNECTED_005, 
		UNCONNECTED_006, UNCONNECTED_007, UNCONNECTED_008, 
		UNCONNECTED_009, UNCONNECTED_010, UNCONNECTED_011, 
		UNCONNECTED_012, n_58201, UNCONNECTED_013, UNCONNECTED_014, 
		UNCONNECTED_015, UNCONNECTED_016, UNCONNECTED_017, 
		UNCONNECTED_018, UNCONNECTED_019, UNCONNECTED_020, 
		UNCONNECTED_021, UNCONNECTED_022, UNCONNECTED_023, 
		UNCONNECTED_024, UNCONNECTED_025, UNCONNECTED_026, 
		UNCONNECTED_027, UNCONNECTED_028, instrc[105], instrc[104]}));
	AWDP_ADD_160 i_896(.O0(nbus_137), .opb({opb[15], opb[14], opb[13], opb[
		12], opb[11], opb[10], opb[9], opb[8], opb[7], opb[6], opb[5], opb
		[4], opb[3], opb[2], opb[1], opb[0]}), .I0({n_58206, 
		UNCONNECTED_029, UNCONNECTED_030, UNCONNECTED_031, 
		UNCONNECTED_032, UNCONNECTED_033, UNCONNECTED_034, 
		UNCONNECTED_035, UNCONNECTED_036, UNCONNECTED_037, 
		UNCONNECTED_038, UNCONNECTED_039, UNCONNECTED_040, 
		UNCONNECTED_041, instrc[105], instrc[104]}));
	AWDP_ADD_177 i_895(.O0(nbus_138), .opa({opa[31], opa[30], opa[29], opa[
		28], opa[27], opa[26], opa[25], opa[24], opa[23], opa[22], opa[
		21], opa[20], opa[19], opa[18], opa[17], opa[16], n_61034, opa[
		14], n_61025, n_61016, opa[11], opa[10], n_61007, opa[8], n_60998
		, n_60989, n_60980, opa[4], n_60971, n_60962, opa[1], n_60953}),
		 .I0({UNCONNECTED_042, UNCONNECTED_043, UNCONNECTED_044, 
		UNCONNECTED_045, UNCONNECTED_046, UNCONNECTED_047, 
		UNCONNECTED_048, UNCONNECTED_049, UNCONNECTED_050, 
		UNCONNECTED_051, UNCONNECTED_052, UNCONNECTED_053, n_58205, 
		UNCONNECTED_054, UNCONNECTED_055, UNCONNECTED_056, 
		UNCONNECTED_057, UNCONNECTED_058, UNCONNECTED_059, 
		UNCONNECTED_060, UNCONNECTED_061, UNCONNECTED_062, 
		UNCONNECTED_063, UNCONNECTED_064, UNCONNECTED_065, 
		UNCONNECTED_066, UNCONNECTED_067, UNCONNECTED_068, 
		UNCONNECTED_069, UNCONNECTED_070, instrc[105], instrc[104]}));
	AWDP_ADD_47 i_894(.O0(nbus_139), .opa({n_61034, opa[14], n_61025, n_61016
		, opa[11], opa[10], n_61007, opa[8], n_60998, n_60989, n_60980, opa
		[4], n_60971, n_60962, opa[1], n_60953}), .I0({UNCONNECTED_071, 
		UNCONNECTED_072, n_58202, UNCONNECTED_073, UNCONNECTED_074, 
		UNCONNECTED_075, UNCONNECTED_076, UNCONNECTED_077, 
		UNCONNECTED_078, UNCONNECTED_079, UNCONNECTED_080, 
		UNCONNECTED_081, UNCONNECTED_082, UNCONNECTED_083, instrc[105], instrc
		[104]}));
	AWDP_SUB_176 i_893(.O0(nbus_140), .opa({opa[31], opa[30], opa[29], opa[
		28], opa[27], opa[26], opa[25], opa[24], opa[23], opa[22], opa[
		21], opa[20], opa[19], opa[18], opa[17], opa[16], n_61034, opa[
		14], n_61025, n_61016, opa[11], opa[10], n_61007, opa[8], n_60998
		, n_60989, n_60980, opa[4], n_60971, n_60962, opa[1], n_60953}),
		 .I0({UNCONNECTED_084, UNCONNECTED_085, UNCONNECTED_086, 
		UNCONNECTED_087, UNCONNECTED_088, UNCONNECTED_089, 
		UNCONNECTED_090, UNCONNECTED_091, UNCONNECTED_092, 
		UNCONNECTED_093, UNCONNECTED_094, UNCONNECTED_095, n_58201, 
		UNCONNECTED_096, UNCONNECTED_097, UNCONNECTED_098, 
		UNCONNECTED_099, UNCONNECTED_100, UNCONNECTED_101, 
		UNCONNECTED_102, UNCONNECTED_103, UNCONNECTED_104, 
		UNCONNECTED_105, UNCONNECTED_106, UNCONNECTED_107, 
		UNCONNECTED_108, UNCONNECTED_109, UNCONNECTED_110, 
		UNCONNECTED_111, UNCONNECTED_112, instrc[105], instrc[104]}));
	AWDP_SUB_237 i_892(.O0(nbus_141), .opa({n_61034, opa[14], n_61025, n_61016
		, opa[11], opa[10], n_61007, opa[8], n_60998, n_60989, n_60980, opa
		[4], n_60971, n_60962, opa[1], n_60953}), .I0({UNCONNECTED_113, 
		UNCONNECTED_114, instrc[106], UNCONNECTED_115, UNCONNECTED_116, 
		UNCONNECTED_117, UNCONNECTED_118, UNCONNECTED_119, 
		UNCONNECTED_120, UNCONNECTED_121, UNCONNECTED_122, 
		UNCONNECTED_123, UNCONNECTED_124, UNCONNECTED_125, instrc[105], instrc
		[104]}));
	AWDP_ADD_198 i_891(.O0(nbus_142), .opd({n_58018, opd[30], n_57937, n_57946
		, n_57956, n_57965, opd[25], opd[24], opd[23], opd[22], opd[21],
		 opd[20], opd[19], opd[18], opd[17], opd[16], opd[15], opd[14], opd
		[13], opd[12], opd[11], opd[10], opd[9], opd[8], opd[7], opd[6],
		 opd[5], opd[4], opd[3], opd[2], opd[1], n_56964}), .I0({
		UNCONNECTED_126, UNCONNECTED_127, UNCONNECTED_128, 
		UNCONNECTED_129, UNCONNECTED_130, UNCONNECTED_131, 
		UNCONNECTED_132, UNCONNECTED_133, UNCONNECTED_134, 
		UNCONNECTED_135, UNCONNECTED_136, UNCONNECTED_137, 
		UNCONNECTED_138, UNCONNECTED_139, UNCONNECTED_140, 
		UNCONNECTED_141, UNCONNECTED_142, UNCONNECTED_143, 
		UNCONNECTED_144, UNCONNECTED_145, UNCONNECTED_146, 
		UNCONNECTED_147, UNCONNECTED_148, UNCONNECTED_149, 
		UNCONNECTED_150, UNCONNECTED_151, UNCONNECTED_152, n_58201, 
		UNCONNECTED_153, UNCONNECTED_154, instrc[105], instrc[104]}));
	AWDP_ADD_239 i_890(.O0(nbus_143), .opd({opd[15], opd[14], opd[13], opd[
		12], opd[11], opd[10], opd[9], opd[8], opd[7], opd[6], n_56982, n_56973
		, n_58783, n_58801, n_56955, n_56964}), .I0({UNCONNECTED_155, 
		UNCONNECTED_156, UNCONNECTED_157, UNCONNECTED_158, 
		UNCONNECTED_159, UNCONNECTED_160, UNCONNECTED_161, 
		UNCONNECTED_162, UNCONNECTED_163, UNCONNECTED_164, 
		UNCONNECTED_165, n_58205, UNCONNECTED_166, UNCONNECTED_167, instrc
		[105], instrc[104]}));
	AWDP_LSH_40 i_889(.O0(nbus_11291), .opb({opb[4], opb[3], opb[2], opb[1],
		 opb[0]}));
	AWDP_ADD_45 i_774(.O0({n_2701, n_2699, n_2697, n_2695, n_2693, n_2691, n_2689
		, n_2687, n_2685, n_2683, n_2681, n_2679, n_2677, n_2675, n_2673
		, n_2671, n_2669, n_2667, n_2665, n_2663, n_2661, n_2659, n_2657
		, n_2655, n_2653, n_2651, n_2649, n_2647, n_2645, n_2643, n_2641
		, n_2639}), .regs_6(regs_6), .opd({n_58018, opd[30], n_57937, n_57946
		, n_57956, n_57965, opd[25], opd[24], opd[23], opd[22], opd[21],
		 opd[20], opd[19], opd[18], opd[17], opd[16], opd[15], opd[14], opd
		[13], opd[12], opd[11], opd[10], opd[9], opd[8], opd[7], opd[6],
		 n_56982, n_56973, n_58783, opd[2], n_56955, n_56964}));
	AWDP_SUB_139 i_773(.O0({n_2702, n_2700, n_2698, n_2696, n_2694, n_2692, n_2690
		, n_2688, n_2686, n_2684, n_2682, n_2680, n_2678, n_2676, n_2674
		, n_2672, n_2670, n_2668, n_2666, n_2664, n_2662, n_2660, n_2658
		, n_2656, n_2654, n_2652, n_2650, n_2648, n_2646, n_2644, n_2642
		, n_2640}), .regs_6(regs_6), .opd({n_58018, opd[30], n_57937, n_57946
		, n_57956, n_57965, opd[25], opd[24], opd[23], opd[22], opd[21],
		 opd[20], opd[19], opd[18], opd[17], opd[16], opd[15], opd[14], opd
		[13], opd[12], opd[11], opd[10], opd[9], opd[8], opd[7], opd[6],
		 opd[5], opd[4], opd[3], opd[2], opd[1], n_56964}));
	AWDP_DEC_236 i_743(.O0({\regs_1_0[31] , \regs_1_0[30] , \regs_1_0[29] , \regs_1_0[28] 
		, \regs_1_0[27] , \regs_1_0[26] , \regs_1_0[25] , \regs_1_0[24] 
		, \regs_1_0[23] , \regs_1_0[22] , \regs_1_0[21] , \regs_1_0[20] 
		, \regs_1_0[19] , \regs_1_0[18] , \regs_1_0[17] , \regs_1_0[16] 
		, n_3487, n_3486, n_3485, n_3484, n_3483, n_3482, n_3481, n_3480
		, n_3479, n_3478, n_3477, n_3476, n_3475, n_3474, n_3473, n_3472
		}), .ecx(ecx));
	AWDP_DEC_206 i_742(.O0({\regs_1[15] , \regs_1[14] , \regs_1[13] , \regs_1[12] 
		, \regs_1[11] , \regs_1[10] , \regs_1[9] , \regs_1[8] , \regs_1[7] 
		, \regs_1[6] , \regs_1[5] , \regs_1[4] , \regs_1[3] , \regs_1[2] 
		, \regs_1[1] , \regs_1[0] }), .cx({ecx[15], ecx[14], ecx[13], ecx
		[12], ecx[11], ecx[10], ecx[9], ecx[8], ecx[7], ecx[6], ecx[5], ecx
		[4], ecx[3], ecx[2], ecx[1], ecx[0]}));
	AWDP_INC_125 i_738(.O0({n_3551, n_3550, n_3549, n_3548, n_3547, n_3546, n_3545
		, n_3544, n_3543, n_3542, n_3541, n_3540, n_3539, n_3538, n_3537
		, n_3536, n_3535, n_3534, n_3533, n_3532, n_3531, n_3530, n_3529
		, n_3528, n_3527, n_3526, n_3525, n_3524, n_3523, n_3522, n_3521
		, n_3520, n_3519, n_3518, n_3517, n_3516, n_3515, n_3514, n_3513
		, n_3512, n_3511, n_3510, n_3509, n_3508, n_3507, n_3506, n_3505
		, n_3504, n_3503, n_3502, n_3501, n_3500, n_3499, n_3498, n_3497
		, n_3496, n_3495, n_3494, n_3493, n_3492, n_3491, n_3490, n_3489
		, n_3488}), .I0({n_60591, n_60611, n_60620, n_60564, n_60573, n_60582
		, n_60510, n_60519, n_60528, n_60537, n_60546, n_60555, n_60483,
		 n_60492, n_60501, n_60474, nbus_11271[15], nbus_11271[14], nbus_11271
		[13], nbus_11271[12], nbus_11271[11], nbus_11271[10], nbus_11271
		[9], nbus_11271[8], nbus_11271[7], nbus_11271[6], nbus_11271[5],
		 nbus_11271[4], nbus_11271[3], nbus_11271[2], nbus_11271[1], nbus_11271
		[0], n_60458, n_58483, n_58474, n_58465, n_58456, n_58447, n_58438
		, n_58429, n_58420, n_58411, n_58402, n_58393, n_58384, n_58375,
		 n_58366, n_58357, n_58348, n_58339, n_58330, n_58321, n_58312, n_58303
		, n_58294, n_58285, n_58275, n_58265, nbus_11273[5], nbus_11273[
		4], n_58256, n_58247, n_58225, n_58238}));
	AWDP_INC_163 i_735(.O0({UNCONNECTED_168, UNCONNECTED_169, 
		UNCONNECTED_170, UNCONNECTED_171, UNCONNECTED_172, 
		UNCONNECTED_173, UNCONNECTED_174, UNCONNECTED_175, 
		UNCONNECTED_176, UNCONNECTED_177, UNCONNECTED_178, 
		UNCONNECTED_179, UNCONNECTED_180, UNCONNECTED_181, 
		UNCONNECTED_182, UNCONNECTED_183, UNCONNECTED_184, 
		UNCONNECTED_185, UNCONNECTED_186, UNCONNECTED_187, 
		UNCONNECTED_188, UNCONNECTED_189, UNCONNECTED_190, 
		UNCONNECTED_191, UNCONNECTED_192, UNCONNECTED_193, 
		UNCONNECTED_194, UNCONNECTED_195, UNCONNECTED_196, 
		UNCONNECTED_197, UNCONNECTED_198, n_3584, n_3583, n_3582, n_3581
		, n_3580, n_3579, n_3578, n_3577, n_3576, n_3575, n_3574, n_3573
		, n_3572, n_3571, n_3570, n_3569, n_3568, n_3567, n_3566, n_3565
		, n_3564, n_3563, n_3562, n_3561, n_3560, n_3559, n_3558, n_3557
		, n_3556, n_3555, n_3554, n_3553, n_3552}), .I0({UNCONNECTED_199
		, UNCONNECTED_200, UNCONNECTED_201, UNCONNECTED_202, 
		UNCONNECTED_203, UNCONNECTED_204, UNCONNECTED_205, 
		UNCONNECTED_206, UNCONNECTED_207, UNCONNECTED_208, 
		UNCONNECTED_209, UNCONNECTED_210, UNCONNECTED_211, 
		UNCONNECTED_212, UNCONNECTED_213, UNCONNECTED_214, 
		UNCONNECTED_215, UNCONNECTED_216, UNCONNECTED_217, 
		UNCONNECTED_218, UNCONNECTED_219, UNCONNECTED_220, 
		UNCONNECTED_221, UNCONNECTED_222, UNCONNECTED_223, 
		UNCONNECTED_224, UNCONNECTED_225, UNCONNECTED_226, 
		UNCONNECTED_227, UNCONNECTED_228, UNCONNECTED_229, 
		UNCONNECTED_230, n_58983, n_58992, n_58947, n_58929, n_58938, n_58911
		, n_58920, n_58893, n_58902, n_58875, n_58884, n_58857, n_58866,
		 n_59077, n_59086, n_59059, n_59068, n_59041, n_58965, n_59050, n_58974
		, n_59023, n_59032, n_59014, \nbus_11290[7] , \nbus_11290[6] , \nbus_11290[5] 
		, \nbus_11290[4] , \nbus_11290[3] , \nbus_11290[2] , n_59001, n_58956
		}));
	AWDP_LE_211 i_734(.O0({n_577}), .divq(divq), .I0({UNCONNECTED_231, divr[
		63], divr[62], divr[61], divr[60], divr[59], divr[58], divr[57],
		 divr[56], divr[55], divr[54], divr[53], divr[52], divr[51], divr
		[50], divr[49], divr[48], divr[47], divr[46], divr[45], divr[44]
		, divr[43], divr[42], divr[41], divr[40], divr[39], divr[38], divr
		[37], divr[36], divr[35], divr[34], divr[33], divr[32], divr[31]
		, divr[30], divr[29], divr[28], divr[27], divr[26], divr[25], divr
		[24], divr[23], divr[22], divr[21], divr[20], divr[19], divr[18]
		, divr[17], divr[16], divr[15], divr[14], divr[13], divr[12], divr
		[11], divr[10], divr[9], divr[8], divr[7], divr[6], divr[5], divr
		[4], divr[3], divr[2], divr[1]}));
	AWDP_SUB_39 i_731(.O0(divr_1), .divr(divr), .divq(divq));
	AWDP_GE_13 i_729(.O0({n_579}), .divr(divr), .divq(divq));
	AWDP_LSH_10 i_728(.O0(nbus_11346), .opd({opd[5], opd[4], opd[3], opd[2],
		 opd[1], opd[0]}));
	AWDP_ADD_11 i_727(.O0(opc_14), .opc({n_60600, opc[30], opc[29], opc[28],
		 opc[27], opc[26], opc[25], opc[24], opc[23], opc[22], opc[21], opc
		[20], opc[19], opc[18], opc[17], opc[16], opc[15], opc[14], opc[
		13], opc[12], opc[11], opc[10], opc[9], opc[8], opc[7], opc[6], opc
		[5], opc[4], opc[3], opc[2], opc[1], n_60467}), .I0(nbus_11346)
		);
	AWDP_INC_210 i_721(.O0({n_3680, n_3679, n_3678, n_3677, n_3676, n_3675, n_3674
		, n_3673, n_3672, n_3671, n_3670, n_3669, n_3668, n_3667, n_3666
		, n_3665, n_3664, n_3663, n_3662, n_3661, n_3660, n_3659, n_3658
		, n_3657, n_3656, n_3655, n_3654, n_3653, n_3652, n_3651, n_3650
		, n_3649}), .I0(nbus_11270));
	AWDP_DEC_7 i_718(.O0({\opc_1[7] , \opc_1[6] , \opc_1[5] , \opc_1[4] , \opc_1[3] 
		, \opc_1[2] , \opc_1[1] , \opc_1[0] }), .opc({opc[7], opc[6], opc
		[5], opc[4], opc[3], opc[2], opc[1], n_60467}));
	AWDP_DEC_143 i_715(.O0({\opc_5[31] , \opc_5[30] , \opc_5[29] , \opc_5[28] 
		, \opc_5[27] , \opc_5[26] , \opc_5[25] , \opc_5[24] , \opc_5[23] 
		, \opc_5[22] , \opc_5[21] , \opc_5[20] , \opc_5[19] , \opc_5[18] 
		, \opc_5[17] , \opc_5[16] , \opc_5[15] , \opc_5[14] , \opc_5[13] 
		, \opc_5[12] , \opc_5[11] , \opc_5[10] , \opc_5[9] , \opc_5[8] ,
		 \opc_5[7] , \opc_5[6] , \opc_5[5] , n_3686, n_3685, n_3684, n_3683
		, n_3682}), .opc({n_60600, opc[30], opc[29], opc[28], opc[27], opc
		[26], opc[25], opc[24], opc[23], opc[22], opc[21], opc[20], opc[
		19], opc[18], opc[17], opc[16], opc[15], opc[14], opc[13], opc[
		12], opc[11], opc[10], opc[9], opc[8], opc[7], opc[6], opc[5], opc
		[4], opc[3], opc[2], opc[1], n_60467}));
	AWDP_EQ_138 i_710(.O0({n_585}), .I0({n_60629, opb[30], opb[29], opb[28],
		 opb[27], opb[26], opb[25], opb[24], opb[23], opb[22], opb[21], opb
		[20], opb[19], opb[18], opb[17], opb[16], opb[15], opb[14], opb[
		13], opb[12], opb[11], opb[10], opb[9], opb[8], opb[7], opb[6], opb
		[5], opb[4], opb[3], opb[2], opb[1], opb[0], n_60600, opc[30], opc
		[29], opc[28], opc[27], opc[26], opc[25], opc[24], opc[23], opc[
		22], opc[21], opc[20], opc[19], opc[18], opc[17], opc[16], opc[
		15], opc[14], opc[13], opc[12], opc[11], opc[10], opc[9], opc[8]
		, opc[7], opc[6], opc[5], opc[4], opc[3], opc[2], opc[1], n_60467
		}), .I1({regs_2[31], regs_2[30], regs_2[29], regs_2[28], regs_2[
		27], regs_2[26], regs_2[25], regs_2[24], regs_2[23], regs_2[22],
		 regs_2[21], regs_2[20], regs_2[19], regs_2[18], regs_2[17], regs_2
		[16], regs_2[15], regs_2[14], regs_2[13], regs_2[12], regs_2[11]
		, regs_2[10], regs_2[9], regs_2[8], regs_2[7], regs_2[6], regs_2
		[5], regs_2[4], regs_2[3], regs_2[2], regs_2[1], regs_2[0], regs_0
		[31], regs_0[30], regs_0[29], regs_0[28], regs_0[27], regs_0[26]
		, regs_0[25], regs_0[24], regs_0[23], regs_0[22], regs_0[21], regs_0
		[20], regs_0[19], regs_0[18], regs_0[17], regs_0[16], regs_0[15]
		, regs_0[14], regs_0[13], regs_0[12], regs_0[11], regs_0[10], regs_0
		[9], regs_0[8], regs_0[7], regs_0[6], regs_0[5], regs_0[4], regs_0
		[3], regs_0[2], regs_0[1], regs_0[0]}));
	AWDP_INC_153 i_702(.O0(opa_0), .I0({n_60458, n_58483, n_58474, n_58465, n_58456
		, n_58447, n_58438, n_58429, n_58420, n_58411, n_58402, n_58393,
		 n_58384, n_58375, n_58366, n_58357, n_58348, n_58339, n_58330, n_58321
		, n_58312, n_58303, n_58294, n_58285, n_58275, n_58265, nbus_11273
		[5], nbus_11273[4], n_58256, n_58247, n_58225, n_58238}));
	AWDP_INC_26111934 i_700(.O0({\opa_1[15] , \opa_1[14] , \opa_1[13] , \opa_1[12] 
		, \opa_1[11] , \opa_1[10] , \opa_1[9] , \opa_1[8] , \opa_1[7] , \opa_1[6] 
		, \opa_1[5] , \opa_1[4] , \opa_1[3] , \opa_1[2] , \opa_1[1] , \opa_1[0] 
		}), .I0({n_58348, n_58339, n_58330, n_58321, n_58312, n_58303, n_58294
		, n_58285, n_58275, n_58265, nbus_11273[5], nbus_11273[4], n_58256
		, n_58247, n_58225, n_58238}));
	AWDP_INC_200 i_689(.O0({n_6290, n_6289, n_6288, n_6287, n_6286, n_6285, n_6284
		, n_6283, n_6282, n_6281, n_6280, n_6279, n_6278, n_6277, n_6276
		, n_6275, n_6274, n_6273, n_6272, n_6271, n_6270, n_6269, n_6268
		, n_6267, n_6266, n_6265, n_6264, n_6263, n_6262, n_6261, n_6260
		, n_6259}), .I0({n_60591, n_60611, n_60620, n_60564, n_60573, n_60582
		, n_60510, n_60519, n_60528, n_60537, n_60546, n_60555, n_60483,
		 n_60492, n_60501, n_60474, nbus_11271[15], nbus_11271[14], nbus_11271
		[13], nbus_11271[12], nbus_11271[11], nbus_11271[10], nbus_11271
		[9], nbus_11271[8], nbus_11271[7], nbus_11271[6], nbus_11271[5],
		 nbus_11271[4], nbus_11271[3], nbus_11271[2], nbus_11271[1], nbus_11271
		[0]}));
	arithbox arithbox(.arithop({\opcode[3] , \opcode[2] , \opcode[1] , \opcode[0] 
		}), .calc_sz(calc_sz), .ci(\eflags[0] ), .co(nCF_arithbox), .af(nAF_arithbox
		), .ai(\eflags[4] ), .sa(opas_arithbox), .sb(opbs_arithbox), .opa
		({opa[31], opa[30], opa[29], opa[28], opa[27], opa[26], opa[25],
		 opa[24], opa[23], opa[22], opa[21], opa[20], opa[19], opa[18], opa
		[17], opa[16], n_61034, opa[14], n_61025, n_61016, opa[11], opa[
		10], n_61007, opa[8], n_60998, n_60989, n_60980, opa[4], n_60971
		, n_60962, opa[1], n_60953}), .opb({n_60629, opb[30], opb[29], opb
		[28], opb[27], opb[26], opb[25], opb[24], opb[23], opb[22], opb[
		21], opb[20], opb[19], opb[18], opb[17], opb[16], opb[15], opb[
		14], opb[13], opb[12], opb[11], opb[10], opb[9], opb[8], opb[7],
		 opb[6], opb[5], opb[4], opb[3], opb[2], opb[1], opb[0]}), .resa
		(resa_arithbox), .cmp(tcmp_arithbox));
	synthetic_op synthetic_op(.clk(clk), .sel({\opcode[2] , \opcode[1] , \opcode[0] 
		}), .opa32({opa[31], opa[30], opa[29], opa[28], opa[27], opa[26]
		, opa[25], opa[24], opa[23], opa[22], opa[21], opa[20], opa[19],
		 opa[18], opa[17], opa[16], n_61034, opa[14], n_61025, n_61016, opa
		[11], opa[10], n_61007, opa[8], n_60998, n_60989, n_60980, opa[4
		], n_60971, n_60962, opa[1], n_60953}), .opb32({n_60629, opb[30]
		, opb[29], opb[28], opb[27], opb[26], opb[25], opb[24], opb[23],
		 opb[22], opb[21], opb[20], opb[19], opb[18], opb[17], opb[16], opb
		[15], opb[14], opb[13], opb[12], opb[11], opb[10], opb[9], opb[8
		], opb[7], opb[6], opb[5], opb[4], opb[3], opb[2], opb[1], opb[0
		]}), .res64(mul64));
	AWDP_ADD_242 i_654(.O0({n_4727, n_4722, n_4717, n_4712, n_4707, n_4702, n_4697
		, n_4692, n_4687, n_4682, n_4677, n_4672, n_4667, n_4662, n_4657
		, n_4652, n_4647, n_4642, n_4637, n_4632, n_4627, n_4622, n_4617
		, n_4612, n_4607, n_4602, n_4597, n_4592, n_4587, n_4582, n_4577
		, n_4572}), .opb({n_60629, opb[30], opb[29], opb[28], opb[27], opb
		[26], opb[25], opb[24], opb[23], opb[22], opb[21], opb[20], opb[
		19], opb[18], opb[17], opb[16], opb[15], opb[14], opb[13], opb[
		12], opb[11], opb[10], opb[9], opb[8], opb[7], opb[6], opb[5], opb
		[4], opb[3], opb[2], opb[1], opb[0]}), .I0({UNCONNECTED_232, 
		UNCONNECTED_233, UNCONNECTED_234, UNCONNECTED_235, 
		UNCONNECTED_236, UNCONNECTED_237, UNCONNECTED_238, 
		UNCONNECTED_239, UNCONNECTED_240, UNCONNECTED_241, 
		UNCONNECTED_242, UNCONNECTED_243, UNCONNECTED_244, 
		UNCONNECTED_245, UNCONNECTED_246, UNCONNECTED_247, 
		UNCONNECTED_248, UNCONNECTED_249, UNCONNECTED_250, 
		UNCONNECTED_251, UNCONNECTED_252, UNCONNECTED_253, 
		UNCONNECTED_254, UNCONNECTED_255, n_60998, n_60989, n_60980, opa
		[4], n_60971, n_60962, opa[1], n_60953}));
	AWDP_ADD_107 i_652(.O0({n_4729, n_4723, n_4718, n_4713, n_4708, n_4703, n_4698
		, n_4693, n_4688, n_4683, n_4678, n_4673, n_4668, n_4663, n_4658
		, n_4653, n_4648, n_4643, n_4638, n_4633, n_4628, n_4623, n_4618
		, n_4613, n_4608, n_4603, n_4598, n_4593, n_4588, n_4583, n_4578
		, n_4573}), .opd({n_58018, opd[30], n_57937, n_57946, n_57956, n_57965
		, opd[25], opd[24], opd[23], opd[22], opd[21], opd[20], opd[19],
		 opd[18], opd[17], opd[16], opd[15], opd[14], opd[13], opd[12], opd
		[11], opd[10], opd[9], opd[8], opd[7], opd[6], n_56982, n_56973,
		 n_58783, n_58801, n_56955, n_56964}), .I0({UNCONNECTED_256, 
		UNCONNECTED_257, UNCONNECTED_258, n_60600, opc[30], opc[29], opc
		[28], opc[27], opc[26], opc[25], opc[24], opc[23], opc[22], opc[
		21], opc[20], opc[19], opc[18], opc[17], opc[16], opc[15], opc[
		14], opc[13], opc[12], opc[11], opc[10], opc[9], opc[8], opc[7],
		 opc[6], opc[5], UNCONNECTED_259, UNCONNECTED_260}));
	AWDP_ADD_189 i_651(.O0({n_4730, n_4724, n_4719, n_4714, n_4709, n_4704, n_4699
		, n_4694, n_4689, n_4684, n_4679, n_4674, n_4669, n_4664, n_4659
		, n_4654, n_4649, n_4644, n_4639, n_4634, n_4629, n_4624, n_4619
		, n_4614, n_4609, n_4604, n_4599, n_4594, n_4589, n_4584, n_4579
		, n_4574}), .opd({n_58018, opd[30], n_57937, n_57946, n_57956, n_57965
		, opd[25], opd[24], opd[23], opd[22], opd[21], opd[20], opd[19],
		 opd[18], opd[17], opd[16], opd[15], opd[14], opd[13], opd[12], opd
		[11], opd[10], opd[9], opd[8], opd[7], opd[6], n_56982, n_56973,
		 n_58783, n_58801, n_56955, n_56964}));
	AWDP_ADD_201 i_617(.O0({n_847, n_845, n_843, n_841, n_839, n_837, n_835,
		 n_833, n_831, n_829, n_827, n_825, n_823, n_821, n_819, n_817, n_815
		, n_813, n_811, n_809, n_807, n_805, n_803, n_801, n_799, n_797,
		 n_795, n_793, n_791, n_789, n_787, n_785}), .ldtr(ldtr), .I0({gs
		[31], gs[30], gs[29], gs[28], gs[27], gs[26], gs[25], gs[24], gs
		[23], gs[22], gs[21], gs[20], gs[19], gs[18], gs[17], gs[16], gs
		[15], gs[14], gs[13], gs[12], gs[11], gs[10], gs[9], gs[8], gs[7
		], gs[6], gs[5], gs[4], gs[3], UNCONNECTED_261, UNCONNECTED_262,
		 UNCONNECTED_263}));
	AWDP_ADD_216 i_615(.O0({n_848, n_846, n_844, n_842, n_840, n_838, n_836,
		 n_834, n_832, n_830, n_828, n_826, n_824, n_822, n_820, n_818, n_816
		, n_814, n_812, n_810, n_808, n_806, n_804, n_802, n_800, n_798,
		 n_796, n_794, n_792, n_790, n_788, n_786}), .gdtr(gdtr), .I0({gs
		[31], gs[30], gs[29], gs[28], gs[27], gs[26], gs[25], gs[24], gs
		[23], gs[22], gs[21], gs[20], gs[19], gs[18], gs[17], gs[16], gs
		[15], gs[14], gs[13], gs[12], gs[11], gs[10], gs[9], gs[8], gs[7
		], gs[6], gs[5], gs[4], gs[3], UNCONNECTED_264, UNCONNECTED_265,
		 UNCONNECTED_266}));
	AWDP_ADD_117 i_612(.O0({n_6675, n_6673, n_6671, n_6669, n_6667, n_6665, n_6663
		, n_6661, n_6659, n_6657, n_6655, n_6653, n_6651, n_6649, n_6647
		, n_6645, n_6643, n_6641, n_6639, n_6637, n_6635, n_6633, n_6631
		, n_6629, n_6627, n_6625, n_6623, n_6621, n_6619, n_6617, n_6615
		, n_6613}), .idtr(idtr), .I0({instrc[95], instrc[94], instrc[93]
		, instrc[92], instrc[91], instrc[90], instrc[89], instrc[88], instrc
		[87], instrc[86], instrc[85], instrc[84], instrc[83], instrc[82]
		, instrc[81], instrc[80], UNCONNECTED_267, UNCONNECTED_268, 
		UNCONNECTED_269}));
	AWDP_ADD_135 i_610(.O0({n_6676, n_6674, n_6672, n_6670, n_6668, n_6666, n_6664
		, n_6662, n_6660, n_6658, n_6656, n_6654, n_6652, n_6650, n_6648
		, n_6646, n_6644, n_6642, n_6640, n_6638, n_6636, n_6634, n_6632
		, n_6630, n_6628, n_6626, n_6624, n_6622, n_6620, n_6618, n_6616
		, n_6614}), .gdtr(gdtr), .I0({\tr[15] , \tr[14] , \tr[13] , \tr[12] 
		, \tr[11] , \tr[10] , \tr[9] , \tr[8] , \tr[7] , \tr[6] , \tr[5] 
		, \tr[4] , \tr[3] , UNCONNECTED_270, UNCONNECTED_271, 
		UNCONNECTED_272}));
	AWDP_SUB_192 i_609(.O0(Daddrs_8), .opd({n_58018, opd[30], n_57937, n_57946
		, n_57956, n_57965, opd[25], opd[24], opd[23], opd[22], opd[21],
		 opd[20], opd[19], opd[18], opd[17], opd[16], opd[15], opd[14], opd
		[13], opd[12], opd[11], opd[10], opd[9], opd[8], opd[7], opd[6],
		 n_56982, n_56973, n_58783, n_58801, n_56955, n_56964}));
	AWDP_ADD_84 i_608(.O0(Daddrs_1), .Daddrs(Daddr));
	AWDP_ADD_74 i_607(.O0(Daddrs_3), .Daddrs(Daddr));
	AWDP_ADD_20 i_605(.O0({n_5311, n_5310, n_5309, n_5308, n_5307, n_5306, n_5305
		, n_5304, n_5303, n_5302, n_5301, n_5300, n_5299, n_5298, n_5297
		, n_5296, n_5295, n_5294, n_5293, n_5292, n_5291, n_5290, n_5289
		, n_5288, n_5287, n_5286, n_5285, n_5284, n_5283, n_5282, n_5281
		, n_5280}), .opd({n_58018, opd[30], n_57937, n_57946, n_57956, n_57965
		, opd[25], opd[24], opd[23], opd[22], opd[21], opd[20], opd[19],
		 opd[18], opd[17], opd[16], opd[15], opd[14], opd[13], opd[12], opd
		[11], opd[10], opd[9], opd[8], opd[7], opd[6], opd[5], opd[4], opd
		[3], opd[2], opd[1], opd[0]}), .desc(desc));
	AWDP_ADD_190 i_571(.O0({n_1442, n_1441, n_1440, n_1439, n_1438, n_1437, n_1436
		, n_1435, n_1434, n_1433, n_1432, n_1431, n_1430, n_1429, n_1428
		, n_1427, n_1426, n_1425, n_1424, n_1423, n_1422, n_1421, n_1420
		, n_1419, n_1418, n_1417, n_1416, n_1415, n_1414, n_1413, n_1412
		, n_1411}), .I0({UNCONNECTED_273, UNCONNECTED_274, 
		UNCONNECTED_275, UNCONNECTED_276, UNCONNECTED_277, 
		UNCONNECTED_278, UNCONNECTED_279, UNCONNECTED_280, 
		UNCONNECTED_281, UNCONNECTED_282, UNCONNECTED_283, 
		UNCONNECTED_284, UNCONNECTED_285, UNCONNECTED_286, 
		UNCONNECTED_287, UNCONNECTED_288, regs_14[15], regs_14[14], regs_14
		[13], regs_14[12], regs_14[11], regs_14[10], regs_14[9], regs_14
		[8], regs_14[7], regs_14[6], regs_14[5], regs_14[4], regs_14[3],
		 regs_14[2], regs_14[1], regs_14[0]}), .I1({\nbus_14543[27] , \nbus_14543[26] 
		, \nbus_14543[25] , \nbus_14543[24] , \nbus_14543[23] , \nbus_14543[22] 
		, \nbus_14543[21] , \nbus_14543[20] , \nbus_14543[19] , \nbus_14543[18] 
		, \nbus_14543[17] , \nbus_14543[16] , \nbus_14543[15] , \nbus_14543[14] 
		, \nbus_14543[13] , \nbus_14543[12] , \nbus_14543[11] , \nbus_14543[10] 
		, \nbus_14543[9] , \nbus_14543[8] , \nbus_14543[7] , \nbus_14543[6] 
		, \nbus_14543[5] , \nbus_14543[4] , \nbus_14543[3] , \nbus_14543[2] 
		, cs[1], cs[0], UNCONNECTED_289, UNCONNECTED_290, 
		UNCONNECTED_291, UNCONNECTED_292}));
endmodule
module cpu(clk, rstn, iack, int_cpu, ivect, cr0, cr2, icr2, cr3, cs, pg_fault, ipg_fault
		, useq_ptr, valid_len, queue, pg_en, pc_out, pc_req, read_req, write_req
		, read_ack, write_ack, flush_Itlb, flush_Dtlb, readio_req, writeio_req
		, readio_ack, writeio_ack, write_data, writeio_data, read_data, readio_data
		, write_sz, read_sz, io_add, Daddr, pt_fault, wr_fault);

	input clk;
	input rstn;
	output iack;
	input int_cpu;
	input [7:0] ivect;
	output [31:0] cr0;
	input [31:0] cr2;
	input [31:0] icr2;
	output [31:0] cr3;
	output [31:0] cs;
	input pg_fault;
	input ipg_fault;
	output [3:0] useq_ptr;
	input [5:0] valid_len;
	input [127:0] queue;
	output pg_en;
	output [31:0] pc_out;
	output pc_req;
	output read_req;
	output write_req;
	input read_ack;
	input write_ack;
	output flush_Itlb;
	output flush_Dtlb;
	output readio_req;
	output writeio_req;
	input readio_ack;
	input writeio_ack;
	output [31:0] write_data;
	output [31:0] writeio_data;
	input [31:0] read_data;
	input [31:0] readio_data;
	output [1:0] write_sz;
	output [1:0] read_sz;
	output [31:0] io_add;
	output [31:0] Daddr;
	input pt_fault;
	input wr_fault;

	wire [2:0] reps;
	wire [2:0] opz;
	wire [127:0] dec2vliw;
	wire [31:0] lenpc;
	wire [31:0] add_src;
	wire [7:0] from_acu;
	wire [63:0] to_acu;
	wire [210:0] deco2acu;



	vliw i_vliw(.clk(clk), .rstn(rstn), .instrc(dec2vliw), .ie(ie), .readio_data
		(readio_data), .io_add({UNCONNECTED_000, UNCONNECTED_001, 
		UNCONNECTED_002, UNCONNECTED_003, UNCONNECTED_004, 
		UNCONNECTED_005, UNCONNECTED_006, UNCONNECTED_007, 
		UNCONNECTED_008, UNCONNECTED_009, UNCONNECTED_010, 
		UNCONNECTED_011, UNCONNECTED_012, UNCONNECTED_013, 
		UNCONNECTED_014, UNCONNECTED_015, io_add[15], io_add[14], io_add
		[13], io_add[12], io_add[11], io_add[10], io_add[9], io_add[8], io_add
		[7], io_add[6], io_add[5], io_add[4], io_add[3], io_add[2], io_add
		[1], io_add[0]}), .writeio_data(writeio_data), .writeio_req(writeio_req
		), .readio_req(readio_req), .writeio_ack(writeio_ack), .readio_ack
		(readio_ack), .read_reqs(read_req), .read_ack(read_ack), .read_data
		(read_data), .over_seg({\over_seg[5] , UNCONNECTED_016, 
		UNCONNECTED_017, UNCONNECTED_018, UNCONNECTED_019, 
		UNCONNECTED_020}), .cr3({cr3[31], cr3[30], cr3[29], cr3[28], cr3
		[27], cr3[26], cr3[25], cr3[24], cr3[23], cr3[22], cr3[21], cr3[
		20], cr3[19], cr3[18], cr3[17], cr3[16], cr3[15], cr3[14], cr3[
		13], cr3[12], UNCONNECTED_021, UNCONNECTED_022, UNCONNECTED_023,
		 UNCONNECTED_024, UNCONNECTED_025, UNCONNECTED_026, 
		UNCONNECTED_027, UNCONNECTED_028, UNCONNECTED_029, 
		UNCONNECTED_030, UNCONNECTED_031, UNCONNECTED_032}), .cr2(cr2), 
		.icr2(icr2), .cr0({UNCONNECTED_033, UNCONNECTED_034, 
		UNCONNECTED_035, UNCONNECTED_036, UNCONNECTED_037, 
		UNCONNECTED_038, UNCONNECTED_039, UNCONNECTED_040, 
		UNCONNECTED_041, UNCONNECTED_042, UNCONNECTED_043, 
		UNCONNECTED_044, UNCONNECTED_045, UNCONNECTED_046, 
		UNCONNECTED_047, cr0[16], UNCONNECTED_048, UNCONNECTED_049, 
		UNCONNECTED_050, UNCONNECTED_051, UNCONNECTED_052, 
		UNCONNECTED_053, UNCONNECTED_054, UNCONNECTED_055, 
		UNCONNECTED_056, UNCONNECTED_057, UNCONNECTED_058, 
		UNCONNECTED_059, UNCONNECTED_060, \cr0[2] , UNCONNECTED_061, \cr0[0] 
		}), .write_reqs(write_req), .write_ack(write_ack), .write_data(write_data
		), .Daddr(Daddr), .write_sz(write_sz), .cs({UNCONNECTED_062, 
		UNCONNECTED_063, UNCONNECTED_064, UNCONNECTED_065, 
		UNCONNECTED_066, UNCONNECTED_067, UNCONNECTED_068, 
		UNCONNECTED_069, UNCONNECTED_070, UNCONNECTED_071, 
		UNCONNECTED_072, UNCONNECTED_073, UNCONNECTED_074, 
		UNCONNECTED_075, UNCONNECTED_076, UNCONNECTED_077, 
		UNCONNECTED_078, UNCONNECTED_079, UNCONNECTED_080, 
		UNCONNECTED_081, UNCONNECTED_082, UNCONNECTED_083, 
		UNCONNECTED_084, UNCONNECTED_085, UNCONNECTED_086, 
		UNCONNECTED_087, UNCONNECTED_088, UNCONNECTED_089, 
		UNCONNECTED_090, UNCONNECTED_091, cs[1], cs[0]}), .add_src(add_src
		), .from_acu(from_acu), .to_acu(to_acu), .pg_en(pg_en), .imm({
		UNCONNECTED_092, UNCONNECTED_093, UNCONNECTED_094, 
		UNCONNECTED_095, UNCONNECTED_096, UNCONNECTED_097, 
		UNCONNECTED_098, UNCONNECTED_099, UNCONNECTED_100, 
		UNCONNECTED_101, UNCONNECTED_102, UNCONNECTED_103, 
		UNCONNECTED_104, UNCONNECTED_105, UNCONNECTED_106, 
		UNCONNECTED_107, \imm[47] , \imm[46] , \imm[45] , \imm[44] , \imm[43] 
		, \imm[42] , \imm[41] , \imm[40] , \imm[39] , \imm[38] , \imm[37] 
		, \imm[36] , \imm[35] , \imm[34] , \imm[33] , \imm[32] , \imm[31] 
		, \imm[30] , \imm[29] , \imm[28] , \imm[27] , \imm[26] , \imm[25] 
		, \imm[24] , \imm[23] , \imm[22] , \imm[21] , \imm[20] , \imm[19] 
		, \imm[18] , \imm[17] , \imm[16] , \imm[15] , \imm[14] , \imm[13] 
		, \imm[12] , \imm[11] , \imm[10] , \imm[9] , \imm[8] , \imm[7] ,
		 \imm[6] , \imm[5] , \imm[4] , \imm[3] , \imm[2] , \imm[1] , \imm[0] 
		}), .lenpc(lenpc), .pc_out(pc_out), .pc_req(pc_req), .opz(opz), 
		.reps(reps), .flush_tlb(flush_Itlb), .flush_Dtlb(flush_Dtlb), .terminate
		(term), .start_up(st), .pg_fault(pg_fault), .ipg_fault(ipg_fault
		), .wr_fault(wr_fault), .pt_fault(pt_fault));
	acu i_acu(.clk(clk), .rstn(rstn), .from_regf(to_acu), .add_src(add_src),
		 .to_regf(from_acu), .from_dec(deco2acu), .db67(\cr0[0] ));
	deco i_deco(.clk(clk), .rstn(rstn), .useq_ptr(useq_ptr), .in128(queue), 
		.adz(\cr0[0] ), .pc_req(pc_req), .ivect(ivect), .int_main(int_cpu
		), .iack(iack), .ie(ie), .pg_fault(pg_fault), .ipg_fault(ipg_fault
		), .cpl({cs[1], cs[0]}), .cr0({UNCONNECTED_108, UNCONNECTED_109,
		 UNCONNECTED_110, UNCONNECTED_111, UNCONNECTED_112, 
		UNCONNECTED_113, UNCONNECTED_114, UNCONNECTED_115, 
		UNCONNECTED_116, UNCONNECTED_117, UNCONNECTED_118, 
		UNCONNECTED_119, UNCONNECTED_120, UNCONNECTED_121, 
		UNCONNECTED_122, UNCONNECTED_123, UNCONNECTED_124, 
		UNCONNECTED_125, UNCONNECTED_126, UNCONNECTED_127, 
		UNCONNECTED_128, UNCONNECTED_129, UNCONNECTED_130, 
		UNCONNECTED_131, UNCONNECTED_132, UNCONNECTED_133, 
		UNCONNECTED_134, UNCONNECTED_135, UNCONNECTED_136, \cr0[2] , 
		UNCONNECTED_137, UNCONNECTED_138}), .valid_len(valid_len), .to_vliw
		(dec2vliw), .lenpc_out(lenpc), .immediate({UNCONNECTED_139, 
		UNCONNECTED_140, UNCONNECTED_141, UNCONNECTED_142, 
		UNCONNECTED_143, UNCONNECTED_144, UNCONNECTED_145, 
		UNCONNECTED_146, UNCONNECTED_147, UNCONNECTED_148, 
		UNCONNECTED_149, UNCONNECTED_150, UNCONNECTED_151, 
		UNCONNECTED_152, UNCONNECTED_153, UNCONNECTED_154, \imm[47] , \imm[46] 
		, \imm[45] , \imm[44] , \imm[43] , \imm[42] , \imm[41] , \imm[40] 
		, \imm[39] , \imm[38] , \imm[37] , \imm[36] , \imm[35] , \imm[34] 
		, \imm[33] , \imm[32] , \imm[31] , \imm[30] , \imm[29] , \imm[28] 
		, \imm[27] , \imm[26] , \imm[25] , \imm[24] , \imm[23] , \imm[22] 
		, \imm[21] , \imm[20] , \imm[19] , \imm[18] , \imm[17] , \imm[16] 
		, \imm[15] , \imm[14] , \imm[13] , \imm[12] , \imm[11] , \imm[10] 
		, \imm[9] , \imm[8] , \imm[7] , \imm[6] , \imm[5] , \imm[4] , \imm[3] 
		, \imm[2] , \imm[1] , \imm[0] }), .to_acu(deco2acu), .operand_size
		(opz), .reps(reps), .over_seg({\over_seg[5] , UNCONNECTED_155, 
		UNCONNECTED_156, UNCONNECTED_157, UNCONNECTED_158, 
		UNCONNECTED_159}), .term(term), .start(st));
endmodule
module AWDP_ADD_27(O0, addrshft, useq_ptr);
    output [6:0] O0;
    input [5:0] addrshft;
    input [3:0] useq_ptr;
    // Line 58
    wire [6:0] O0;
    // Line 81
    wire [6:0] N861;

    // Line 58
    assign O0 = N861;
    // Line 81
    assign N861 = useq_ptr + addrshft;
endmodule

module AWDP_ADD_9(O0, addr);

	output [31:0] O0;
	input [31:0] addr;

	wire \addr[4] ;
	wire \addr[5] ;
	wire \addr[6] ;
	wire \addr[7] ;
	wire \addr[8] ;
	wire \addr[9] ;
	wire \addr[10] ;
	wire \addr[11] ;
	wire \addr[12] ;
	wire \addr[13] ;
	wire \addr[14] ;
	wire \addr[15] ;
	wire \addr[16] ;
	wire \addr[17] ;
	wire \addr[18] ;
	wire \addr[19] ;
	wire \addr[20] ;
	wire \addr[21] ;
	wire \addr[22] ;
	wire \addr[23] ;
	wire \addr[24] ;
	wire \addr[25] ;
	wire \addr[26] ;
	wire \addr[27] ;
	wire \addr[28] ;
	wire \addr[29] ;
	wire \addr[30] ;
	wire \addr[31] ;


	assign O0[0] = addr[0];
	assign O0[1] = addr[1];
	assign O0[2] = addr[2];
	assign O0[3] = addr[3];
	assign \addr[4]  = addr[4];
	assign \addr[5]  = addr[5];
	assign \addr[6]  = addr[6];
	assign \addr[7]  = addr[7];
	assign \addr[8]  = addr[8];
	assign \addr[9]  = addr[9];
	assign \addr[10]  = addr[10];
	assign \addr[11]  = addr[11];
	assign \addr[12]  = addr[12];
	assign \addr[13]  = addr[13];
	assign \addr[14]  = addr[14];
	assign \addr[15]  = addr[15];
	assign \addr[16]  = addr[16];
	assign \addr[17]  = addr[17];
	assign \addr[18]  = addr[18];
	assign \addr[19]  = addr[19];
	assign \addr[20]  = addr[20];
	assign \addr[21]  = addr[21];
	assign \addr[22]  = addr[22];
	assign \addr[23]  = addr[23];
	assign \addr[24]  = addr[24];
	assign \addr[25]  = addr[25];
	assign \addr[26]  = addr[26];
	assign \addr[27]  = addr[27];
	assign \addr[28]  = addr[28];
	assign \addr[29]  = addr[29];
	assign \addr[30]  = addr[30];
	assign \addr[31]  = addr[31];

	notech_ha2 i_27(.A(\addr[31] ), .B(n_300), .Z(O0[31]));
	notech_ha2 i_26(.A(\addr[30] ), .B(n_298), .Z(O0[30]), .CO(n_300));
	notech_ha2 i_25(.A(\addr[29] ), .B(n_296), .Z(O0[29]), .CO(n_298));
	notech_ha2 i_24(.A(\addr[28] ), .B(n_294), .Z(O0[28]), .CO(n_296));
	notech_ha2 i_23(.A(\addr[27] ), .B(n_292), .Z(O0[27]), .CO(n_294));
	notech_ha2 i_22(.A(\addr[26] ), .B(n_290), .Z(O0[26]), .CO(n_292));
	notech_ha2 i_21(.A(\addr[25] ), .B(n_288), .Z(O0[25]), .CO(n_290));
	notech_ha2 i_20(.A(\addr[24] ), .B(n_286), .Z(O0[24]), .CO(n_288));
	notech_ha2 i_19(.A(\addr[23] ), .B(n_284), .Z(O0[23]), .CO(n_286));
	notech_ha2 i_18(.A(\addr[22] ), .B(n_282), .Z(O0[22]), .CO(n_284));
	notech_ha2 i_17(.A(\addr[21] ), .B(n_280), .Z(O0[21]), .CO(n_282));
	notech_ha2 i_16(.A(\addr[20] ), .B(n_278), .Z(O0[20]), .CO(n_280));
	notech_ha2 i_15(.A(\addr[19] ), .B(n_276), .Z(O0[19]), .CO(n_278));
	notech_ha2 i_14(.A(\addr[18] ), .B(n_274), .Z(O0[18]), .CO(n_276));
	notech_ha2 i_13(.A(\addr[17] ), .B(n_272), .Z(O0[17]), .CO(n_274));
	notech_ha2 i_12(.A(\addr[16] ), .B(n_270), .Z(O0[16]), .CO(n_272));
	notech_ha2 i_11(.A(\addr[15] ), .B(n_268), .Z(O0[15]), .CO(n_270));
	notech_ha2 i_10(.A(\addr[14] ), .B(n_266), .Z(O0[14]), .CO(n_268));
	notech_ha2 i_9(.A(\addr[13] ), .B(n_264), .Z(O0[13]), .CO(n_266));
	notech_ha2 i_8(.A(\addr[12] ), .B(n_262), .Z(O0[12]), .CO(n_264));
	notech_ha2 i_7(.A(\addr[11] ), .B(n_260), .Z(O0[11]), .CO(n_262));
	notech_ha2 i_6(.A(\addr[10] ), .B(n_258), .Z(O0[10]), .CO(n_260));
	notech_ha2 i_5(.A(\addr[9] ), .B(n_256), .Z(O0[9]), .CO(n_258));
	notech_ha2 i_4(.A(\addr[8] ), .B(n_254), .Z(O0[8]), .CO(n_256));
	notech_ha2 i_3(.A(\addr[7] ), .B(n_252), .Z(O0[7]), .CO(n_254));
	notech_ha2 i_2(.A(\addr[6] ), .B(n_250), .Z(O0[6]), .CO(n_252));
	notech_ha2 i_1(.A(\addr[5] ), .B(\addr[4] ), .Z(O0[5]), .CO(n_250));
	notech_inv i_0(.A(\addr[4] ), .Z(O0[4]));
endmodule
module AWDP_EQ_228374(O0, tagA, addr);
    output [0:0] O0;
    input [17:0] tagA;
    input [31:14] addr;
    // Line 128
    wire [0:0] N875;
    // Line 128
    wire [0:0] O0;

    // Line 128
    assign N875 = tagA == addr;
    // Line 128
    assign O0 = N875;
endmodule

module AWDP_EQ_328640(O0, addr, addrf);
    output [0:0] O0;
    input [31:0] addr;
    input [31:0] addrf;
    // Line 58
    wire [0:0] O0;
    // Line 85
    wire [0:0] N886;

    // Line 58
    assign O0 = N886;
    // Line 85
    assign N886 = addr == addrf;
endmodule

module AWDP_INC_10(O0, purge_cnt);

	output [10:0] O0;
	input [10:0] purge_cnt;




	notech_ha2 i_10(.A(purge_cnt[10]), .B(n_106), .Z(O0[10]));
	notech_ha2 i_9(.A(purge_cnt[9]), .B(n_104), .Z(O0[9]), .CO(n_106));
	notech_ha2 i_8(.A(purge_cnt[8]), .B(n_102), .Z(O0[8]), .CO(n_104));
	notech_ha2 i_7(.A(purge_cnt[7]), .B(n_100), .Z(O0[7]), .CO(n_102));
	notech_ha2 i_6(.A(purge_cnt[6]), .B(n_98), .Z(O0[6]), .CO(n_100));
	notech_ha2 i_5(.A(purge_cnt[5]), .B(n_96), .Z(O0[5]), .CO(n_98));
	notech_ha2 i_4(.A(purge_cnt[4]), .B(n_94), .Z(O0[4]), .CO(n_96));
	notech_ha2 i_3(.A(purge_cnt[3]), .B(n_92), .Z(O0[3]), .CO(n_94));
	notech_ha2 i_2(.A(purge_cnt[2]), .B(n_90), .Z(O0[2]), .CO(n_92));
	notech_ha2 i_1(.A(purge_cnt[1]), .B(purge_cnt[0]), .Z(O0[1]), .CO(n_90)
		);
	notech_inv i_0(.A(purge_cnt[0]), .Z(O0[0]));
endmodule
module useq(iaddr, idata, code_req, code_ack, clk, rstn, useq_ptr, squeue, pc_in
		, pc_req, cs, pg_en, pg_fault, pc_pg_fault, valid_len, busy_ram
		);

	output [31:0] iaddr;
	input [127:0] idata;
	output code_req;
	input code_ack;
	input clk;
	input rstn;
	input [3:0] useq_ptr;
	output [127:0] squeue;
	input [31:0] pc_in;
	input pc_req;
	input [31:0] cs;
	input pg_en;
	input pg_fault;
	output pc_pg_fault;
	output [5:0] valid_len;
	input busy_ram;

	wire [1:0] wptr;
	wire [255:0] queue;
	wire [1:0] fault_wptr;
	wire [3:0] tagV;
	wire [17:0] tagA;
	wire [31:0] addr_0;
	wire [9:0] cacheA;
	wire [149:0] cacheD;
	wire [6:0] nbus_12105;
	wire [31:0] addrf;
	wire [5:0] addrshft;
	wire [10:0] purge_cnt;

	supply0 AMBIT_GND;
	supply1 AMBIT_VDD;


	notech_inv i_15646(.A(n_63813), .Z(n_63814));
	notech_inv i_15645(.A(n_63808), .Z(n_63813));
	notech_inv i_15644(.A(n_63811), .Z(n_63812));
	notech_inv i_15643(.A(n_63804), .Z(n_63811));
	notech_inv i_15642(.A(n_63809), .Z(n_63810));
	notech_inv i_15641(.A(n_63802), .Z(n_63809));
	notech_inv i_15640(.A(n_63807), .Z(n_63808));
	notech_inv i_15639(.A(n_63810), .Z(n_63807));
	notech_inv i_15638(.A(n_63805), .Z(n_63806));
	notech_inv i_15637(.A(cacheD[148]), .Z(n_63805));
	notech_inv i_15636(.A(n_63803), .Z(n_63804));
	notech_inv i_15635(.A(n_63806), .Z(n_63803));
	notech_inv i_15634(.A(n_63801), .Z(n_63802));
	notech_inv i_15633(.A(n_63812), .Z(n_63801));
	notech_inv i_15510(.A(n_63677), .Z(n_63678));
	notech_inv i_15509(.A(n_63628), .Z(n_63677));
	notech_inv i_15468(.A(n_63635), .Z(n_63636));
	notech_inv i_15467(.A(n_63560), .Z(n_63635));
	notech_inv i_15466(.A(n_63633), .Z(n_63634));
	notech_inv i_15465(.A(n_63554), .Z(n_63633));
	notech_inv i_15464(.A(n_63631), .Z(n_63632));
	notech_inv i_15463(.A(n_63550), .Z(n_63631));
	notech_inv i_15462(.A(n_63629), .Z(n_63630));
	notech_inv i_15461(.A(n_63548), .Z(n_63629));
	notech_inv i_15460(.A(n_63627), .Z(n_63628));
	notech_inv i_15459(.A(n_63630), .Z(n_63627));
	notech_inv i_15396(.A(n_63563), .Z(n_63564));
	notech_inv i_15395(.A(n_63488), .Z(n_63563));
	notech_inv i_15394(.A(n_63561), .Z(n_63562));
	notech_inv i_15393(.A(n_63486), .Z(n_63561));
	notech_inv i_15392(.A(n_63559), .Z(n_63560));
	notech_inv i_15391(.A(n_63562), .Z(n_63559));
	notech_inv i_15390(.A(n_63557), .Z(n_63558));
	notech_inv i_15389(.A(n_63482), .Z(n_63557));
	notech_inv i_15388(.A(n_63555), .Z(n_63556));
	notech_inv i_15387(.A(n_63480), .Z(n_63555));
	notech_inv i_15386(.A(n_63553), .Z(n_63554));
	notech_inv i_15385(.A(n_63556), .Z(n_63553));
	notech_inv i_15384(.A(n_63551), .Z(n_63552));
	notech_inv i_15383(.A(n_63478), .Z(n_63551));
	notech_inv i_15382(.A(n_63549), .Z(n_63550));
	notech_inv i_15381(.A(n_63552), .Z(n_63549));
	notech_inv i_15380(.A(n_63547), .Z(n_63548));
	notech_inv i_15379(.A(n_63632), .Z(n_63547));
	notech_inv i_15322(.A(n_63489), .Z(n_63490));
	notech_inv i_15321(.A(clk), .Z(n_63489));
	notech_inv i_15320(.A(n_63487), .Z(n_63488));
	notech_inv i_15319(.A(n_63490), .Z(n_63487));
	notech_inv i_15318(.A(n_63485), .Z(n_63486));
	notech_inv i_15317(.A(n_63564), .Z(n_63485));
	notech_inv i_15316(.A(n_63483), .Z(n_63484));
	notech_inv i_15315(.A(n_63396), .Z(n_63483));
	notech_inv i_15314(.A(n_63481), .Z(n_63482));
	notech_inv i_15313(.A(n_63484), .Z(n_63481));
	notech_inv i_15312(.A(n_63479), .Z(n_63480));
	notech_inv i_15311(.A(n_63558), .Z(n_63479));
	notech_inv i_15310(.A(n_63477), .Z(n_63478));
	notech_inv i_15309(.A(n_63634), .Z(n_63477));
	notech_inv i_15228(.A(n_63395), .Z(n_63396));
	notech_inv i_15227(.A(n_63636), .Z(n_63395));
	notech_inv i_14702(.A(n_62839), .Z(n_62861));
	notech_inv i_14700(.A(n_62839), .Z(n_62859));
	notech_inv i_14699(.A(n_62839), .Z(n_62858));
	notech_inv i_14695(.A(n_62839), .Z(n_62854));
	notech_inv i_14693(.A(n_62839), .Z(n_62852));
	notech_inv i_14690(.A(n_62839), .Z(n_62849));
	notech_inv i_14688(.A(n_62839), .Z(n_62847));
	notech_inv i_14687(.A(n_62839), .Z(n_62846));
	notech_inv i_14682(.A(n_62839), .Z(n_62841));
	notech_inv i_14681(.A(n_62839), .Z(code_req));
	notech_inv i_14680(.A(n_62863), .Z(n_62839));
	notech_inv i_14561(.A(n_62686), .Z(n_62709));
	notech_inv i_14560(.A(n_62686), .Z(n_62708));
	notech_inv i_14559(.A(n_62686), .Z(n_62707));
	notech_inv i_14558(.A(n_62686), .Z(n_62706));
	notech_inv i_14557(.A(n_62686), .Z(n_62705));
	notech_inv i_14555(.A(n_62686), .Z(n_62703));
	notech_inv i_14554(.A(n_62686), .Z(n_62702));
	notech_inv i_14553(.A(n_62686), .Z(n_62701));
	notech_inv i_14552(.A(n_62686), .Z(n_62700));
	notech_inv i_14551(.A(n_62686), .Z(n_62699));
	notech_inv i_14549(.A(n_62686), .Z(n_62697));
	notech_inv i_14548(.A(n_62686), .Z(n_62696));
	notech_inv i_14547(.A(n_62686), .Z(n_62695));
	notech_inv i_14546(.A(n_62686), .Z(n_62694));
	notech_inv i_14545(.A(n_62686), .Z(n_62693));
	notech_inv i_14543(.A(n_62686), .Z(n_62691));
	notech_inv i_14542(.A(n_62686), .Z(n_62690));
	notech_inv i_14541(.A(n_62686), .Z(n_62689));
	notech_inv i_14540(.A(n_62686), .Z(n_62688));
	notech_inv i_14539(.A(n_62686), .Z(n_62687));
	notech_inv i_14538(.A(rstn), .Z(n_62686));
	notech_inv i_14537(.A(n_62680), .Z(n_62685));
	notech_inv i_14536(.A(n_62680), .Z(n_62684));
	notech_inv i_14535(.A(n_62680), .Z(n_62683));
	notech_inv i_14534(.A(n_62680), .Z(n_62682));
	notech_inv i_14533(.A(n_62680), .Z(n_62681));
	notech_inv i_14532(.A(rstn), .Z(n_62680));
	notech_inv i_13403(.A(n_61558), .Z(n_61567));
	notech_inv i_13399(.A(n_61558), .Z(n_61563));
	notech_inv i_13395(.A(n_61558), .Z(n_61559));
	notech_inv i_13394(.A(pc_req), .Z(n_61558));
	notech_inv i_13368(.A(n_61436), .Z(n_61438));
	notech_inv i_13367(.A(n_61436), .Z(pc_pg_fault));
	notech_inv i_13366(.A(n_61444), .Z(n_61436));
	notech_inv i_13364(.A(n_61417), .Z(n_61433));
	notech_inv i_13362(.A(n_61417), .Z(n_61431));
	notech_inv i_13361(.A(n_61417), .Z(n_61430));
	notech_inv i_13357(.A(n_61417), .Z(n_61426));
	notech_inv i_13355(.A(n_61417), .Z(n_61424));
	notech_inv i_13352(.A(n_61417), .Z(n_61421));
	notech_inv i_13350(.A(n_61417), .Z(n_61419));
	notech_inv i_13349(.A(n_61417), .Z(n_61418));
	notech_inv i_13348(.A(wptr[1]), .Z(n_61417));
	notech_inv i_13341(.A(n_61404), .Z(n_61409));
	notech_inv i_13337(.A(n_61404), .Z(n_61405));
	notech_inv i_13336(.A(n_3086), .Z(n_61404));
	notech_inv i_13334(.A(n_61385), .Z(n_61401));
	notech_inv i_13332(.A(n_61385), .Z(n_61399));
	notech_inv i_13331(.A(n_61385), .Z(n_61398));
	notech_inv i_13327(.A(n_61385), .Z(n_61394));
	notech_inv i_13325(.A(n_61385), .Z(n_61392));
	notech_inv i_13323(.A(n_61385), .Z(n_61390));
	notech_inv i_13321(.A(n_61385), .Z(n_61388));
	notech_inv i_13319(.A(n_61385), .Z(n_61386));
	notech_inv i_13318(.A(n_14258715), .Z(n_61385));
	notech_inv i_13311(.A(n_61376), .Z(n_61377));
	notech_inv i_13310(.A(n_14228712), .Z(n_61376));
	notech_inv i_13306(.A(n_61376), .Z(n_61372));
	notech_inv i_13302(.A(n_61376), .Z(n_61368));
	notech_inv i_13297(.A(n_61376), .Z(n_61363));
	notech_inv i_13293(.A(n_61376), .Z(n_61359));
	notech_inv i_13283(.A(n_61348), .Z(n_61349));
	notech_inv i_13282(.A(n_61329), .Z(n_61348));
	notech_inv i_13278(.A(n_61348), .Z(n_61344));
	notech_inv i_13274(.A(n_61348), .Z(n_61340));
	notech_inv i_13269(.A(n_61348), .Z(n_61335));
	notech_inv i_13265(.A(n_61348), .Z(n_61331));
	notech_inv i_13263(.A(n_61376), .Z(n_61329));
	notech_inv i_13255(.A(n_61320), .Z(n_61321));
	notech_inv i_13254(.A(n_61301), .Z(n_61320));
	notech_inv i_13250(.A(n_61320), .Z(n_61316));
	notech_inv i_13246(.A(n_61320), .Z(n_61312));
	notech_inv i_13241(.A(n_61320), .Z(n_61307));
	notech_inv i_13237(.A(n_61320), .Z(n_61303));
	notech_inv i_13235(.A(n_61376), .Z(n_61301));
	notech_inv i_13225(.A(n_61289), .Z(n_61290));
	notech_inv i_13224(.A(\nbus_12122[0] ), .Z(n_61289));
	notech_inv i_13105(.A(n_61390), .Z(n_61160));
	notech_inv i_13103(.A(n_61390), .Z(n_61158));
	notech_inv i_13102(.A(n_61390), .Z(n_61157));
	notech_inv i_13098(.A(n_61390), .Z(n_61153));
	notech_inv i_13096(.A(n_61390), .Z(n_61151));
	notech_inv i_13093(.A(n_61390), .Z(n_61148));
	notech_inv i_13091(.A(n_61390), .Z(n_61146));
	notech_inv i_13090(.A(n_61390), .Z(n_61145));
	notech_inv i_12071(.A(n_60096), .Z(n_60101));
	notech_inv i_12067(.A(n_60096), .Z(n_60097));
	notech_inv i_12066(.A(n_3082), .Z(n_60096));
	notech_inv i_12064(.A(n_60080), .Z(n_60093));
	notech_inv i_12062(.A(n_60080), .Z(n_60091));
	notech_inv i_12058(.A(n_60080), .Z(n_60087));
	notech_inv i_12052(.A(n_60080), .Z(n_60081));
	notech_inv i_12051(.A(n_1304), .Z(n_60080));
	notech_inv i_12049(.A(n_60064), .Z(n_60077));
	notech_inv i_12047(.A(n_60064), .Z(n_60075));
	notech_inv i_12043(.A(n_60064), .Z(n_60071));
	notech_inv i_12037(.A(n_60064), .Z(n_60065));
	notech_inv i_12036(.A(n_1305), .Z(n_60064));
	notech_inv i_12034(.A(n_60048), .Z(n_60061));
	notech_inv i_12032(.A(n_60048), .Z(n_60059));
	notech_inv i_12028(.A(n_60048), .Z(n_60055));
	notech_inv i_12022(.A(n_60048), .Z(n_60049));
	notech_inv i_12021(.A(n_1296), .Z(n_60048));
	notech_inv i_12019(.A(n_60032), .Z(n_60045));
	notech_inv i_12017(.A(n_60032), .Z(n_60043));
	notech_inv i_12013(.A(n_60032), .Z(n_60039));
	notech_inv i_12007(.A(n_60032), .Z(n_60033));
	notech_inv i_12006(.A(n_1297), .Z(n_60032));
	notech_inv i_12004(.A(n_60016), .Z(n_60029));
	notech_inv i_12002(.A(n_60016), .Z(n_60027));
	notech_inv i_11998(.A(n_60016), .Z(n_60023));
	notech_inv i_11992(.A(n_60016), .Z(n_60017));
	notech_inv i_11991(.A(n_1300), .Z(n_60016));
	notech_inv i_11989(.A(n_60000), .Z(n_60013));
	notech_inv i_11987(.A(n_60000), .Z(n_60011));
	notech_inv i_11983(.A(n_60000), .Z(n_60007));
	notech_inv i_11977(.A(n_60000), .Z(n_60001));
	notech_inv i_11976(.A(n_1301), .Z(n_60000));
	notech_inv i_11973(.A(n_59981), .Z(n_59996));
	notech_inv i_11971(.A(n_59981), .Z(n_59994));
	notech_inv i_11966(.A(n_59981), .Z(n_59989));
	notech_inv i_11965(.A(n_59981), .Z(n_59988));
	notech_inv i_11959(.A(n_59981), .Z(n_59982));
	notech_inv i_11958(.A(n_1290), .Z(n_59981));
	notech_inv i_11956(.A(n_59962), .Z(n_59978));
	notech_inv i_11954(.A(n_59962), .Z(n_59976));
	notech_inv i_11953(.A(n_59962), .Z(n_59975));
	notech_inv i_11949(.A(n_59962), .Z(n_59971));
	notech_inv i_11947(.A(n_59962), .Z(n_59969));
	notech_inv i_11944(.A(n_59962), .Z(n_59966));
	notech_inv i_11942(.A(n_59962), .Z(n_59964));
	notech_inv i_11941(.A(n_59962), .Z(n_59963));
	notech_inv i_11940(.A(n_1291), .Z(n_59962));
	notech_inv i_11938(.A(n_59943), .Z(n_59959));
	notech_inv i_11936(.A(n_59943), .Z(n_59957));
	notech_inv i_11935(.A(n_59943), .Z(n_59956));
	notech_inv i_11931(.A(n_59943), .Z(n_59952));
	notech_inv i_11929(.A(n_59943), .Z(n_59950));
	notech_inv i_11926(.A(n_59943), .Z(n_59947));
	notech_inv i_11924(.A(n_59943), .Z(n_59945));
	notech_inv i_11923(.A(n_59943), .Z(n_59944));
	notech_inv i_11922(.A(n_1292), .Z(n_59943));
	notech_inv i_11920(.A(n_59924), .Z(n_59940));
	notech_inv i_11918(.A(n_59924), .Z(n_59938));
	notech_inv i_11917(.A(n_59924), .Z(n_59937));
	notech_inv i_11913(.A(n_59924), .Z(n_59933));
	notech_inv i_11911(.A(n_59924), .Z(n_59931));
	notech_inv i_11908(.A(n_59924), .Z(n_59928));
	notech_inv i_11906(.A(n_59924), .Z(n_59926));
	notech_inv i_11905(.A(n_59924), .Z(n_59925));
	notech_inv i_11904(.A(n_1989), .Z(n_59924));
	notech_inv i_11897(.A(n_59911), .Z(n_59916));
	notech_inv i_11893(.A(n_59911), .Z(n_59912));
	notech_inv i_11892(.A(n_2006), .Z(n_59911));
	notech_inv i_11885(.A(n_59898), .Z(n_59903));
	notech_inv i_11881(.A(n_59898), .Z(n_59899));
	notech_inv i_11880(.A(n_2005), .Z(n_59898));
	notech_inv i_11873(.A(n_59885), .Z(n_59890));
	notech_inv i_11869(.A(n_59885), .Z(n_59886));
	notech_inv i_11868(.A(n_2003), .Z(n_59885));
	notech_inv i_11861(.A(n_59872), .Z(n_59877));
	notech_inv i_11857(.A(n_59872), .Z(n_59873));
	notech_inv i_11856(.A(n_2002), .Z(n_59872));
	notech_inv i_11849(.A(n_59859), .Z(n_59864));
	notech_inv i_11845(.A(n_59859), .Z(n_59860));
	notech_inv i_11844(.A(n_1986), .Z(n_59859));
	notech_inv i_11837(.A(n_59846), .Z(n_59851));
	notech_inv i_11833(.A(n_59846), .Z(n_59847));
	notech_inv i_11832(.A(n_1985), .Z(n_59846));
	notech_inv i_11825(.A(n_59833), .Z(n_59838));
	notech_inv i_11821(.A(n_59833), .Z(n_59834));
	notech_inv i_11820(.A(n_1991), .Z(n_59833));
	notech_inv i_11813(.A(n_59820), .Z(n_59825));
	notech_inv i_11809(.A(n_59820), .Z(n_59821));
	notech_inv i_11808(.A(n_1990), .Z(n_59820));
	notech_inv i_11801(.A(n_59807), .Z(n_59812));
	notech_inv i_11797(.A(n_59807), .Z(n_59808));
	notech_inv i_11796(.A(n_1998), .Z(n_59807));
	notech_inv i_11789(.A(n_59794), .Z(n_59799));
	notech_inv i_11785(.A(n_59794), .Z(n_59795));
	notech_inv i_11784(.A(n_1997), .Z(n_59794));
	notech_inv i_11777(.A(n_59781), .Z(n_59786));
	notech_inv i_11773(.A(n_59781), .Z(n_59782));
	notech_inv i_11772(.A(n_1995), .Z(n_59781));
	notech_inv i_11765(.A(n_59768), .Z(n_59773));
	notech_inv i_11761(.A(n_59768), .Z(n_59769));
	notech_inv i_11760(.A(n_1994), .Z(n_59768));
	notech_inv i_11758(.A(n_59752), .Z(n_59765));
	notech_inv i_11756(.A(n_59752), .Z(n_59763));
	notech_inv i_11752(.A(n_59752), .Z(n_59759));
	notech_inv i_11746(.A(n_59752), .Z(n_59753));
	notech_inv i_11745(.A(n_1318), .Z(n_59752));
	notech_inv i_11743(.A(n_59736), .Z(n_59749));
	notech_inv i_11741(.A(n_59736), .Z(n_59747));
	notech_inv i_11737(.A(n_59736), .Z(n_59743));
	notech_inv i_11731(.A(n_59736), .Z(n_59737));
	notech_inv i_11730(.A(n_1321), .Z(n_59736));
	notech_inv i_11728(.A(n_59720), .Z(n_59733));
	notech_inv i_11726(.A(n_59720), .Z(n_59731));
	notech_inv i_11722(.A(n_59720), .Z(n_59727));
	notech_inv i_11716(.A(n_59720), .Z(n_59721));
	notech_inv i_11715(.A(n_1310), .Z(n_59720));
	notech_inv i_11713(.A(n_59704), .Z(n_59717));
	notech_inv i_11711(.A(n_59704), .Z(n_59715));
	notech_inv i_11707(.A(n_59704), .Z(n_59711));
	notech_inv i_11701(.A(n_59704), .Z(n_59705));
	notech_inv i_11700(.A(n_1311), .Z(n_59704));
	notech_inv i_11698(.A(n_59688), .Z(n_59701));
	notech_inv i_11696(.A(n_59688), .Z(n_59699));
	notech_inv i_11692(.A(n_59688), .Z(n_59695));
	notech_inv i_11686(.A(n_59688), .Z(n_59689));
	notech_inv i_11685(.A(n_1314), .Z(n_59688));
	notech_inv i_11683(.A(n_59672), .Z(n_59685));
	notech_inv i_11681(.A(n_59672), .Z(n_59683));
	notech_inv i_11677(.A(n_59672), .Z(n_59679));
	notech_inv i_11671(.A(n_59672), .Z(n_59673));
	notech_inv i_11670(.A(n_1315), .Z(n_59672));
	notech_inv i_11668(.A(n_59651), .Z(n_59669));
	notech_inv i_11666(.A(n_59651), .Z(n_59667));
	notech_inv i_11663(.A(n_59651), .Z(n_59664));
	notech_inv i_11661(.A(n_59651), .Z(n_59662));
	notech_inv i_11658(.A(n_59651), .Z(n_59659));
	notech_inv i_11656(.A(n_59651), .Z(n_59657));
	notech_inv i_11653(.A(n_59651), .Z(n_59654));
	notech_inv i_11651(.A(n_59651), .Z(n_59652));
	notech_inv i_11650(.A(n_3081), .Z(n_59651));
	notech_inv i_8797(.A(\nbus_12119[0] ), .Z(n_56608));
	notech_inv i_8795(.A(\nbus_12119[0] ), .Z(n_56606));
	notech_inv i_8792(.A(\nbus_12119[0] ), .Z(n_56603));
	notech_inv i_8790(.A(\nbus_12119[0] ), .Z(n_56601));
	notech_inv i_8787(.A(\nbus_12119[0] ), .Z(n_56598));
	notech_inv i_8785(.A(\nbus_12119[0] ), .Z(n_56596));
	notech_inv i_8782(.A(\nbus_12119[0] ), .Z(n_56593));
	notech_inv i_8780(.A(\nbus_12119[0] ), .Z(n_56591));
	notech_inv i_8777(.A(\nbus_12119[128] ), .Z(n_56587));
	notech_inv i_8775(.A(\nbus_12119[128] ), .Z(n_56585));
	notech_inv i_8772(.A(\nbus_12119[128] ), .Z(n_56582));
	notech_inv i_8770(.A(\nbus_12119[128] ), .Z(n_56580));
	notech_inv i_8767(.A(\nbus_12119[128] ), .Z(n_56577));
	notech_inv i_8765(.A(\nbus_12119[128] ), .Z(n_56575));
	notech_inv i_8762(.A(\nbus_12119[128] ), .Z(n_56572));
	notech_inv i_8760(.A(\nbus_12119[128] ), .Z(n_56570));
	notech_inv i_8757(.A(n_56548), .Z(n_56566));
	notech_inv i_8755(.A(n_56548), .Z(n_56564));
	notech_inv i_8752(.A(n_56548), .Z(n_56561));
	notech_inv i_8750(.A(n_56548), .Z(n_56559));
	notech_inv i_8747(.A(n_56548), .Z(n_56556));
	notech_inv i_8745(.A(n_56548), .Z(n_56554));
	notech_inv i_8742(.A(n_56548), .Z(n_56551));
	notech_inv i_8740(.A(n_56548), .Z(n_56549));
	notech_inv i_8739(.A(n_309759578), .Z(n_56548));
	notech_ao4 i_129033640(.A(n_1991), .B(n_17414), .C(n_1990), .D(n_17475),
		 .Z(n_2546));
	notech_and4 i_129333637(.A(n_2542), .B(n_2544), .C(n_2546), .D(n_1785), 
		.Z(n_2547));
	notech_ao4 i_128433646(.A(n_1995), .B(n_17382), .C(n_1994), .D(n_17398),
		 .Z(n_2548));
	notech_ao4 i_128533645(.A(n_1998), .B(n_17406), .C(n_1997), .D(n_17390),
		 .Z(n_2549));
	notech_and3 i_129133639(.A(n_2549), .B(n_2548), .C(n_1798), .Z(n_2551)
		);
	notech_ao4 i_128833642(.A(n_2003), .B(n_17427), .C(n_2002), .D(n_17491),
		 .Z(n_2552));
	notech_ao4 i_128933641(.A(n_2006), .B(n_17459), .C(n_2005), .D(n_17443),
		 .Z(n_2553));
	notech_ao4 i_131233618(.A(n_59975), .B(n_17351), .C(n_59956), .D(n_17359
		), .Z(n_2556));
	notech_ao4 i_131433616(.A(n_1986), .B(n_17367), .C(n_1985), .D(n_17375),
		 .Z(n_2558));
	notech_ao4 i_132133609(.A(n_1991), .B(n_17415), .C(n_1990), .D(n_17477),
		 .Z(n_2560));
	notech_and4 i_132433606(.A(n_2556), .B(n_2558), .C(n_2560), .D(n_1801), 
		.Z(n_2561));
	notech_ao4 i_131533615(.A(n_1995), .B(n_17383), .C(n_1994), .D(n_17399),
		 .Z(n_2562));
	notech_ao4 i_131633614(.A(n_1998), .B(n_17407), .C(n_1997), .D(n_17391),
		 .Z(n_2563));
	notech_and3 i_132233608(.A(n_2563), .B(n_2562), .C(n_1814), .Z(n_2565)
		);
	notech_ao4 i_131933611(.A(n_2003), .B(n_17429), .C(n_2002), .D(n_17493),
		 .Z(n_2566));
	notech_ao4 i_132033610(.A(n_2006), .B(n_17461), .C(n_2005), .D(n_17445),
		 .Z(n_2567));
	notech_ao4 i_134333587(.A(n_59975), .B(n_17352), .C(n_59956), .D(n_17360
		), .Z(n_2570));
	notech_ao4 i_134533585(.A(n_1986), .B(n_17368), .C(n_1985), .D(n_17376),
		 .Z(n_2572));
	notech_ao4 i_135233578(.A(n_59838), .B(n_17416), .C(n_59825), .D(n_17479
		), .Z(n_2574));
	notech_and4 i_135533575(.A(n_2570), .B(n_2572), .C(n_2574), .D(n_1817), 
		.Z(n_2575));
	notech_ao4 i_134633584(.A(n_59786), .B(n_17384), .C(n_59773), .D(n_17400
		), .Z(n_2576));
	notech_ao4 i_134733583(.A(n_59812), .B(n_17408), .C(n_59799), .D(n_17392
		), .Z(n_2577));
	notech_and3 i_135333577(.A(n_2577), .B(n_2576), .C(n_1830), .Z(n_2579)
		);
	notech_ao4 i_135033580(.A(n_59890), .B(n_17431), .C(n_59877), .D(n_17495
		), .Z(n_2580));
	notech_ao4 i_135133579(.A(n_59916), .B(n_17463), .C(n_59903), .D(n_17447
		), .Z(n_2581));
	notech_ao4 i_137433556(.A(n_59975), .B(n_17353), .C(n_59956), .D(n_17361
		), .Z(n_2584));
	notech_ao4 i_137633554(.A(n_59864), .B(n_17369), .C(n_59851), .D(n_17377
		), .Z(n_2586));
	notech_ao4 i_138333547(.A(n_1991), .B(n_17417), .C(n_1990), .D(n_17481),
		 .Z(n_2588));
	notech_and4 i_138633544(.A(n_2584), .B(n_2586), .C(n_2588), .D(n_1833), 
		.Z(n_2589));
	notech_ao4 i_137733553(.A(n_1995), .B(n_17385), .C(n_1994), .D(n_17401),
		 .Z(n_2590));
	notech_ao4 i_137833552(.A(n_1998), .B(n_17409), .C(n_1997), .D(n_17393),
		 .Z(n_2591));
	notech_and3 i_138433546(.A(n_2591), .B(n_2590), .C(n_1846), .Z(n_2593)
		);
	notech_ao4 i_138133549(.A(n_2003), .B(n_17433), .C(n_2002), .D(n_17497),
		 .Z(n_2594));
	notech_ao4 i_138233548(.A(n_2006), .B(n_17465), .C(n_2005), .D(n_17449),
		 .Z(n_2595));
	notech_ao4 i_140533525(.A(n_59975), .B(n_17354), .C(n_59956), .D(n_17362
		), .Z(n_2598));
	notech_ao4 i_140733523(.A(n_1986), .B(n_17370), .C(n_1985), .D(n_17378),
		 .Z(n_2600));
	notech_ao4 i_141433516(.A(n_1991), .B(n_17418), .C(n_1990), .D(n_17483),
		 .Z(n_2602));
	notech_and4 i_141733513(.A(n_2598), .B(n_2600), .C(n_2602), .D(n_1849), 
		.Z(n_2603));
	notech_ao4 i_140833522(.A(n_1995), .B(n_17386), .C(n_1994), .D(n_17402),
		 .Z(n_2604));
	notech_ao4 i_140933521(.A(n_1998), .B(n_17410), .C(n_1997), .D(n_17394),
		 .Z(n_2605));
	notech_and3 i_141533515(.A(n_2605), .B(n_2604), .C(n_1862), .Z(n_2607)
		);
	notech_ao4 i_141233518(.A(n_2003), .B(n_17435), .C(n_2002), .D(n_17499),
		 .Z(n_2608));
	notech_ao4 i_141333517(.A(n_2006), .B(n_17467), .C(n_2005), .D(n_17451),
		 .Z(n_2609));
	notech_ao4 i_143633494(.A(n_59956), .B(n_17363), .C(n_59994), .D(n_17347
		), .Z(n_2612));
	notech_ao4 i_143833492(.A(n_1986), .B(n_17371), .C(n_1985), .D(n_17379),
		 .Z(n_2614));
	notech_ao4 i_144533485(.A(n_1991), .B(n_17421), .C(n_1990), .D(n_17485),
		 .Z(n_2616));
	notech_and4 i_144833482(.A(n_2612), .B(n_2614), .C(n_2616), .D(n_1865), 
		.Z(n_2617));
	notech_ao4 i_143933491(.A(n_1995), .B(n_17387), .C(n_1994), .D(n_17403),
		 .Z(n_2618));
	notech_ao4 i_144033490(.A(n_1998), .B(n_17411), .C(n_1997), .D(n_17395),
		 .Z(n_2619));
	notech_and3 i_144633484(.A(n_2619), .B(n_2618), .C(n_1878), .Z(n_2621)
		);
	notech_ao4 i_144333487(.A(n_2003), .B(n_17437), .C(n_2002), .D(n_17501),
		 .Z(n_2622));
	notech_ao4 i_144433486(.A(n_2006), .B(n_17469), .C(n_2005), .D(n_17453),
		 .Z(n_2623));
	notech_ao4 i_146733463(.A(n_59975), .B(n_17356), .C(n_59956), .D(n_17364
		), .Z(n_2626));
	notech_ao4 i_146933461(.A(n_1986), .B(n_17372), .C(n_1985), .D(n_17380),
		 .Z(n_2628));
	notech_ao4 i_147633454(.A(n_59838), .B(n_17423), .C(n_59825), .D(n_17487
		), .Z(n_2630));
	notech_and4 i_147933451(.A(n_2626), .B(n_2628), .C(n_2630), .D(n_1881), 
		.Z(n_2631));
	notech_ao4 i_147033460(.A(n_59786), .B(n_17388), .C(n_59773), .D(n_17404
		), .Z(n_2632));
	notech_ao4 i_147133459(.A(n_59812), .B(n_17412), .C(n_59799), .D(n_17396
		), .Z(n_2633));
	notech_and3 i_147733453(.A(n_2633), .B(n_2632), .C(n_1894), .Z(n_2635)
		);
	notech_ao4 i_147433456(.A(n_59890), .B(n_17439), .C(n_59877), .D(n_17503
		), .Z(n_2636));
	notech_ao4 i_147533455(.A(n_59916), .B(n_17471), .C(n_59903), .D(n_17455
		), .Z(n_2637));
	notech_ao4 i_149833432(.A(n_59975), .B(n_17357), .C(n_59956), .D(n_17365
		), .Z(n_2640));
	notech_ao4 i_150033430(.A(n_59864), .B(n_17373), .C(n_59851), .D(n_17381
		), .Z(n_2642));
	notech_ao4 i_150733423(.A(n_59838), .B(n_17425), .C(n_59825), .D(n_17489
		), .Z(n_2644));
	notech_and4 i_151033420(.A(n_2640), .B(n_2642), .C(n_2644), .D(n_1897), 
		.Z(n_2645));
	notech_ao4 i_150133429(.A(n_59786), .B(n_17389), .C(n_59773), .D(n_17405
		), .Z(n_2646));
	notech_ao4 i_150233428(.A(n_59812), .B(n_17413), .C(n_59799), .D(n_17397
		), .Z(n_2647));
	notech_and3 i_150833422(.A(n_2647), .B(n_2646), .C(n_1910), .Z(n_2649)
		);
	notech_ao4 i_150533425(.A(n_59890), .B(n_17441), .C(n_59877), .D(n_17505
		), .Z(n_2650));
	notech_ao4 i_150633424(.A(n_59916), .B(n_17473), .C(n_59903), .D(n_17457
		), .Z(n_2651));
	notech_ao4 i_152933401(.A(n_59975), .B(n_17358), .C(n_59956), .D(n_17366
		), .Z(n_2654));
	notech_ao4 i_153133399(.A(n_59864), .B(n_17374), .C(n_59851), .D(n_17382
		), .Z(n_2656));
	notech_ao4 i_153833392(.A(n_59838), .B(n_17427), .C(n_59825), .D(n_17491
		), .Z(n_2658));
	notech_and4 i_154133389(.A(n_2654), .B(n_2656), .C(n_2658), .D(n_1913), 
		.Z(n_2659));
	notech_ao4 i_153233398(.A(n_59786), .B(n_17390), .C(n_59773), .D(n_17406
		), .Z(n_2660));
	notech_ao4 i_153333397(.A(n_59812), .B(n_17414), .C(n_59799), .D(n_17398
		), .Z(n_2661));
	notech_and3 i_153933391(.A(n_2661), .B(n_2660), .C(n_1926), .Z(n_2663)
		);
	notech_ao4 i_153633394(.A(n_59890), .B(n_17443), .C(n_59877), .D(n_17507
		), .Z(n_2664));
	notech_ao4 i_153733393(.A(n_59916), .B(n_17475), .C(n_59903), .D(n_17459
		), .Z(n_2665));
	notech_ao4 i_156033370(.A(n_59975), .B(n_17359), .C(n_59957), .D(n_17367
		), .Z(n_2668));
	notech_ao4 i_156233368(.A(n_59864), .B(n_17375), .C(n_59851), .D(n_17383
		), .Z(n_2670));
	notech_ao4 i_156933361(.A(n_59838), .B(n_17429), .C(n_59825), .D(n_17493
		), .Z(n_2672));
	notech_and4 i_157233358(.A(n_2668), .B(n_2670), .C(n_2672), .D(n_1929), 
		.Z(n_2673));
	notech_ao4 i_156333367(.A(n_59786), .B(n_17391), .C(n_59773), .D(n_17407
		), .Z(n_2674));
	notech_ao4 i_156433366(.A(n_59812), .B(n_17415), .C(n_59799), .D(n_17399
		), .Z(n_2675));
	notech_and3 i_157033360(.A(n_2675), .B(n_2674), .C(n_1942), .Z(n_2677)
		);
	notech_ao4 i_156733363(.A(n_59890), .B(n_17445), .C(n_59877), .D(n_17509
		), .Z(n_2678));
	notech_ao4 i_156833362(.A(n_59916), .B(n_17477), .C(n_59903), .D(n_17461
		), .Z(n_2679));
	notech_ao4 i_159133339(.A(n_59976), .B(n_17360), .C(n_59957), .D(n_17368
		), .Z(n_2682));
	notech_ao4 i_159333337(.A(n_59864), .B(n_17376), .C(n_59851), .D(n_17384
		), .Z(n_2684));
	notech_ao4 i_160033330(.A(n_59838), .B(n_17431), .C(n_59825), .D(n_17495
		), .Z(n_2686));
	notech_and4 i_160333327(.A(n_2682), .B(n_2684), .C(n_2686), .D(n_1945), 
		.Z(n_2687));
	notech_ao4 i_159433336(.A(n_59786), .B(n_17392), .C(n_59773), .D(n_17408
		), .Z(n_2688));
	notech_ao4 i_159533335(.A(n_59812), .B(n_17416), .C(n_59799), .D(n_17400
		), .Z(n_2689));
	notech_and3 i_160133329(.A(n_2689), .B(n_2688), .C(n_1958), .Z(n_2691)
		);
	notech_ao4 i_159833332(.A(n_59890), .B(n_17447), .C(n_59877), .D(n_17511
		), .Z(n_2692));
	notech_ao4 i_159933331(.A(n_59916), .B(n_17479), .C(n_59903), .D(n_17463
		), .Z(n_2693));
	notech_ao4 i_162233308(.A(n_59976), .B(n_17372), .C(n_59957), .D(n_17380
		), .Z(n_2696));
	notech_ao4 i_162433306(.A(n_59864), .B(n_17388), .C(n_59851), .D(n_17396
		), .Z(n_2698));
	notech_ao4 i_163133299(.A(n_59838), .B(n_17455), .C(n_59825), .D(n_17519
		), .Z(n_2700));
	notech_and4 i_163433296(.A(n_2696), .B(n_2698), .C(n_2700), .D(n_1961), 
		.Z(n_2701));
	notech_ao4 i_162533305(.A(n_59786), .B(n_17404), .C(n_59773), .D(n_17423
		), .Z(n_2702));
	notech_ao4 i_162633304(.A(n_59812), .B(n_17439), .C(n_59799), .D(n_17412
		), .Z(n_2703));
	notech_and3 i_163233298(.A(n_2703), .B(n_2702), .C(n_1974), .Z(n_2705)
		);
	notech_ao4 i_162933301(.A(n_59890), .B(n_17471), .C(n_59877), .D(n_17535
		), .Z(n_2706));
	notech_ao4 i_163033300(.A(n_59916), .B(n_17503), .C(n_59903), .D(n_17487
		), .Z(n_2707));
	notech_ao4 i_216032776(.A(n_61359), .B(n_17760), .C(n_61153), .D(n_17475
		), .Z(n_2710));
	notech_ao4 i_219232744(.A(n_61359), .B(n_17752), .C(n_61153), .D(n_17459
		), .Z(n_2711));
	notech_ao4 i_222432712(.A(n_61359), .B(n_17744), .C(n_61153), .D(n_17443
		), .Z(n_2712));
	notech_ao4 i_225632680(.A(n_61359), .B(n_17736), .C(n_61153), .D(n_17427
		), .Z(n_2713));
	notech_nand3 i_68(.A(n_59664), .B(n_59937), .C(queue[14]), .Z(n_2714));
	notech_or2 i_69(.A(n_59957), .B(n_17329), .Z(n_2729));
	notech_nand3 i_1524981(.A(n_3104), .B(n_3097), .C(n_2714), .Z(squeue[14]
		));
	notech_nand3 i_161(.A(n_59664), .B(n_59937), .C(queue[54]), .Z(n_2730)
		);
	notech_or2 i_162(.A(n_59956), .B(n_17369), .Z(n_2745));
	notech_nand3 i_5525021(.A(n_3118), .B(n_3111), .C(n_2730), .Z(squeue[54]
		));
	notech_nand3 i_347(.A(n_59664), .B(n_59937), .C(queue[60]), .Z(n_2746)
		);
	notech_or2 i_348(.A(n_59956), .B(n_17375), .Z(n_2761));
	notech_nand3 i_6125027(.A(n_3132), .B(n_3125), .C(n_2746), .Z(squeue[60]
		));
	notech_nand3 i_409(.A(n_59664), .B(n_59937), .C(queue[62]), .Z(n_2762)
		);
	notech_or2 i_410(.A(n_59956), .B(n_17377), .Z(n_2777));
	notech_nand3 i_6325029(.A(n_3146), .B(n_3139), .C(n_2762), .Z(squeue[62]
		));
	notech_nand3 i_471(.A(n_59664), .B(n_59937), .C(queue[64]), .Z(n_2778)
		);
	notech_or2 i_472(.A(n_59956), .B(n_17379), .Z(n_2793));
	notech_nand3 i_6525031(.A(n_3160), .B(n_3153), .C(n_2778), .Z(squeue[64]
		));
	notech_nand3 i_564(.A(n_59664), .B(n_59937), .C(queue[68]), .Z(n_2794)
		);
	notech_or2 i_565(.A(n_59952), .B(n_17383), .Z(n_2809));
	notech_nand3 i_6925035(.A(n_3174), .B(n_3167), .C(n_2794), .Z(squeue[68]
		));
	notech_nand3 i_626(.A(n_59664), .B(n_59937), .C(queue[70]), .Z(n_2810)
		);
	notech_or2 i_627(.A(n_59952), .B(n_17385), .Z(n_2825));
	notech_nand3 i_7125037(.A(n_3188), .B(n_3181), .C(n_2810), .Z(squeue[70]
		));
	notech_nand3 i_781(.A(n_59664), .B(n_59937), .C(queue[75]), .Z(n_2826)
		);
	notech_or2 i_782(.A(n_59952), .B(n_17390), .Z(n_2841));
	notech_nand3 i_7625042(.A(n_3202), .B(n_3195), .C(n_2826), .Z(squeue[75]
		));
	notech_nand3 i_812(.A(n_59664), .B(n_59937), .C(queue[76]), .Z(n_2842)
		);
	notech_or2 i_813(.A(n_59952), .B(n_17391), .Z(n_2857));
	notech_nand3 i_7725043(.A(n_3216), .B(n_3209), .C(n_2842), .Z(squeue[76]
		));
	notech_nand3 i_874(.A(n_59664), .B(n_59937), .C(queue[78]), .Z(n_2858)
		);
	notech_or2 i_875(.A(n_59952), .B(n_17393), .Z(n_2873));
	notech_nand3 i_7925045(.A(n_3230), .B(n_3223), .C(n_2858), .Z(squeue[78]
		));
	notech_nand3 i_1060(.A(n_59664), .B(n_59938), .C(queue[84]), .Z(n_2874)
		);
	notech_or2 i_1061(.A(n_59952), .B(n_17399), .Z(n_2889));
	notech_nand3 i_8525051(.A(n_3244), .B(n_3237), .C(n_2874), .Z(squeue[84]
		));
	notech_nand3 i_1122(.A(n_59664), .B(n_59938), .C(queue[86]), .Z(n_2890)
		);
	notech_or2 i_1123(.A(n_59952), .B(n_17401), .Z(n_2905));
	notech_nand3 i_8725053(.A(n_3258), .B(n_3251), .C(n_2890), .Z(squeue[86]
		));
	notech_nand3 i_1308(.A(n_59664), .B(n_59937), .C(queue[92]), .Z(n_2906)
		);
	notech_or2 i_1309(.A(n_59952), .B(n_17407), .Z(n_2921));
	notech_nand3 i_9325059(.A(n_3272), .B(n_3265), .C(n_2906), .Z(squeue[92]
		));
	notech_nand3 i_1370(.A(n_59664), .B(n_59937), .C(queue[94]), .Z(n_2922)
		);
	notech_or2 i_1371(.A(n_59956), .B(n_17409), .Z(n_2937));
	notech_nand3 i_9525061(.A(n_3286), .B(n_3279), .C(n_2922), .Z(squeue[94]
		));
	notech_nand3 i_1556(.A(n_59664), .B(n_59937), .C(queue[100]), .Z(n_2938)
		);
	notech_or2 i_1557(.A(n_59956), .B(n_17415), .Z(n_2956));
	notech_nand3 i_10125067(.A(n_3300), .B(n_3293), .C(n_2938), .Z(squeue[
		100]));
	notech_nand3 i_1618(.A(n_59664), .B(n_59937), .C(queue[102]), .Z(n_2957)
		);
	notech_or2 i_1619(.A(n_59956), .B(n_17417), .Z(n_2972));
	notech_nand3 i_10325069(.A(n_3314), .B(n_3307), .C(n_2957), .Z(squeue[
		102]));
	notech_nand3 i_1804(.A(n_59662), .B(n_59937), .C(queue[108]), .Z(n_2973)
		);
	notech_or2 i_1805(.A(n_59956), .B(n_17429), .Z(n_2988));
	notech_nand3 i_10925075(.A(n_3328), .B(n_3321), .C(n_2973), .Z(squeue[
		108]));
	notech_nand3 i_1866(.A(n_59662), .B(n_59933), .C(queue[110]), .Z(n_2989)
		);
	notech_or2 i_1867(.A(n_59952), .B(n_17433), .Z(n_3004));
	notech_nand3 i_11125077(.A(n_3342), .B(n_3335), .C(n_2989), .Z(squeue[
		110]));
	notech_nand3 i_2052(.A(n_59662), .B(n_59933), .C(queue[116]), .Z(n_3005)
		);
	notech_or2 i_2053(.A(n_59952), .B(n_17445), .Z(n_3020));
	notech_nand3 i_11725083(.A(n_3356), .B(n_3349), .C(n_3005), .Z(squeue[
		116]));
	notech_nand3 i_2114(.A(n_59662), .B(n_59933), .C(queue[118]), .Z(n_3021)
		);
	notech_or2 i_2115(.A(n_59956), .B(n_17449), .Z(n_3036));
	notech_nand3 i_11925085(.A(n_3370), .B(n_3363), .C(n_3021), .Z(squeue[
		118]));
	notech_nand3 i_2300(.A(n_59662), .B(n_59933), .C(queue[124]), .Z(n_3037)
		);
	notech_or2 i_2301(.A(n_59956), .B(n_17461), .Z(n_3052));
	notech_nand3 i_12525091(.A(n_3384), .B(n_3377), .C(n_3037), .Z(squeue[
		124]));
	notech_nand3 i_2362(.A(n_59662), .B(n_59933), .C(queue[126]), .Z(n_3053)
		);
	notech_or2 i_2363(.A(n_59959), .B(n_17465), .Z(n_3068));
	notech_nand3 i_12725093(.A(n_3398), .B(n_3391), .C(n_3053), .Z(squeue[
		126]));
	notech_and2 i_1(.A(addrshft[1]), .B(n_17679), .Z(n_3069));
	notech_nor2 i_60(.A(addrshft[5]), .B(addrshft[4]), .Z(n_3070));
	notech_and3 i_6(.A(addrshft[0]), .B(n_3070), .C(addrshft[3]), .Z(n_3072)
		);
	notech_nao3 i_1331200(.A(addrshft[1]), .B(n_3072), .C(addrshft[2]), .Z(n_1321
		));
	notech_ao3 i_9(.A(addrshft[3]), .B(n_3070), .C(addrshft[0]), .Z(n_3074)
		);
	notech_nao3 i_1331195(.A(addrshft[1]), .B(n_3074), .C(addrshft[2]), .Z(n_1318
		));
	notech_and2 i_5(.A(addrshft[1]), .B(addrshft[2]), .Z(n_3076));
	notech_nand3 i_1331220(.A(addrshft[1]), .B(addrshft[2]), .C(n_3072), .Z(n_1315
		));
	notech_nand3 i_1331215(.A(addrshft[1]), .B(addrshft[2]), .C(n_3074), .Z(n_1314
		));
	notech_and2 i_7(.A(addrshft[2]), .B(n_17678), .Z(n_3078));
	notech_nao3 i_1331210(.A(addrshft[2]), .B(n_3072), .C(addrshft[1]), .Z(n_1311
		));
	notech_nao3 i_1331205(.A(addrshft[2]), .B(n_3074), .C(addrshft[1]), .Z(n_1310
		));
	notech_and4 i_18(.A(n_59731), .B(n_59715), .C(n_59699), .D(n_59683), .Z(n_3080
		));
	notech_and3 i_5303(.A(n_59763), .B(n_59747), .C(n_3080), .Z(n_3081));
	notech_ao3 i_2(.A(addrshft[0]), .B(n_3070), .C(addrshft[3]), .Z(n_3082)
		);
	notech_nand3 i_1331180(.A(n_3082), .B(addrshft[1]), .C(addrshft[2]), .Z(n_1305
		));
	notech_nand3 i_1331170(.A(n_60101), .B(addrshft[2]), .C(n_17678), .Z(n_1304
		));
	notech_or4 i_10(.A(addrshft[5]), .B(addrshft[4]), .C(addrshft[0]), .D(addrshft
		[3]), .Z(n_3084));
	notech_nao3 i_1331175(.A(addrshft[1]), .B(addrshft[2]), .C(n_3084), .Z(n_1301
		));
	notech_nao3 i_1331165(.A(addrshft[2]), .B(n_17678), .C(n_3084), .Z(n_1300
		));
	notech_and2 i_8(.A(n_17678), .B(n_17679), .Z(n_3086));
	notech_nand2 i_1331190(.A(n_3086), .B(n_3072), .Z(n_1297));
	notech_nand2 i_1331185(.A(n_61409), .B(n_3074), .Z(n_1296));
	notech_and4 i_14(.A(n_60059), .B(n_60043), .C(n_60027), .D(n_60011), .Z(n_3088
		));
	notech_nand3 i_3(.A(n_3082), .B(addrshft[1]), .C(n_17679), .Z(n_1292));
	notech_nao3 i_1331155(.A(addrshft[1]), .B(n_17679), .C(n_3084), .Z(n_1291
		));
	notech_nand3 i_1331150(.A(n_3082), .B(n_17678), .C(n_17679), .Z(n_1290)
		);
	notech_and3 i_5322(.A(n_59994), .B(n_59976), .C(n_59959), .Z(n_3091));
	notech_ao4 i_70(.A(n_60027), .B(n_17337), .C(n_60011), .D(n_17353), .Z(n_3092
		));
	notech_ao4 i_71(.A(n_59976), .B(n_17321), .C(n_59683), .D(n_17433), .Z(n_3094
		));
	notech_ao4 i_72(.A(n_59715), .B(n_17409), .C(n_59699), .D(n_17417), .Z(n_3095
		));
	notech_and4 i_81(.A(n_3095), .B(n_3094), .C(n_3092), .D(n_2729), .Z(n_3097
		));
	notech_ao4 i_73(.A(n_59747), .B(n_17393), .C(n_59731), .D(n_17401), .Z(n_3098
		));
	notech_ao4 i_74(.A(n_60043), .B(n_17377), .C(n_59763), .D(n_17385), .Z(n_3099
		));
	notech_ao4 i_75(.A(n_60075), .B(n_17361), .C(n_60059), .D(n_17369), .Z(n_3101
		));
	notech_ao4 i_76(.A(n_59994), .B(n_17313), .C(n_60091), .D(n_17345), .Z(n_3102
		));
	notech_and4 i_82(.A(n_3102), .B(n_3101), .C(n_3099), .D(n_3098), .Z(n_3104
		));
	notech_ao4 i_163(.A(n_60023), .B(n_17377), .C(n_60007), .D(n_17393), .Z(n_3106
		));
	notech_ao4 i_164(.A(n_59975), .B(n_17361), .C(n_59679), .D(n_17513), .Z(n_3108
		));
	notech_ao4 i_165(.A(n_59711), .B(n_17481), .C(n_59695), .D(n_17497), .Z(n_3109
		));
	notech_and4 i_174(.A(n_3109), .B(n_3108), .C(n_3106), .D(n_2745), .Z(n_3111
		));
	notech_ao4 i_166(.A(n_59743), .B(n_17449), .C(n_59727), .D(n_17465), .Z(n_3112
		));
	notech_ao4 i_167(.A(n_60039), .B(n_17417), .C(n_59759), .D(n_17433), .Z(n_3113
		));
	notech_ao4 i_168(.A(n_60075), .B(n_17401), .C(n_60055), .D(n_17409), .Z(n_3115
		));
	notech_ao4 i_169(.A(n_59994), .B(n_17353), .C(n_60091), .D(n_17385), .Z(n_3116
		));
	notech_and4 i_175(.A(n_3116), .B(n_3115), .C(n_3113), .D(n_3112), .Z(n_3118
		));
	notech_ao4 i_349(.A(n_60027), .B(n_17383), .C(n_60011), .D(n_17399), .Z(n_3120
		));
	notech_ao4 i_350(.A(n_59975), .B(n_17367), .C(n_59683), .D(n_17525), .Z(n_3122
		));
	notech_ao4 i_351(.A(n_59715), .B(n_17493), .C(n_59699), .D(n_17509), .Z(n_3123
		));
	notech_and4 i_360(.A(n_3123), .B(n_3122), .C(n_3120), .D(n_2761), .Z(n_3125
		));
	notech_ao4 i_352(.A(n_59747), .B(n_17461), .C(n_59731), .D(n_17477), .Z(n_3126
		));
	notech_ao4 i_353(.A(n_60043), .B(n_17429), .C(n_59763), .D(n_17445), .Z(n_3127
		));
	notech_ao4 i_354(.A(n_60071), .B(n_17407), .C(n_60059), .D(n_17415), .Z(n_3129
		));
	notech_ao4 i_355(.A(n_59994), .B(n_17359), .C(n_60087), .D(n_17391), .Z(n_3130
		));
	notech_and4 i_361(.A(n_3130), .B(n_3129), .C(n_3127), .D(n_3126), .Z(n_3132
		));
	notech_ao4 i_411(.A(n_60027), .B(n_17385), .C(n_60011), .D(n_17401), .Z(n_3134
		));
	notech_ao4 i_412(.A(n_59975), .B(n_17369), .C(n_59683), .D(n_17529), .Z(n_3136
		));
	notech_ao4 i_413(.A(n_59715), .B(n_17497), .C(n_59699), .D(n_17513), .Z(n_3137
		));
	notech_and4 i_422(.A(n_3137), .B(n_3136), .C(n_3134), .D(n_2777), .Z(n_3139
		));
	notech_ao4 i_414(.A(n_59747), .B(n_17465), .C(n_59731), .D(n_17481), .Z(n_3140
		));
	notech_ao4 i_415(.A(n_60043), .B(n_17433), .C(n_59763), .D(n_17449), .Z(n_3141
		));
	notech_ao4 i_416(.A(n_60075), .B(n_17409), .C(n_60059), .D(n_17417), .Z(n_3143
		));
	notech_ao4 i_417(.A(n_59994), .B(n_17361), .C(n_60091), .D(n_17393), .Z(n_3144
		));
	notech_and4 i_423(.A(n_3144), .B(n_3143), .C(n_3141), .D(n_3140), .Z(n_3146
		));
	notech_ao4 i_473(.A(n_60027), .B(n_17387), .C(n_60011), .D(n_17403), .Z(n_3148
		));
	notech_ao4 i_474(.A(n_59975), .B(n_17371), .C(n_59683), .D(n_17533), .Z(n_3150
		));
	notech_ao4 i_475(.A(n_59715), .B(n_17501), .C(n_59699), .D(n_17517), .Z(n_3151
		));
	notech_and4 i_484(.A(n_3151), .B(n_3150), .C(n_3148), .D(n_2793), .Z(n_3153
		));
	notech_ao4 i_476(.A(n_59747), .B(n_17469), .C(n_59731), .D(n_17485), .Z(n_3154
		));
	notech_ao4 i_477(.A(n_60043), .B(n_17437), .C(n_59763), .D(n_17453), .Z(n_3155
		));
	notech_ao4 i_478(.A(n_60075), .B(n_17411), .C(n_60059), .D(n_17421), .Z(n_3157
		));
	notech_ao4 i_479(.A(n_59994), .B(n_17363), .C(n_60091), .D(n_17395), .Z(n_3158
		));
	notech_and4 i_485(.A(n_3158), .B(n_3157), .C(n_3155), .D(n_3154), .Z(n_3160
		));
	notech_ao4 i_566(.A(n_60027), .B(n_17391), .C(n_60011), .D(n_17407), .Z(n_3162
		));
	notech_ao4 i_567(.A(n_59971), .B(n_17375), .C(n_59683), .D(n_17541), .Z(n_3164
		));
	notech_ao4 i_568(.A(n_59715), .B(n_17509), .C(n_59699), .D(n_17525), .Z(n_3165
		));
	notech_and4 i_577(.A(n_3165), .B(n_3164), .C(n_3162), .D(n_2809), .Z(n_3167
		));
	notech_ao4 i_569(.A(n_59747), .B(n_17477), .C(n_59731), .D(n_17493), .Z(n_3168
		));
	notech_ao4 i_570(.A(n_60043), .B(n_17445), .C(n_59763), .D(n_17461), .Z(n_3169
		));
	notech_ao4 i_571(.A(n_60075), .B(n_17415), .C(n_60059), .D(n_17429), .Z(n_3171
		));
	notech_ao4 i_572(.A(n_59994), .B(n_17367), .C(n_60091), .D(n_17399), .Z(n_3172
		));
	notech_and4 i_578(.A(n_3172), .B(n_3171), .C(n_3169), .D(n_3168), .Z(n_3174
		));
	notech_ao4 i_628(.A(n_60027), .B(n_17393), .C(n_60011), .D(n_17409), .Z(n_3176
		));
	notech_ao4 i_629(.A(n_59971), .B(n_17377), .C(n_59683), .D(n_17545), .Z(n_3178
		));
	notech_ao4 i_630(.A(n_59715), .B(n_17513), .C(n_59699), .D(n_17529), .Z(n_3179
		));
	notech_and4 i_639(.A(n_3179), .B(n_3178), .C(n_3176), .D(n_2825), .Z(n_3181
		));
	notech_ao4 i_631(.A(n_59747), .B(n_17481), .C(n_59731), .D(n_17497), .Z(n_3182
		));
	notech_ao4 i_632(.A(n_60043), .B(n_17449), .C(n_59763), .D(n_17465), .Z(n_3183
		));
	notech_ao4 i_633(.A(n_60075), .B(n_17417), .C(n_60059), .D(n_17433), .Z(n_3185
		));
	notech_ao4 i_634(.A(n_59994), .B(n_17369), .C(n_60091), .D(n_17401), .Z(n_3186
		));
	notech_and4 i_640(.A(n_3186), .B(n_3185), .C(n_3183), .D(n_3182), .Z(n_3188
		));
	notech_ao4 i_783(.A(n_60027), .B(n_17398), .C(n_60011), .D(n_17414), .Z(n_3190
		));
	notech_ao4 i_784(.A(n_59971), .B(n_17382), .C(n_59683), .D(n_17555), .Z(n_3192
		));
	notech_ao4 i_785(.A(n_59715), .B(n_17523), .C(n_59699), .D(n_17539), .Z(n_3193
		));
	notech_and4 i_794(.A(n_3193), .B(n_3192), .C(n_3190), .D(n_2841), .Z(n_3195
		));
	notech_ao4 i_786(.A(n_59747), .B(n_17491), .C(n_59731), .D(n_17507), .Z(n_3196
		));
	notech_ao4 i_787(.A(n_60043), .B(n_17459), .C(n_59763), .D(n_17475), .Z(n_3197
		));
	notech_ao4 i_788(.A(n_60075), .B(n_17427), .C(n_60059), .D(n_17443), .Z(n_3199
		));
	notech_ao4 i_789(.A(n_59994), .B(n_17374), .C(n_60091), .D(n_17406), .Z(n_3200
		));
	notech_and4 i_795(.A(n_3200), .B(n_3199), .C(n_3197), .D(n_3196), .Z(n_3202
		));
	notech_ao4 i_814(.A(n_60023), .B(n_17399), .C(n_60007), .D(n_17415), .Z(n_3204
		));
	notech_ao4 i_815(.A(n_59971), .B(n_17383), .C(n_59679), .D(n_17557), .Z(n_3206
		));
	notech_ao4 i_816(.A(n_59711), .B(n_17525), .C(n_59695), .D(n_17541), .Z(n_3207
		));
	notech_and4 i_825(.A(n_3207), .B(n_3206), .C(n_3204), .D(n_2857), .Z(n_3209
		));
	notech_ao4 i_817(.A(n_59743), .B(n_17493), .C(n_59727), .D(n_17509), .Z(n_3210
		));
	notech_ao4 i_818(.A(n_60039), .B(n_17461), .C(n_59759), .D(n_17477), .Z(n_3211
		));
	notech_ao4 i_819(.A(n_60075), .B(n_17429), .C(n_60055), .D(n_17445), .Z(n_3213
		));
	notech_ao4 i_820(.A(n_59994), .B(n_17375), .C(n_60091), .D(n_17407), .Z(n_3214
		));
	notech_and4 i_826(.A(n_3214), .B(n_3213), .C(n_3211), .D(n_3210), .Z(n_3216
		));
	notech_ao4 i_876(.A(n_60023), .B(n_17401), .C(n_60007), .D(n_17417), .Z(n_3218
		));
	notech_ao4 i_877(.A(n_59971), .B(n_17385), .C(n_59679), .D(n_17561), .Z(n_3220
		));
	notech_ao4 i_878(.A(n_59711), .B(n_17529), .C(n_59695), .D(n_17545), .Z(n_3221
		));
	notech_and4 i_887(.A(n_3221), .B(n_3220), .C(n_3218), .D(n_2873), .Z(n_3223
		));
	notech_ao4 i_879(.A(n_59743), .B(n_17497), .C(n_59727), .D(n_17513), .Z(n_3224
		));
	notech_ao4 i_880(.A(n_60039), .B(n_17465), .C(n_59759), .D(n_17481), .Z(n_3225
		));
	notech_ao4 i_881(.A(n_60071), .B(n_17433), .C(n_60055), .D(n_17449), .Z(n_3227
		));
	notech_ao4 i_882(.A(n_59989), .B(n_17377), .C(n_60087), .D(n_17409), .Z(n_3228
		));
	notech_and4 i_888(.A(n_3228), .B(n_3227), .C(n_3225), .D(n_3224), .Z(n_3230
		));
	notech_ao4 i_1062(.A(n_60023), .B(n_17407), .C(n_60007), .D(n_17429), .Z
		(n_3232));
	notech_ao4 i_1063(.A(n_59971), .B(n_17391), .C(n_59679), .D(n_17573), .Z
		(n_3234));
	notech_ao4 i_1064(.A(n_59711), .B(n_17541), .C(n_59695), .D(n_17557), .Z
		(n_3235));
	notech_and4 i_1073(.A(n_3235), .B(n_3234), .C(n_3232), .D(n_2889), .Z(n_3237
		));
	notech_ao4 i_1065(.A(n_59743), .B(n_17509), .C(n_59727), .D(n_17525), .Z
		(n_3238));
	notech_ao4 i_1066(.A(n_60039), .B(n_17477), .C(n_59759), .D(n_17493), .Z
		(n_3239));
	notech_ao4 i_1067(.A(n_60071), .B(n_17445), .C(n_60055), .D(n_17461), .Z
		(n_3241));
	notech_ao4 i_1068(.A(n_59989), .B(n_17383), .C(n_60087), .D(n_17415), .Z
		(n_3242));
	notech_and4 i_1074(.A(n_3242), .B(n_3241), .C(n_3239), .D(n_3238), .Z(n_3244
		));
	notech_ao4 i_1124(.A(n_60023), .B(n_17409), .C(n_60007), .D(n_17433), .Z
		(n_3246));
	notech_ao4 i_1125(.A(n_59971), .B(n_17393), .C(n_59679), .D(n_17577), .Z
		(n_3248));
	notech_ao4 i_1126(.A(n_59711), .B(n_17545), .C(n_59695), .D(n_17561), .Z
		(n_3249));
	notech_and4 i_1135(.A(n_3249), .B(n_3248), .C(n_3246), .D(n_2905), .Z(n_3251
		));
	notech_ao4 i_1127(.A(n_59743), .B(n_17513), .C(n_59727), .D(n_17529), .Z
		(n_3252));
	notech_ao4 i_1128(.A(n_60039), .B(n_17481), .C(n_59759), .D(n_17497), .Z
		(n_3253));
	notech_ao4 i_1129(.A(n_60071), .B(n_17449), .C(n_60055), .D(n_17465), .Z
		(n_3255));
	notech_ao4 i_1130(.A(n_59989), .B(n_17385), .C(n_60087), .D(n_17417), .Z
		(n_3256));
	notech_and4 i_1136(.A(n_3256), .B(n_3255), .C(n_3253), .D(n_3252), .Z(n_3258
		));
	notech_ao4 i_1310(.A(n_60023), .B(n_17415), .C(n_60007), .D(n_17445), .Z
		(n_3260));
	notech_ao4 i_1311(.A(n_59971), .B(n_17399), .C(n_59679), .D(n_17589), .Z
		(n_3262));
	notech_ao4 i_1312(.A(n_59711), .B(n_17557), .C(n_59695), .D(n_17573), .Z
		(n_3263));
	notech_and4 i_1321(.A(n_3263), .B(n_3262), .C(n_3260), .D(n_2921), .Z(n_3265
		));
	notech_ao4 i_1313(.A(n_59743), .B(n_17525), .C(n_59727), .D(n_17541), .Z
		(n_3266));
	notech_ao4 i_1314(.A(n_60039), .B(n_17493), .C(n_59759), .D(n_17509), .Z
		(n_3267));
	notech_ao4 i_1315(.A(n_60071), .B(n_17461), .C(n_60055), .D(n_17477), .Z
		(n_3269));
	notech_ao4 i_1316(.A(n_59989), .B(n_17391), .C(n_60087), .D(n_17429), .Z
		(n_3270));
	notech_and4 i_1322(.A(n_3270), .B(n_3269), .C(n_3267), .D(n_3266), .Z(n_3272
		));
	notech_ao4 i_1372(.A(n_60023), .B(n_17417), .C(n_60007), .D(n_17449), .Z
		(n_3274));
	notech_ao4 i_1373(.A(n_59975), .B(n_17401), .C(n_59679), .D(n_17593), .Z
		(n_3276));
	notech_ao4 i_1374(.A(n_59711), .B(n_17561), .C(n_59695), .D(n_17577), .Z
		(n_3277));
	notech_and4 i_1383(.A(n_3277), .B(n_3276), .C(n_3274), .D(n_2937), .Z(n_3279
		));
	notech_ao4 i_1375(.A(n_59743), .B(n_17529), .C(n_59727), .D(n_17545), .Z
		(n_3280));
	notech_ao4 i_1376(.A(n_60039), .B(n_17497), .C(n_59759), .D(n_17513), .Z
		(n_3281));
	notech_ao4 i_1377(.A(n_60071), .B(n_17465), .C(n_60055), .D(n_17481), .Z
		(n_3283));
	notech_ao4 i_1378(.A(n_59989), .B(n_17393), .C(n_60087), .D(n_17433), .Z
		(n_3284));
	notech_and4 i_1384(.A(n_3284), .B(n_3283), .C(n_3281), .D(n_3280), .Z(n_3286
		));
	notech_ao4 i_1558(.A(n_60023), .B(n_17429), .C(n_60007), .D(n_17461), .Z
		(n_3288));
	notech_ao4 i_1559(.A(n_59975), .B(n_17407), .C(n_59679), .D(n_17605), .Z
		(n_3290));
	notech_ao4 i_1560(.A(n_59711), .B(n_17573), .C(n_59695), .D(n_17589), .Z
		(n_3291));
	notech_and4 i_1569(.A(n_3291), .B(n_3290), .C(n_3288), .D(n_2956), .Z(n_3293
		));
	notech_ao4 i_1561(.A(n_59743), .B(n_17541), .C(n_59727), .D(n_17557), .Z
		(n_3294));
	notech_ao4 i_1562(.A(n_60039), .B(n_17509), .C(n_59759), .D(n_17525), .Z
		(n_3295));
	notech_ao4 i_1563(.A(n_60071), .B(n_17477), .C(n_60055), .D(n_17493), .Z
		(n_3297));
	notech_ao4 i_1564(.A(n_59989), .B(n_17399), .C(n_60087), .D(n_17445), .Z
		(n_3298));
	notech_and4 i_1570(.A(n_3298), .B(n_3297), .C(n_3295), .D(n_3294), .Z(n_3300
		));
	notech_ao4 i_1620(.A(n_60023), .B(n_17433), .C(n_60007), .D(n_17465), .Z
		(n_3302));
	notech_ao4 i_1621(.A(n_59975), .B(n_17409), .C(n_59679), .D(n_17609), .Z
		(n_3304));
	notech_ao4 i_1622(.A(n_59711), .B(n_17577), .C(n_59695), .D(n_17593), .Z
		(n_3305));
	notech_and4 i_1631(.A(n_3305), .B(n_3304), .C(n_3302), .D(n_2972), .Z(n_3307
		));
	notech_ao4 i_1623(.A(n_59743), .B(n_17545), .C(n_59727), .D(n_17561), .Z
		(n_3308));
	notech_ao4 i_1624(.A(n_60039), .B(n_17513), .C(n_59759), .D(n_17529), .Z
		(n_3309));
	notech_ao4 i_1625(.A(n_60071), .B(n_17481), .C(n_60055), .D(n_17497), .Z
		(n_3311));
	notech_ao4 i_1626(.A(n_59994), .B(n_17401), .C(n_60087), .D(n_17449), .Z
		(n_3312));
	notech_and4 i_1632(.A(n_3312), .B(n_3311), .C(n_3309), .D(n_3308), .Z(n_3314
		));
	notech_ao4 i_1806(.A(n_60023), .B(n_17445), .C(n_60007), .D(n_17477), .Z
		(n_3316));
	notech_ao4 i_1807(.A(n_59975), .B(n_17415), .C(n_59679), .D(n_17621), .Z
		(n_3318));
	notech_ao4 i_1808(.A(n_59711), .B(n_17589), .C(n_59695), .D(n_17605), .Z
		(n_3319));
	notech_and4 i_1817(.A(n_3319), .B(n_3318), .C(n_3316), .D(n_2988), .Z(n_3321
		));
	notech_ao4 i_1809(.A(n_59743), .B(n_17557), .C(n_59727), .D(n_17573), .Z
		(n_3322));
	notech_ao4 i_1810(.A(n_60039), .B(n_17525), .C(n_59759), .D(n_17541), .Z
		(n_3323));
	notech_ao4 i_1811(.A(n_60071), .B(n_17493), .C(n_60055), .D(n_17509), .Z
		(n_3325));
	notech_ao4 i_1812(.A(n_59994), .B(n_17407), .C(n_60087), .D(n_17461), .Z
		(n_3326));
	notech_and4 i_1818(.A(n_3326), .B(n_3325), .C(n_3323), .D(n_3322), .Z(n_3328
		));
	notech_ao4 i_1868(.A(n_60023), .B(n_17449), .C(n_60007), .D(n_17481), .Z
		(n_3330));
	notech_ao4 i_1869(.A(n_59971), .B(n_17417), .C(n_59679), .D(n_17625), .Z
		(n_3332));
	notech_ao4 i_1870(.A(n_59711), .B(n_17593), .C(n_59695), .D(n_17609), .Z
		(n_3333));
	notech_and4 i_1879(.A(n_3333), .B(n_3332), .C(n_3330), .D(n_3004), .Z(n_3335
		));
	notech_ao4 i_1871(.A(n_59743), .B(n_17561), .C(n_59727), .D(n_17577), .Z
		(n_3336));
	notech_ao4 i_1872(.A(n_60039), .B(n_17529), .C(n_59759), .D(n_17545), .Z
		(n_3337));
	notech_ao4 i_1873(.A(n_60071), .B(n_17497), .C(n_60055), .D(n_17513), .Z
		(n_3339));
	notech_ao4 i_1874(.A(n_59989), .B(n_17409), .C(n_60087), .D(n_17465), .Z
		(n_3340));
	notech_and4 i_1880(.A(n_3340), .B(n_3339), .C(n_3337), .D(n_3336), .Z(n_3342
		));
	notech_ao4 i_2054(.A(n_60027), .B(n_17461), .C(n_60011), .D(n_17493), .Z
		(n_3344));
	notech_ao4 i_2055(.A(n_59971), .B(n_17429), .C(n_59683), .D(n_17637), .Z
		(n_3346));
	notech_ao4 i_2056(.A(n_59715), .B(n_17605), .C(n_59699), .D(n_17621), .Z
		(n_3347));
	notech_and4 i_2065(.A(n_3347), .B(n_3346), .C(n_3344), .D(n_3020), .Z(n_3349
		));
	notech_ao4 i_2057(.A(n_59747), .B(n_17573), .C(n_59731), .D(n_17589), .Z
		(n_3350));
	notech_ao4 i_2058(.A(n_60043), .B(n_17541), .C(n_59763), .D(n_17557), .Z
		(n_3351));
	notech_ao4 i_2059(.A(n_60071), .B(n_17509), .C(n_60059), .D(n_17525), .Z
		(n_3353));
	notech_ao4 i_2060(.A(n_59989), .B(n_17415), .C(n_60087), .D(n_17477), .Z
		(n_3354));
	notech_and4 i_2066(.A(n_3354), .B(n_3353), .C(n_3351), .D(n_3350), .Z(n_3356
		));
	notech_ao4 i_2116(.A(n_60029), .B(n_17465), .C(n_60013), .D(n_17497), .Z
		(n_3358));
	notech_ao4 i_2117(.A(n_59975), .B(n_17433), .C(n_59685), .D(n_17641), .Z
		(n_3360));
	notech_ao4 i_2118(.A(n_59717), .B(n_17609), .C(n_59701), .D(n_17625), .Z
		(n_3361));
	notech_and4 i_2127(.A(n_3361), .B(n_3360), .C(n_3358), .D(n_3036), .Z(n_3363
		));
	notech_ao4 i_2119(.A(n_59749), .B(n_17577), .C(n_59733), .D(n_17593), .Z
		(n_3364));
	notech_ao4 i_2120(.A(n_60045), .B(n_17545), .C(n_59765), .D(n_17561), .Z
		(n_3365));
	notech_ao4 i_2121(.A(n_60075), .B(n_17513), .C(n_60061), .D(n_17529), .Z
		(n_3367));
	notech_ao4 i_2122(.A(n_59989), .B(n_17417), .C(n_60091), .D(n_17481), .Z
		(n_3368));
	notech_and4 i_2128(.A(n_3368), .B(n_3367), .C(n_3365), .D(n_3364), .Z(n_3370
		));
	notech_ao4 i_2302(.A(n_60029), .B(n_17477), .C(n_60013), .D(n_17509), .Z
		(n_3372));
	notech_ao4 i_2303(.A(n_59975), .B(n_17445), .C(n_59685), .D(n_17653), .Z
		(n_3374));
	notech_ao4 i_2304(.A(n_59717), .B(n_17621), .C(n_59701), .D(n_17637), .Z
		(n_3375));
	notech_and4 i_2313(.A(n_3375), .B(n_3374), .C(n_3372), .D(n_3052), .Z(n_3377
		));
	notech_ao4 i_2305(.A(n_59749), .B(n_17589), .C(n_59733), .D(n_17605), .Z
		(n_3378));
	notech_ao4 i_2306(.A(n_60045), .B(n_17557), .C(n_59765), .D(n_17573), .Z
		(n_3379));
	notech_ao4 i_2307(.A(n_60077), .B(n_17525), .C(n_60061), .D(n_17541), .Z
		(n_3381));
	notech_ao4 i_2308(.A(n_59994), .B(n_17429), .C(n_60093), .D(n_17493), .Z
		(n_3382));
	notech_and4 i_2314(.A(n_3382), .B(n_3381), .C(n_3379), .D(n_3378), .Z(n_3384
		));
	notech_ao4 i_2364(.A(n_60029), .B(n_17481), .C(n_60013), .D(n_17513), .Z
		(n_3386));
	notech_ao4 i_2365(.A(n_59978), .B(n_17449), .C(n_59685), .D(n_17657), .Z
		(n_3388));
	notech_ao4 i_2366(.A(n_59717), .B(n_17625), .C(n_59701), .D(n_17641), .Z
		(n_3389));
	notech_and4 i_2375(.A(n_3389), .B(n_3388), .C(n_3386), .D(n_3068), .Z(n_3391
		));
	notech_ao4 i_2367(.A(n_59749), .B(n_17593), .C(n_59733), .D(n_17609), .Z
		(n_3392));
	notech_ao4 i_2368(.A(n_60045), .B(n_17561), .C(n_59765), .D(n_17577), .Z
		(n_3393));
	notech_ao4 i_2369(.A(n_60077), .B(n_17529), .C(n_60061), .D(n_17545), .Z
		(n_3395));
	notech_ao4 i_2370(.A(n_59996), .B(n_17433), .C(n_60093), .D(n_17497), .Z
		(n_3396));
	notech_and4 i_2376(.A(n_3396), .B(n_3395), .C(n_3393), .D(n_3392), .Z(n_3398
		));
	notech_ao4 i_227159(.A(n_1129), .B(addrshft[1]), .C(n_113256518), .D(n_113356519
		), .Z(valid_len_1101034));
	notech_ao4 i_327160(.A(n_3400), .B(addrshft[2]), .C(n_113256518), .D(n_1123
		), .Z(valid_len_2101033));
	notech_ao4 i_427161(.A(n_1129), .B(addrshft[3]), .C(n_113256518), .D(n_1114
		), .Z(valid_len_3101032));
	notech_ao3 i_627163(.A(n_61430), .B(addrshft[5]), .C(wptr[0]), .Z(valid_len
		[5]));
	notech_ao4 i_128333647(.A(n_59864), .B(n_17366), .C(n_59851), .D(n_17374
		), .Z(n_2544));
	notech_nand2 i_331122(.A(n_61430), .B(n_17300), .Z(n_3400));
	notech_ao4 i_128133649(.A(n_59978), .B(n_17350), .C(n_59959), .D(n_17358
		), .Z(n_2542));
	notech_ao4 i_125833672(.A(n_2006), .B(n_17457), .C(n_2005), .D(n_17441),
		 .Z(n_2539));
	notech_ao4 i_125733673(.A(n_2003), .B(n_17425), .C(n_2002), .D(n_17489),
		 .Z(n_2538));
	notech_and3 i_126033670(.A(n_2535), .B(n_2534), .C(n_1782), .Z(n_2537)
		);
	notech_ao4 i_125433676(.A(n_1998), .B(n_17405), .C(n_1997), .D(n_17389),
		 .Z(n_2535));
	notech_ao4 i_125333677(.A(n_1995), .B(n_17381), .C(n_1994), .D(n_17397),
		 .Z(n_2534));
	notech_and4 i_126233668(.A(n_2528), .B(n_2530), .C(n_2532), .D(n_1769), 
		.Z(n_2533));
	notech_ao4 i_125933671(.A(n_1991), .B(n_17413), .C(n_1990), .D(n_17473),
		 .Z(n_2532));
	notech_ao4 i_125233678(.A(n_1986), .B(n_17365), .C(n_1985), .D(n_17373),
		 .Z(n_2530));
	notech_ao4 i_125033680(.A(n_59978), .B(n_17349), .C(n_59959), .D(n_17357
		), .Z(n_2528));
	notech_ao4 i_122733703(.A(n_2006), .B(n_17455), .C(n_2005), .D(n_17439),
		 .Z(n_2525));
	notech_ao4 i_122633704(.A(n_2003), .B(n_17423), .C(n_2002), .D(n_17487),
		 .Z(n_2524));
	notech_and3 i_122933701(.A(n_2521), .B(n_2520), .C(n_1766), .Z(n_2523)
		);
	notech_ao4 i_122333707(.A(n_1998), .B(n_17404), .C(n_1997), .D(n_17388),
		 .Z(n_2521));
	notech_ao4 i_122233708(.A(n_1995), .B(n_17380), .C(n_1994), .D(n_17396),
		 .Z(n_2520));
	notech_and4 i_123133699(.A(n_2514), .B(n_2516), .C(n_2518), .D(n_1753), 
		.Z(n_2519));
	notech_ao4 i_122833702(.A(n_1991), .B(n_17412), .C(n_1990), .D(n_17471),
		 .Z(n_2518));
	notech_ao4 i_122133709(.A(n_1986), .B(n_17364), .C(n_1985), .D(n_17372),
		 .Z(n_2516));
	notech_ao4 i_121933711(.A(n_59978), .B(n_17348), .C(n_59959), .D(n_17356
		), .Z(n_2514));
	notech_ao4 i_119633734(.A(n_2006), .B(n_17453), .C(n_2005), .D(n_17437),
		 .Z(n_2511));
	notech_ao4 i_119533735(.A(n_2003), .B(n_17421), .C(n_2002), .D(n_17485),
		 .Z(n_2510));
	notech_and3 i_119833732(.A(n_2507), .B(n_2506), .C(n_1750), .Z(n_2509)
		);
	notech_ao4 i_119233738(.A(n_1998), .B(n_17403), .C(n_1997), .D(n_17387),
		 .Z(n_2507));
	notech_ao4 i_119133739(.A(n_1995), .B(n_17379), .C(n_1994), .D(n_17395),
		 .Z(n_2506));
	notech_and4 i_120033730(.A(n_2500), .B(n_2502), .C(n_2504), .D(n_1737), 
		.Z(n_2505));
	notech_ao4 i_119733733(.A(n_1991), .B(n_17411), .C(n_1990), .D(n_17469),
		 .Z(n_2504));
	notech_ao4 i_119033740(.A(n_1986), .B(n_17363), .C(n_1985), .D(n_17371),
		 .Z(n_2502));
	notech_ao4 i_118833742(.A(n_59978), .B(n_17347), .C(n_59996), .D(n_17339
		), .Z(n_2500));
	notech_ao4 i_116533765(.A(n_2006), .B(n_17451), .C(n_2005), .D(n_17435),
		 .Z(n_2497));
	notech_ao4 i_116433766(.A(n_2003), .B(n_17418), .C(n_2002), .D(n_17483),
		 .Z(n_2496));
	notech_and3 i_116733763(.A(n_2493), .B(n_2492), .C(n_1734), .Z(n_2495)
		);
	notech_ao4 i_116133769(.A(n_1998), .B(n_17402), .C(n_1997), .D(n_17386),
		 .Z(n_2493));
	notech_ao4 i_116033770(.A(n_1995), .B(n_17378), .C(n_1994), .D(n_17394),
		 .Z(n_2492));
	notech_and4 i_116933761(.A(n_2486), .B(n_2488), .C(n_2490), .D(n_1721), 
		.Z(n_2491));
	notech_ao4 i_116633764(.A(n_1991), .B(n_17410), .C(n_1990), .D(n_17467),
		 .Z(n_2490));
	notech_ao4 i_115933771(.A(n_1986), .B(n_17362), .C(n_1985), .D(n_17370),
		 .Z(n_2488));
	notech_ao4 i_115733773(.A(n_59978), .B(n_17346), .C(n_59959), .D(n_17354
		), .Z(n_2486));
	notech_ao4 i_113433796(.A(n_2006), .B(n_17449), .C(n_2005), .D(n_17433),
		 .Z(n_2483));
	notech_ao4 i_113333797(.A(n_2003), .B(n_17417), .C(n_2002), .D(n_17481),
		 .Z(n_2482));
	notech_and3 i_113633794(.A(n_2479), .B(n_2478), .C(n_1718), .Z(n_2481)
		);
	notech_ao4 i_113033800(.A(n_1998), .B(n_17401), .C(n_1997), .D(n_17385),
		 .Z(n_2479));
	notech_ao4 i_112933801(.A(n_1995), .B(n_17377), .C(n_1994), .D(n_17393),
		 .Z(n_2478));
	notech_and4 i_113833792(.A(n_2472), .B(n_2474), .C(n_2476), .D(n_1705), 
		.Z(n_2477));
	notech_ao4 i_113533795(.A(n_1991), .B(n_17409), .C(n_1990), .D(n_17465),
		 .Z(n_2476));
	notech_ao4 i_112833802(.A(n_1986), .B(n_17361), .C(n_1985), .D(n_17369),
		 .Z(n_2474));
	notech_ao4 i_112633804(.A(n_59978), .B(n_17345), .C(n_59959), .D(n_17353
		), .Z(n_2472));
	notech_ao4 i_110333827(.A(n_2006), .B(n_17445), .C(n_2005), .D(n_17429),
		 .Z(n_2469));
	notech_ao4 i_110233828(.A(n_2003), .B(n_17415), .C(n_2002), .D(n_17477),
		 .Z(n_2468));
	notech_and3 i_110533825(.A(n_2465), .B(n_2464), .C(n_1702), .Z(n_2467)
		);
	notech_ao4 i_109933831(.A(n_1998), .B(n_17399), .C(n_1997), .D(n_17383),
		 .Z(n_2465));
	notech_ao4 i_109833832(.A(n_1995), .B(n_17375), .C(n_1994), .D(n_17391),
		 .Z(n_2464));
	notech_and4 i_110733823(.A(n_2458), .B(n_2460), .C(n_2462), .D(n_1689), 
		.Z(n_2463));
	notech_ao4 i_110433826(.A(n_1991), .B(n_17407), .C(n_1990), .D(n_17461),
		 .Z(n_2462));
	notech_ao4 i_109733833(.A(n_1986), .B(n_17359), .C(n_1985), .D(n_17367),
		 .Z(n_2460));
	notech_ao4 i_109533835(.A(n_59978), .B(n_17343), .C(n_59959), .D(n_17351
		), .Z(n_2458));
	notech_ao4 i_107233858(.A(n_2006), .B(n_17443), .C(n_2005), .D(n_17427),
		 .Z(n_2455));
	notech_ao4 i_107133859(.A(n_2003), .B(n_17414), .C(n_2002), .D(n_17475),
		 .Z(n_2454));
	notech_and3 i_107433856(.A(n_2451), .B(n_2450), .C(n_1686), .Z(n_2453)
		);
	notech_ao4 i_106833862(.A(n_1998), .B(n_17398), .C(n_1997), .D(n_17382),
		 .Z(n_2451));
	notech_ao4 i_106733863(.A(n_1995), .B(n_17374), .C(n_1994), .D(n_17390),
		 .Z(n_2450));
	notech_and4 i_107633854(.A(n_2444), .B(n_2446), .C(n_2448), .D(n_1673), 
		.Z(n_2449));
	notech_ao4 i_107333857(.A(n_1991), .B(n_17406), .C(n_1990), .D(n_17459),
		 .Z(n_2448));
	notech_ao4 i_106633864(.A(n_1986), .B(n_17358), .C(n_1985), .D(n_17366),
		 .Z(n_2446));
	notech_ao4 i_106433866(.A(n_59978), .B(n_17342), .C(n_59959), .D(n_17350
		), .Z(n_2444));
	notech_ao4 i_104133889(.A(n_2006), .B(n_17441), .C(n_2005), .D(n_17425),
		 .Z(n_2441));
	notech_ao4 i_104033890(.A(n_2003), .B(n_17413), .C(n_2002), .D(n_17473),
		 .Z(n_2440));
	notech_and3 i_104333887(.A(n_2437), .B(n_2436), .C(n_1670), .Z(n_2439)
		);
	notech_ao4 i_103733893(.A(n_1998), .B(n_17397), .C(n_1997), .D(n_17381),
		 .Z(n_2437));
	notech_ao4 i_103633894(.A(n_1995), .B(n_17373), .C(n_1994), .D(n_17389),
		 .Z(n_2436));
	notech_and4 i_104533885(.A(n_2430), .B(n_2432), .C(n_2434), .D(n_1657), 
		.Z(n_2435));
	notech_ao4 i_104233888(.A(n_1991), .B(n_17405), .C(n_1990), .D(n_17457),
		 .Z(n_2434));
	notech_ao4 i_103533895(.A(n_1986), .B(n_17357), .C(n_1985), .D(n_17365),
		 .Z(n_2432));
	notech_ao4 i_103333897(.A(n_59978), .B(n_17341), .C(n_59959), .D(n_17349
		), .Z(n_2430));
	notech_ao4 i_101033920(.A(n_2006), .B(n_17439), .C(n_2005), .D(n_17423),
		 .Z(n_2427));
	notech_ao4 i_100933921(.A(n_2003), .B(n_17412), .C(n_2002), .D(n_17471),
		 .Z(n_2426));
	notech_and3 i_101233918(.A(n_2423), .B(n_2422), .C(n_1654), .Z(n_2425)
		);
	notech_ao4 i_100633924(.A(n_1998), .B(n_17396), .C(n_1997), .D(n_17380),
		 .Z(n_2423));
	notech_ao4 i_100533925(.A(n_1995), .B(n_17372), .C(n_1994), .D(n_17388),
		 .Z(n_2422));
	notech_and4 i_101433916(.A(n_2416), .B(n_2418), .C(n_2420), .D(n_1641), 
		.Z(n_2421));
	notech_ao4 i_101133919(.A(n_1991), .B(n_17404), .C(n_1990), .D(n_17455),
		 .Z(n_2420));
	notech_ao4 i_100433926(.A(n_1986), .B(n_17356), .C(n_1985), .D(n_17364),
		 .Z(n_2418));
	notech_ao4 i_100233928(.A(n_59978), .B(n_17340), .C(n_59959), .D(n_17348
		), .Z(n_2416));
	notech_ao4 i_97933951(.A(n_2006), .B(n_17437), .C(n_2005), .D(n_17421), 
		.Z(n_2413));
	notech_ao4 i_97833952(.A(n_2003), .B(n_17411), .C(n_2002), .D(n_17469), 
		.Z(n_2412));
	notech_and3 i_98133949(.A(n_2409), .B(n_2408), .C(n_1638), .Z(n_2411));
	notech_ao4 i_97533955(.A(n_1998), .B(n_17395), .C(n_1997), .D(n_17379), 
		.Z(n_2409));
	notech_ao4 i_97433956(.A(n_1995), .B(n_17371), .C(n_1994), .D(n_17387), 
		.Z(n_2408));
	notech_and4 i_98333947(.A(n_2402), .B(n_2404), .C(n_2406), .D(n_1625), .Z
		(n_2407));
	notech_ao4 i_98033950(.A(n_1991), .B(n_17403), .C(n_1990), .D(n_17453), 
		.Z(n_2406));
	notech_ao4 i_97333957(.A(n_1986), .B(n_17355), .C(n_1985), .D(n_17363), 
		.Z(n_2404));
	notech_ao4 i_97133959(.A(n_59959), .B(n_17347), .C(n_59978), .D(n_17339)
		, .Z(n_2402));
	notech_ao4 i_94833982(.A(n_2006), .B(n_17435), .C(n_2005), .D(n_17418), 
		.Z(n_2399));
	notech_ao4 i_94733983(.A(n_2003), .B(n_17410), .C(n_2002), .D(n_17467), 
		.Z(n_2398));
	notech_and3 i_95033980(.A(n_2395), .B(n_2394), .C(n_1622), .Z(n_2397));
	notech_ao4 i_94433986(.A(n_1998), .B(n_17394), .C(n_1997), .D(n_17378), 
		.Z(n_2395));
	notech_ao4 i_94333987(.A(n_1995), .B(n_17370), .C(n_1994), .D(n_17386), 
		.Z(n_2394));
	notech_and4 i_95233978(.A(n_2388), .B(n_2390), .C(n_2392), .D(n_1609), .Z
		(n_2393));
	notech_ao4 i_94933981(.A(n_1991), .B(n_17402), .C(n_1990), .D(n_17451), 
		.Z(n_2392));
	notech_ao4 i_94233988(.A(n_1986), .B(n_17354), .C(n_1985), .D(n_17362), 
		.Z(n_2390));
	notech_ao4 i_94033990(.A(n_59978), .B(n_17338), .C(n_59959), .D(n_17346)
		, .Z(n_2388));
	notech_ao4 i_91734013(.A(n_2006), .B(n_17433), .C(n_2005), .D(n_17417), 
		.Z(n_2385));
	notech_ao4 i_91634014(.A(n_2003), .B(n_17409), .C(n_2002), .D(n_17465), 
		.Z(n_2384));
	notech_and3 i_91934011(.A(n_2381), .B(n_2380), .C(n_1606), .Z(n_2383));
	notech_ao4 i_91334017(.A(n_1998), .B(n_17393), .C(n_1997), .D(n_17377), 
		.Z(n_2381));
	notech_ao4 i_91234018(.A(n_1995), .B(n_17369), .C(n_1994), .D(n_17385), 
		.Z(n_2380));
	notech_and4 i_92134009(.A(n_2374), .B(n_2376), .C(n_2378), .D(n_1593), .Z
		(n_2379));
	notech_ao4 i_91834012(.A(n_1991), .B(n_17401), .C(n_1990), .D(n_17449), 
		.Z(n_2378));
	notech_ao4 i_91134019(.A(n_1986), .B(n_17353), .C(n_1985), .D(n_17361), 
		.Z(n_2376));
	notech_ao4 i_90934021(.A(n_59978), .B(n_17337), .C(n_59959), .D(n_17345)
		, .Z(n_2374));
	notech_ao4 i_88634044(.A(n_2006), .B(n_17429), .C(n_2005), .D(n_17415), 
		.Z(n_2371));
	notech_ao4 i_88534045(.A(n_2003), .B(n_17407), .C(n_2002), .D(n_17461), 
		.Z(n_2370));
	notech_and3 i_88834042(.A(n_2367), .B(n_2366), .C(n_1590), .Z(n_2369));
	notech_ao4 i_88234048(.A(n_1998), .B(n_17391), .C(n_1997), .D(n_17375), 
		.Z(n_2367));
	notech_ao4 i_88134049(.A(n_1995), .B(n_17367), .C(n_1994), .D(n_17383), 
		.Z(n_2366));
	notech_and4 i_89034040(.A(n_2360), .B(n_2362), .C(n_2364), .D(n_1577), .Z
		(n_2365));
	notech_ao4 i_88734043(.A(n_1991), .B(n_17399), .C(n_1990), .D(n_17445), 
		.Z(n_2364));
	notech_ao4 i_88034050(.A(n_1986), .B(n_17351), .C(n_1985), .D(n_17359), 
		.Z(n_2362));
	notech_ao4 i_87834052(.A(n_59978), .B(n_17335), .C(n_59959), .D(n_17343)
		, .Z(n_2360));
	notech_ao4 i_85534075(.A(n_59916), .B(n_17427), .C(n_59903), .D(n_17414)
		, .Z(n_2357));
	notech_ao4 i_85434076(.A(n_59890), .B(n_17406), .C(n_59877), .D(n_17459)
		, .Z(n_2356));
	notech_and3 i_85734073(.A(n_2353), .B(n_2352), .C(n_1574), .Z(n_2355));
	notech_ao4 i_85134079(.A(n_59812), .B(n_17390), .C(n_59799), .D(n_17374)
		, .Z(n_2353));
	notech_ao4 i_85034080(.A(n_59786), .B(n_17366), .C(n_59773), .D(n_17382)
		, .Z(n_2352));
	notech_and4 i_85934071(.A(n_2346), .B(n_2348), .C(n_2350), .D(n_1561), .Z
		(n_2351));
	notech_ao4 i_85634074(.A(n_59838), .B(n_17398), .C(n_59825), .D(n_17443)
		, .Z(n_2350));
	notech_ao4 i_84934081(.A(n_59864), .B(n_17350), .C(n_59851), .D(n_17358)
		, .Z(n_2348));
	notech_ao4 i_84734083(.A(n_59978), .B(n_17334), .C(n_59959), .D(n_17342)
		, .Z(n_2346));
	notech_ao4 i_82434106(.A(n_59912), .B(n_17425), .C(n_59899), .D(n_17413)
		, .Z(n_2343));
	notech_ao4 i_82334107(.A(n_59886), .B(n_17405), .C(n_59873), .D(n_17457)
		, .Z(n_2342));
	notech_and3 i_82634104(.A(n_2339), .B(n_2338), .C(n_1558), .Z(n_2341));
	notech_ao4 i_82034110(.A(n_59808), .B(n_17389), .C(n_59795), .D(n_17373)
		, .Z(n_2339));
	notech_ao4 i_81934111(.A(n_59782), .B(n_17365), .C(n_59769), .D(n_17381)
		, .Z(n_2338));
	notech_and4 i_82834102(.A(n_2332), .B(n_2334), .C(n_2336), .D(n_1545), .Z
		(n_2337));
	notech_ao4 i_82534105(.A(n_59834), .B(n_17397), .C(n_59821), .D(n_17441)
		, .Z(n_2336));
	notech_ao4 i_81834112(.A(n_59860), .B(n_17349), .C(n_59847), .D(n_17357)
		, .Z(n_2334));
	notech_ao4 i_81634114(.A(n_59976), .B(n_17333), .C(n_59957), .D(n_17341)
		, .Z(n_2332));
	notech_ao4 i_79334137(.A(n_59912), .B(n_17423), .C(n_59899), .D(n_17412)
		, .Z(n_2329));
	notech_ao4 i_79234138(.A(n_59886), .B(n_17404), .C(n_59873), .D(n_17455)
		, .Z(n_2328));
	notech_and3 i_79534135(.A(n_2325), .B(n_2324), .C(n_1542), .Z(n_2327));
	notech_ao4 i_78934141(.A(n_59808), .B(n_17388), .C(n_59795), .D(n_17372)
		, .Z(n_2325));
	notech_ao4 i_78834142(.A(n_59782), .B(n_17364), .C(n_59769), .D(n_17380)
		, .Z(n_2324));
	notech_and4 i_79734133(.A(n_2318), .B(n_2320), .C(n_2322), .D(n_1529), .Z
		(n_2323));
	notech_ao4 i_79434136(.A(n_59834), .B(n_17396), .C(n_59821), .D(n_17439)
		, .Z(n_2322));
	notech_ao4 i_78734143(.A(n_59860), .B(n_17348), .C(n_59847), .D(n_17356)
		, .Z(n_2320));
	notech_ao4 i_78534145(.A(n_59976), .B(n_17332), .C(n_59957), .D(n_17340)
		, .Z(n_2318));
	notech_ao4 i_76234168(.A(n_59912), .B(n_17421), .C(n_59899), .D(n_17411)
		, .Z(n_2315));
	notech_ao4 i_76134169(.A(n_59886), .B(n_17403), .C(n_59873), .D(n_17453)
		, .Z(n_2314));
	notech_and3 i_76434166(.A(n_2311), .B(n_2310), .C(n_1526), .Z(n_2313));
	notech_ao4 i_75834172(.A(n_59808), .B(n_17387), .C(n_59795), .D(n_17371)
		, .Z(n_2311));
	notech_ao4 i_75734173(.A(n_59782), .B(n_17363), .C(n_59769), .D(n_17379)
		, .Z(n_2310));
	notech_and4 i_76634164(.A(n_2304), .B(n_2306), .C(n_2308), .D(n_1513), .Z
		(n_2309));
	notech_ao4 i_76334167(.A(n_59834), .B(n_17395), .C(n_59821), .D(n_17437)
		, .Z(n_2308));
	notech_ao4 i_75634174(.A(n_59860), .B(n_17347), .C(n_59847), .D(n_17355)
		, .Z(n_2306));
	notech_ao4 i_75434176(.A(n_59976), .B(n_17331), .C(n_59957), .D(n_17339)
		, .Z(n_2304));
	notech_ao4 i_73134199(.A(n_59912), .B(n_17418), .C(n_59899), .D(n_17410)
		, .Z(n_2301));
	notech_ao4 i_73034200(.A(n_59886), .B(n_17402), .C(n_59873), .D(n_17451)
		, .Z(n_2300));
	notech_and3 i_73334197(.A(n_2297), .B(n_2296), .C(n_1510), .Z(n_2299));
	notech_ao4 i_72734203(.A(n_59808), .B(n_17386), .C(n_59795), .D(n_17370)
		, .Z(n_2297));
	notech_ao4 i_72634204(.A(n_59782), .B(n_17362), .C(n_59769), .D(n_17378)
		, .Z(n_2296));
	notech_and4 i_73534195(.A(n_2290), .B(n_2292), .C(n_2294), .D(n_1497), .Z
		(n_2295));
	notech_ao4 i_73234198(.A(n_59834), .B(n_17394), .C(n_59821), .D(n_17435)
		, .Z(n_2294));
	notech_ao4 i_72534205(.A(n_59860), .B(n_17346), .C(n_59847), .D(n_17354)
		, .Z(n_2292));
	notech_ao4 i_72334207(.A(n_59976), .B(n_17330), .C(n_59957), .D(n_17338)
		, .Z(n_2290));
	notech_ao4 i_70034230(.A(n_59912), .B(n_17417), .C(n_59899), .D(n_17409)
		, .Z(n_2287));
	notech_ao4 i_69934231(.A(n_59886), .B(n_17401), .C(n_59873), .D(n_17449)
		, .Z(n_2286));
	notech_and3 i_70234228(.A(n_2283), .B(n_2282), .C(n_1494), .Z(n_2285));
	notech_ao4 i_69634234(.A(n_59808), .B(n_17385), .C(n_59795), .D(n_17369)
		, .Z(n_2283));
	notech_ao4 i_69534235(.A(n_59782), .B(n_17361), .C(n_59769), .D(n_17377)
		, .Z(n_2282));
	notech_and4 i_70434226(.A(n_2276), .B(n_2278), .C(n_2280), .D(n_1481), .Z
		(n_2281));
	notech_ao4 i_70134229(.A(n_59834), .B(n_17393), .C(n_59821), .D(n_17433)
		, .Z(n_2280));
	notech_ao4 i_69434236(.A(n_59860), .B(n_17345), .C(n_59847), .D(n_17353)
		, .Z(n_2278));
	notech_ao4 i_69234238(.A(n_59976), .B(n_17329), .C(n_59957), .D(n_17337)
		, .Z(n_2276));
	notech_ao4 i_66934261(.A(n_59912), .B(n_17416), .C(n_59899), .D(n_17408)
		, .Z(n_2273));
	notech_ao4 i_66834262(.A(n_59886), .B(n_17400), .C(n_59873), .D(n_17447)
		, .Z(n_2272));
	notech_and3 i_67134259(.A(n_2269), .B(n_2268), .C(n_1478), .Z(n_2271));
	notech_ao4 i_66534265(.A(n_59808), .B(n_17384), .C(n_59795), .D(n_17368)
		, .Z(n_2269));
	notech_ao4 i_66434266(.A(n_59782), .B(n_17360), .C(n_59769), .D(n_17376)
		, .Z(n_2268));
	notech_and4 i_67334257(.A(n_2262), .B(n_2264), .C(n_2266), .D(n_1465), .Z
		(n_2267));
	notech_ao4 i_67034260(.A(n_59834), .B(n_17392), .C(n_59821), .D(n_17431)
		, .Z(n_2266));
	notech_ao4 i_66334267(.A(n_59860), .B(n_17344), .C(n_59847), .D(n_17352)
		, .Z(n_2264));
	notech_ao4 i_66134269(.A(n_59976), .B(n_17328), .C(n_59957), .D(n_17336)
		, .Z(n_2262));
	notech_ao4 i_63834292(.A(n_59912), .B(n_17415), .C(n_59899), .D(n_17407)
		, .Z(n_2259));
	notech_ao4 i_63734293(.A(n_59886), .B(n_17399), .C(n_59873), .D(n_17445)
		, .Z(n_2258));
	notech_and3 i_64034290(.A(n_2255), .B(n_2254), .C(n_1462), .Z(n_2257));
	notech_ao4 i_63434296(.A(n_59808), .B(n_17383), .C(n_59795), .D(n_17367)
		, .Z(n_2255));
	notech_ao4 i_63334297(.A(n_59782), .B(n_17359), .C(n_59769), .D(n_17375)
		, .Z(n_2254));
	notech_and4 i_64234288(.A(n_2248), .B(n_2250), .C(n_2252), .D(n_1449), .Z
		(n_2253));
	notech_ao4 i_63934291(.A(n_59834), .B(n_17391), .C(n_59821), .D(n_17429)
		, .Z(n_2252));
	notech_ao4 i_63234298(.A(n_59860), .B(n_17343), .C(n_59847), .D(n_17351)
		, .Z(n_2250));
	notech_ao4 i_63034300(.A(n_59976), .B(n_17327), .C(n_59957), .D(n_17335)
		, .Z(n_2248));
	notech_ao4 i_60734323(.A(n_59912), .B(n_17414), .C(n_59899), .D(n_17406)
		, .Z(n_2245));
	notech_ao4 i_60634324(.A(n_59886), .B(n_17398), .C(n_59873), .D(n_17443)
		, .Z(n_2244));
	notech_and3 i_60934321(.A(n_2241), .B(n_2240), .C(n_1446), .Z(n_2243));
	notech_ao4 i_60334327(.A(n_59808), .B(n_17382), .C(n_59795), .D(n_17366)
		, .Z(n_2241));
	notech_ao4 i_60234328(.A(n_59782), .B(n_17358), .C(n_59769), .D(n_17374)
		, .Z(n_2240));
	notech_and4 i_61134319(.A(n_2234), .B(n_2236), .C(n_2238), .D(n_1433), .Z
		(n_2239));
	notech_ao4 i_60834322(.A(n_59834), .B(n_17390), .C(n_59821), .D(n_17427)
		, .Z(n_2238));
	notech_ao4 i_60134329(.A(n_59860), .B(n_17342), .C(n_59847), .D(n_17350)
		, .Z(n_2236));
	notech_ao4 i_59934331(.A(n_59976), .B(n_17326), .C(n_59957), .D(n_17334)
		, .Z(n_2234));
	notech_ao4 i_57634354(.A(n_59912), .B(n_17413), .C(n_59899), .D(n_17405)
		, .Z(n_2231));
	notech_ao4 i_57534355(.A(n_59886), .B(n_17397), .C(n_59873), .D(n_17441)
		, .Z(n_2230));
	notech_and3 i_57834352(.A(n_2227), .B(n_2226), .C(n_1430), .Z(n_2229));
	notech_ao4 i_57234358(.A(n_59808), .B(n_17381), .C(n_59795), .D(n_17365)
		, .Z(n_2227));
	notech_ao4 i_57134359(.A(n_59782), .B(n_17357), .C(n_59769), .D(n_17373)
		, .Z(n_2226));
	notech_and4 i_58034350(.A(n_2220), .B(n_2222), .C(n_2224), .D(n_1417), .Z
		(n_2225));
	notech_ao4 i_57734353(.A(n_59834), .B(n_17389), .C(n_59821), .D(n_17425)
		, .Z(n_2224));
	notech_ao4 i_57034360(.A(n_59860), .B(n_17341), .C(n_59847), .D(n_17349)
		, .Z(n_2222));
	notech_ao4 i_56834362(.A(n_59976), .B(n_17325), .C(n_59957), .D(n_17333)
		, .Z(n_2220));
	notech_ao4 i_54534385(.A(n_59912), .B(n_17412), .C(n_59899), .D(n_17404)
		, .Z(n_2217));
	notech_ao4 i_54434386(.A(n_59886), .B(n_17396), .C(n_59873), .D(n_17439)
		, .Z(n_2216));
	notech_and3 i_54734383(.A(n_2213), .B(n_2212), .C(n_1414), .Z(n_2215));
	notech_ao4 i_54134389(.A(n_59808), .B(n_17380), .C(n_59795), .D(n_17364)
		, .Z(n_2213));
	notech_ao4 i_54034390(.A(n_59782), .B(n_17356), .C(n_59769), .D(n_17372)
		, .Z(n_2212));
	notech_and4 i_54934381(.A(n_2206), .B(n_2208), .C(n_2210), .D(n_1401), .Z
		(n_2211));
	notech_ao4 i_54634384(.A(n_59834), .B(n_17388), .C(n_59821), .D(n_17423)
		, .Z(n_2210));
	notech_ao4 i_53934391(.A(n_59860), .B(n_17340), .C(n_59847), .D(n_17348)
		, .Z(n_2208));
	notech_ao4 i_53734393(.A(n_59976), .B(n_17324), .C(n_59957), .D(n_17332)
		, .Z(n_2206));
	notech_ao4 i_51434416(.A(n_59912), .B(n_17411), .C(n_59899), .D(n_17403)
		, .Z(n_2203));
	notech_ao4 i_51334417(.A(n_59886), .B(n_17395), .C(n_59873), .D(n_17437)
		, .Z(n_2202));
	notech_and3 i_51634414(.A(n_2199), .B(n_2198), .C(n_1398), .Z(n_2201));
	notech_ao4 i_51034420(.A(n_59808), .B(n_17379), .C(n_59795), .D(n_17363)
		, .Z(n_2199));
	notech_ao4 i_50934421(.A(n_59782), .B(n_17355), .C(n_59769), .D(n_17371)
		, .Z(n_2198));
	notech_and4 i_51834412(.A(n_2192), .B(n_2194), .C(n_2196), .D(n_1385), .Z
		(n_2197));
	notech_ao4 i_51534415(.A(n_59834), .B(n_17387), .C(n_59821), .D(n_17421)
		, .Z(n_2196));
	notech_ao4 i_50834422(.A(n_59860), .B(n_17339), .C(n_59847), .D(n_17347)
		, .Z(n_2194));
	notech_ao4 i_50634424(.A(n_59959), .B(n_17331), .C(n_59996), .D(n_17315)
		, .Z(n_2192));
	notech_ao4 i_48334447(.A(n_17410), .B(n_59912), .C(n_17402), .D(n_59899)
		, .Z(n_2189));
	notech_ao4 i_48234448(.A(n_17394), .B(n_59886), .C(n_17435), .D(n_59873)
		, .Z(n_2188));
	notech_and3 i_48534445(.A(n_2185), .B(n_2184), .C(n_1382), .Z(n_2187));
	notech_ao4 i_47934451(.A(n_17378), .B(n_59808), .C(n_17362), .D(n_59795)
		, .Z(n_2185));
	notech_ao4 i_47834452(.A(n_17354), .B(n_59782), .C(n_17370), .D(n_59769)
		, .Z(n_2184));
	notech_and4 i_48734443(.A(n_2178), .B(n_2180), .C(n_2182), .D(n_1369), .Z
		(n_2183));
	notech_ao4 i_48434446(.A(n_17386), .B(n_59834), .C(n_17418), .D(n_59821)
		, .Z(n_2182));
	notech_ao4 i_47734453(.A(n_17338), .B(n_59860), .C(n_17346), .D(n_59847)
		, .Z(n_2180));
	notech_ao4 i_47534455(.A(n_59978), .B(n_17322), .C(n_59959), .D(n_17330)
		, .Z(n_2178));
	notech_ao4 i_45234478(.A(n_59912), .B(n_17408), .C(n_59899), .D(n_17400)
		, .Z(n_2175));
	notech_ao4 i_45134479(.A(n_59886), .B(n_17392), .C(n_59873), .D(n_17431)
		, .Z(n_2174));
	notech_and3 i_45434476(.A(n_2171), .B(n_2170), .C(n_1366), .Z(n_2173));
	notech_ao4 i_44834482(.A(n_59808), .B(n_17376), .C(n_59795), .D(n_17360)
		, .Z(n_2171));
	notech_ao4 i_44734483(.A(n_59782), .B(n_17352), .C(n_59769), .D(n_17368)
		, .Z(n_2170));
	notech_and4 i_45634474(.A(n_2164), .B(n_2166), .C(n_2168), .D(n_1353), .Z
		(n_2169));
	notech_ao4 i_45334477(.A(n_59834), .B(n_17384), .C(n_59821), .D(n_17416)
		, .Z(n_2168));
	notech_ao4 i_44634484(.A(n_59860), .B(n_17336), .C(n_59847), .D(n_17344)
		, .Z(n_2166));
	notech_ao4 i_44434486(.A(n_59978), .B(n_17320), .C(n_59957), .D(n_17328)
		, .Z(n_2164));
	notech_ao4 i_42134509(.A(n_59916), .B(n_17407), .C(n_59903), .D(n_17399)
		, .Z(n_2161));
	notech_ao4 i_42034510(.A(n_59890), .B(n_17391), .C(n_59877), .D(n_17429)
		, .Z(n_2160));
	notech_and3 i_42334507(.A(n_2157), .B(n_2156), .C(n_1350), .Z(n_2159));
	notech_ao4 i_41734513(.A(n_59812), .B(n_17375), .C(n_59799), .D(n_17359)
		, .Z(n_2157));
	notech_ao4 i_41634514(.A(n_59786), .B(n_17351), .C(n_59773), .D(n_17367)
		, .Z(n_2156));
	notech_and4 i_42534505(.A(n_2150), .B(n_2152), .C(n_2154), .D(n_1337), .Z
		(n_2155));
	notech_ao4 i_42234508(.A(n_59838), .B(n_17383), .C(n_59825), .D(n_17415)
		, .Z(n_2154));
	notech_ao4 i_41534515(.A(n_59864), .B(n_17335), .C(n_59851), .D(n_17343)
		, .Z(n_2152));
	notech_ao4 i_41334517(.A(n_59976), .B(n_17319), .C(n_59957), .D(n_17327)
		, .Z(n_2150));
	notech_ao4 i_39034540(.A(n_59916), .B(n_17406), .C(n_59903), .D(n_17398)
		, .Z(n_2147));
	notech_ao4 i_38934541(.A(n_59890), .B(n_17390), .C(n_59877), .D(n_17427)
		, .Z(n_2146));
	notech_and3 i_39234538(.A(n_2143), .B(n_2142), .C(n_1334), .Z(n_2145));
	notech_ao4 i_38634544(.A(n_59812), .B(n_17374), .C(n_59799), .D(n_17358)
		, .Z(n_2143));
	notech_ao4 i_38534545(.A(n_59786), .B(n_17350), .C(n_59773), .D(n_17366)
		, .Z(n_2142));
	notech_and4 i_39434536(.A(n_2136), .B(n_2138), .C(n_2140), .D(n_1320), .Z
		(n_2141));
	notech_ao4 i_39134539(.A(n_59838), .B(n_17382), .C(n_59825), .D(n_17414)
		, .Z(n_2140));
	notech_ao4 i_38434546(.A(n_59864), .B(n_17334), .C(n_59851), .D(n_17342)
		, .Z(n_2138));
	notech_ao4 i_38234548(.A(n_59976), .B(n_17318), .C(n_59957), .D(n_17326)
		, .Z(n_2136));
	notech_ao4 i_35934571(.A(n_59916), .B(n_17405), .C(n_59903), .D(n_17397)
		, .Z(n_2133));
	notech_ao4 i_35834572(.A(n_59890), .B(n_17389), .C(n_59877), .D(n_17425)
		, .Z(n_2132));
	notech_and3 i_36134569(.A(n_2129), .B(n_2128), .C(n_1316), .Z(n_2131));
	notech_ao4 i_35534575(.A(n_59812), .B(n_17373), .C(n_59799), .D(n_17357)
		, .Z(n_2129));
	notech_ao4 i_35434576(.A(n_59786), .B(n_17349), .C(n_59773), .D(n_17365)
		, .Z(n_2128));
	notech_and4 i_36334567(.A(n_2122), .B(n_2124), .C(n_2126), .D(n_1293), .Z
		(n_2127));
	notech_ao4 i_36034570(.A(n_59838), .B(n_17381), .C(n_59825), .D(n_17413)
		, .Z(n_2126));
	notech_ao4 i_35334577(.A(n_59864), .B(n_17333), .C(n_59851), .D(n_17341)
		, .Z(n_2124));
	notech_ao4 i_35134579(.A(n_59976), .B(n_17317), .C(n_59957), .D(n_17325)
		, .Z(n_2122));
	notech_ao4 i_32834602(.A(n_59916), .B(n_17404), .C(n_59903), .D(n_17396)
		, .Z(n_2119));
	notech_ao4 i_32734603(.A(n_59890), .B(n_17388), .C(n_59877), .D(n_17423)
		, .Z(n_2118));
	notech_and3 i_33034600(.A(n_2115), .B(n_2114), .C(n_1287), .Z(n_2117));
	notech_ao4 i_32434606(.A(n_59812), .B(n_17372), .C(n_59799), .D(n_17356)
		, .Z(n_2115));
	notech_ao4 i_32334607(.A(n_59786), .B(n_17348), .C(n_59773), .D(n_17364)
		, .Z(n_2114));
	notech_and4 i_33234598(.A(n_2108), .B(n_2110), .C(n_2112), .D(n_1273), .Z
		(n_2113));
	notech_ao4 i_32934601(.A(n_59838), .B(n_17380), .C(n_59825), .D(n_17412)
		, .Z(n_2112));
	notech_ao4 i_32234608(.A(n_59864), .B(n_17332), .C(n_59851), .D(n_17340)
		, .Z(n_2110));
	notech_ao4 i_32034610(.A(n_59976), .B(n_17316), .C(n_59952), .D(n_17324)
		, .Z(n_2108));
	notech_ao4 i_29734633(.A(n_59916), .B(n_17403), .C(n_59903), .D(n_17395)
		, .Z(n_2105));
	notech_ao4 i_29634634(.A(n_59890), .B(n_17387), .C(n_59877), .D(n_17421)
		, .Z(n_2104));
	notech_and3 i_29934631(.A(n_2101), .B(n_2100), .C(n_1270), .Z(n_2103));
	notech_ao4 i_29334637(.A(n_59812), .B(n_17371), .C(n_59799), .D(n_17355)
		, .Z(n_2101));
	notech_ao4 i_29234638(.A(n_59786), .B(n_17347), .C(n_59773), .D(n_17363)
		, .Z(n_2100));
	notech_and4 i_30134629(.A(n_2094), .B(n_2096), .C(n_2098), .D(n_1257), .Z
		(n_2099));
	notech_ao4 i_29834632(.A(n_59838), .B(n_17379), .C(n_59825), .D(n_17411)
		, .Z(n_2098));
	notech_ao4 i_29134639(.A(n_59864), .B(n_17331), .C(n_59851), .D(n_17339)
		, .Z(n_2096));
	notech_ao4 i_28934641(.A(n_59996), .B(n_17307), .C(n_59971), .D(n_17315)
		, .Z(n_2094));
	notech_ao4 i_26634664(.A(n_59916), .B(n_17401), .C(n_59903), .D(n_17393)
		, .Z(n_2091));
	notech_ao4 i_26534665(.A(n_59890), .B(n_17385), .C(n_59877), .D(n_17417)
		, .Z(n_2090));
	notech_and3 i_26834662(.A(n_2087), .B(n_2086), .C(n_1254), .Z(n_2089));
	notech_ao4 i_26234668(.A(n_59812), .B(n_17369), .C(n_59799), .D(n_17353)
		, .Z(n_2087));
	notech_ao4 i_26134669(.A(n_59786), .B(n_17345), .C(n_59773), .D(n_17361)
		, .Z(n_2086));
	notech_and4 i_27034660(.A(n_2080), .B(n_2082), .C(n_2084), .D(n_1241), .Z
		(n_2085));
	notech_ao4 i_26734663(.A(n_59838), .B(n_17377), .C(n_59825), .D(n_17409)
		, .Z(n_2084));
	notech_ao4 i_26034670(.A(n_59864), .B(n_17329), .C(n_59851), .D(n_17337)
		, .Z(n_2082));
	notech_ao4 i_25834672(.A(n_59964), .B(n_17313), .C(n_59945), .D(n_17321)
		, .Z(n_2080));
	notech_ao4 i_23534695(.A(n_59916), .B(n_17400), .C(n_59903), .D(n_17392)
		, .Z(n_2077));
	notech_ao4 i_23434696(.A(n_59890), .B(n_17384), .C(n_59877), .D(n_17416)
		, .Z(n_2076));
	notech_and3 i_23734693(.A(n_2073), .B(n_2072), .C(n_1238), .Z(n_2075));
	notech_ao4 i_23134699(.A(n_59812), .B(n_17368), .C(n_59799), .D(n_17352)
		, .Z(n_2073));
	notech_ao4 i_23034700(.A(n_59786), .B(n_17344), .C(n_59773), .D(n_17360)
		, .Z(n_2072));
	notech_and4 i_23934691(.A(n_2066), .B(n_2068), .C(n_2070), .D(n_122560143
		), .Z(n_2071));
	notech_ao4 i_23634694(.A(n_59838), .B(n_17376), .C(n_59825), .D(n_17408)
		, .Z(n_2070));
	notech_ao4 i_22934701(.A(n_59864), .B(n_17328), .C(n_59851), .D(n_17336)
		, .Z(n_2068));
	notech_ao4 i_22734703(.A(n_59964), .B(n_17312), .C(n_59945), .D(n_17320)
		, .Z(n_2066));
	notech_ao4 i_20434726(.A(n_59912), .B(n_17399), .C(n_59899), .D(n_17391)
		, .Z(n_2063));
	notech_ao4 i_20334727(.A(n_59886), .B(n_17383), .C(n_59873), .D(n_17415)
		, .Z(n_2062));
	notech_and3 i_20634724(.A(n_2059), .B(n_2058), .C(n_122260146), .Z(n_2061
		));
	notech_ao4 i_20034730(.A(n_59808), .B(n_17367), .C(n_59795), .D(n_17351)
		, .Z(n_2059));
	notech_ao4 i_19934731(.A(n_59782), .B(n_17343), .C(n_59769), .D(n_17359)
		, .Z(n_2058));
	notech_and4 i_20834722(.A(n_2052), .B(n_2054), .C(n_2056), .D(n_120960159
		), .Z(n_2057));
	notech_ao4 i_20534725(.A(n_59834), .B(n_17375), .C(n_59821), .D(n_17407)
		, .Z(n_2056));
	notech_ao4 i_19834732(.A(n_59860), .B(n_17327), .C(n_59847), .D(n_17335)
		, .Z(n_2054));
	notech_ao4 i_19634734(.A(n_59964), .B(n_17311), .C(n_59945), .D(n_17319)
		, .Z(n_2052));
	notech_ao4 i_17334757(.A(n_59912), .B(n_17398), .C(n_59899), .D(n_17390)
		, .Z(n_2049));
	notech_ao4 i_17234758(.A(n_59886), .B(n_17382), .C(n_59873), .D(n_17414)
		, .Z(n_2048));
	notech_and3 i_17534755(.A(n_2045), .B(n_2044), .C(n_120660162), .Z(n_2047
		));
	notech_ao4 i_16934761(.A(n_59808), .B(n_17366), .C(n_59795), .D(n_17350)
		, .Z(n_2045));
	notech_ao4 i_16834762(.A(n_59782), .B(n_17342), .C(n_59769), .D(n_17358)
		, .Z(n_2044));
	notech_and4 i_17734753(.A(n_2038), .B(n_2040), .C(n_2042), .D(n_119360175
		), .Z(n_2043));
	notech_ao4 i_17434756(.A(n_59834), .B(n_17374), .C(n_59821), .D(n_17406)
		, .Z(n_2042));
	notech_ao4 i_16734763(.A(n_59860), .B(n_17326), .C(n_59847), .D(n_17334)
		, .Z(n_2040));
	notech_ao4 i_16534765(.A(n_59964), .B(n_17310), .C(n_59945), .D(n_17318)
		, .Z(n_2038));
	notech_ao4 i_14234788(.A(n_59916), .B(n_17397), .C(n_59903), .D(n_17389)
		, .Z(n_2035));
	notech_ao4 i_14134789(.A(n_59890), .B(n_17381), .C(n_59877), .D(n_17413)
		, .Z(n_2034));
	notech_and3 i_14434786(.A(n_2031), .B(n_2030), .C(n_119060178), .Z(n_2033
		));
	notech_ao4 i_13834792(.A(n_59812), .B(n_17365), .C(n_59799), .D(n_17349)
		, .Z(n_2031));
	notech_ao4 i_13734793(.A(n_59786), .B(n_17341), .C(n_59773), .D(n_17357)
		, .Z(n_2030));
	notech_and4 i_14634784(.A(n_2024), .B(n_2026), .C(n_2028), .D(n_1177), .Z
		(n_2029));
	notech_ao4 i_14334787(.A(n_59838), .B(n_17373), .C(n_59825), .D(n_17405)
		, .Z(n_2028));
	notech_ao4 i_13634794(.A(n_59864), .B(n_17325), .C(n_59851), .D(n_17333)
		, .Z(n_2026));
	notech_ao4 i_13434796(.A(n_59964), .B(n_17309), .C(n_59945), .D(n_17317)
		, .Z(n_2024));
	notech_ao4 i_11134819(.A(n_59916), .B(n_17396), .C(n_59903), .D(n_17388)
		, .Z(n_2021));
	notech_ao4 i_11034820(.A(n_59890), .B(n_17380), .C(n_59877), .D(n_17412)
		, .Z(n_2020));
	notech_and3 i_11334817(.A(n_2017), .B(n_2016), .C(n_1174), .Z(n_2019));
	notech_ao4 i_10734823(.A(n_59812), .B(n_17364), .C(n_59799), .D(n_17348)
		, .Z(n_2017));
	notech_ao4 i_10634824(.A(n_59786), .B(n_17340), .C(n_59773), .D(n_17356)
		, .Z(n_2016));
	notech_and4 i_11534815(.A(n_2010), .B(n_2012), .C(n_2014), .D(n_1161), .Z
		(n_2015));
	notech_ao4 i_11234818(.A(n_59838), .B(n_17372), .C(n_59825), .D(n_17404)
		, .Z(n_2014));
	notech_ao4 i_10534825(.A(n_59864), .B(n_17324), .C(n_59851), .D(n_17332)
		, .Z(n_2012));
	notech_ao4 i_10334827(.A(n_59964), .B(n_17308), .C(n_59945), .D(n_17316)
		, .Z(n_2010));
	notech_ao4 i_7934850(.A(n_59916), .B(n_17395), .C(n_59903), .D(n_17387),
		 .Z(n_2007));
	notech_nand3 i_1034912(.A(n_59933), .B(n_3078), .C(n_3072), .Z(n_2006)
		);
	notech_nand3 i_934913(.A(n_3078), .B(n_3074), .C(n_59933), .Z(n_2005));
	notech_ao4 i_7834851(.A(n_59890), .B(n_17379), .C(n_59877), .D(n_17411),
		 .Z(n_2004));
	notech_nand3 i_834914(.A(n_3072), .B(n_3069), .C(n_59933), .Z(n_2003));
	notech_nand3 i_434918(.A(n_3076), .B(n_3072), .C(n_59937), .Z(n_2002));
	notech_and3 i_8234848(.A(n_1999), .B(n_1996), .C(n_1158), .Z(n_2001));
	notech_ao4 i_7534854(.A(n_59812), .B(n_17363), .C(n_59799), .D(n_17347),
		 .Z(n_1999));
	notech_nand3 i_734915(.A(n_3086), .B(n_3072), .C(n_3091), .Z(n_1998));
	notech_nand3 i_634916(.A(n_3082), .B(n_3076), .C(n_3091), .Z(n_1997));
	notech_ao4 i_7434855(.A(n_59786), .B(n_17339), .C(n_59773), .D(n_17355),
		 .Z(n_1996));
	notech_nao3 i_534917(.A(n_3076), .B(n_3091), .C(n_3084), .Z(n_1995));
	notech_nand3 i_334919(.A(n_3086), .B(n_3074), .C(n_3091), .Z(n_1994));
	notech_and4 i_8434846(.A(n_1983), .B(n_1987), .C(n_1992), .D(n_1145), .Z
		(n_1993));
	notech_ao4 i_8134849(.A(n_59838), .B(n_17371), .C(n_59825), .D(n_17403),
		 .Z(n_1992));
	notech_nand3 i_1234910(.A(n_3074), .B(n_59933), .C(n_3069), .Z(n_1991)
		);
	notech_nand3 i_1134911(.A(n_59937), .B(n_3076), .C(n_3074), .Z(n_1990)
		);
	notech_and4 i_1834904(.A(n_60093), .B(n_60077), .C(n_3088), .D(n_3091), 
		.Z(n_1989));
	notech_ao4 i_7334856(.A(n_59864), .B(n_17323), .C(n_59851), .D(n_17331),
		 .Z(n_1987));
	notech_nao3 i_134920(.A(n_3078), .B(n_3091), .C(n_3084), .Z(n_1986));
	notech_nand3 i_034921(.A(n_60101), .B(n_3078), .C(n_3091), .Z(n_1985));
	notech_ao4 i_7034858(.A(n_59964), .B(n_17307), .C(n_59945), .D(n_17315),
		 .Z(n_1983));
	notech_nand2 i_428391(.A(n_2713), .B(n_1981), .Z(n_35399));
	notech_or4 i_225432682(.A(n_62854), .B(n_61430), .C(n_61398), .D(n_17871
		), .Z(n_1981));
	notech_nand2 i_1228399(.A(n_2712), .B(n_1979), .Z(n_35447));
	notech_or4 i_222232714(.A(n_62854), .B(n_61430), .C(n_61398), .D(n_17870
		), .Z(n_1979));
	notech_nand2 i_2028407(.A(n_2711), .B(n_1977), .Z(n_35495));
	notech_or4 i_219032746(.A(n_62854), .B(n_61430), .C(n_61398), .D(n_17869
		), .Z(n_1977));
	notech_nand2 i_2828415(.A(n_2710), .B(n_1975), .Z(n_35543));
	notech_or4 i_215832778(.A(n_62854), .B(n_61430), .C(n_61398), .D(n_17868
		), .Z(n_1975));
	notech_and4 i_6625032(.A(n_2707), .B(n_2706), .C(n_2701), .D(n_2705), .Z
		(squeue_65101035));
	notech_nand3 i_162133309(.A(n_59662), .B(n_59937), .C(queue[65]), .Z(n_1974
		));
	notech_nand3 i_160833322(.A(n_3086), .B(n_60101), .C(queue[73]), .Z(n_1961
		));
	notech_and4 i_5425020(.A(n_2693), .B(n_2692), .C(n_2687), .D(n_2691), .Z
		(squeue_53101036));
	notech_nand3 i_159033340(.A(n_59662), .B(n_59933), .C(queue[53]), .Z(n_1958
		));
	notech_nand3 i_157733353(.A(n_61409), .B(n_60101), .C(queue[61]), .Z(n_1945
		));
	notech_and4 i_5325019(.A(n_2679), .B(n_2678), .C(n_2673), .D(n_2677), .Z
		(squeue_52101037));
	notech_nand3 i_155933371(.A(n_59662), .B(n_59933), .C(queue[52]), .Z(n_1942
		));
	notech_nand3 i_154633384(.A(n_61409), .B(n_60101), .C(queue[60]), .Z(n_1929
		));
	notech_and4 i_5225018(.A(n_2665), .B(n_2664), .C(n_2659), .D(n_2663), .Z
		(squeue_51101038));
	notech_nand3 i_152833402(.A(n_59662), .B(n_59933), .C(queue[51]), .Z(n_1926
		));
	notech_nand3 i_151533415(.A(n_61409), .B(n_60101), .C(queue[59]), .Z(n_1913
		));
	notech_and4 i_5125017(.A(n_2651), .B(n_2650), .C(n_2645), .D(n_2649), .Z
		(squeue_50101039));
	notech_nand3 i_149733433(.A(n_59662), .B(n_59933), .C(queue[50]), .Z(n_1910
		));
	notech_nand3 i_148433446(.A(n_61409), .B(n_60101), .C(queue[58]), .Z(n_1897
		));
	notech_and4 i_5025016(.A(n_2637), .B(n_2636), .C(n_2631), .D(n_2635), .Z
		(squeue_49101040));
	notech_nand3 i_146633464(.A(n_59662), .B(n_59938), .C(queue[49]), .Z(n_1894
		));
	notech_nand3 i_145333477(.A(n_61409), .B(n_3082), .C(queue[57]), .Z(n_1881
		));
	notech_and4 i_4925015(.A(n_2623), .B(n_2622), .C(n_2617), .D(n_2621), .Z
		(squeue_48101041));
	notech_nand3 i_143533495(.A(n_59662), .B(n_59940), .C(queue[48]), .Z(n_1878
		));
	notech_or2 i_142233508(.A(n_59964), .B(n_17355), .Z(n_1865));
	notech_and4 i_4825014(.A(n_2609), .B(n_2608), .C(n_2603), .D(n_2607), .Z
		(squeue_47101042));
	notech_nand3 i_140433526(.A(n_59662), .B(n_59940), .C(queue[47]), .Z(n_1862
		));
	notech_or2 i_139133539(.A(n_59996), .B(n_17346), .Z(n_1849));
	notech_and4 i_4725013(.A(n_2595), .B(n_2594), .C(n_2589), .D(n_2593), .Z
		(squeue_46101043));
	notech_nand3 i_137333557(.A(n_59662), .B(n_59940), .C(queue[46]), .Z(n_1846
		));
	notech_or2 i_136033570(.A(n_59996), .B(n_17345), .Z(n_1833));
	notech_and4 i_4625012(.A(n_2581), .B(n_2580), .C(n_2575), .D(n_2579), .Z
		(squeue_45101044));
	notech_nand3 i_134233588(.A(n_59662), .B(n_59940), .C(queue[45]), .Z(n_1830
		));
	notech_nand3 i_132933601(.A(n_61409), .B(n_3082), .C(queue[53]), .Z(n_1817
		));
	notech_and4 i_4525011(.A(n_2567), .B(n_2566), .C(n_2561), .D(n_2565), .Z
		(squeue_44101045));
	notech_nand3 i_131133619(.A(n_59669), .B(n_59940), .C(queue[44]), .Z(n_1814
		));
	notech_nand3 i_129833632(.A(n_3086), .B(n_3082), .C(queue[52]), .Z(n_1801
		));
	notech_and4 i_4425010(.A(n_2553), .B(n_2552), .C(n_2547), .D(n_2551), .Z
		(squeue_43101046));
	notech_nand3 i_128033650(.A(n_59669), .B(n_59940), .C(queue[43]), .Z(n_1798
		));
	notech_nand3 i_126733663(.A(n_3086), .B(n_3082), .C(queue[51]), .Z(n_1785
		));
	notech_and4 i_4325009(.A(n_2539), .B(n_2538), .C(n_2533), .D(n_2537), .Z
		(squeue_42101047));
	notech_nand3 i_124933681(.A(n_59669), .B(n_59940), .C(queue[42]), .Z(n_1782
		));
	notech_nand3 i_123633694(.A(n_3086), .B(n_3082), .C(queue[50]), .Z(n_1769
		));
	notech_and4 i_4225008(.A(n_2525), .B(n_2524), .C(n_2519), .D(n_2523), .Z
		(squeue_41101048));
	notech_nand3 i_121833712(.A(n_59669), .B(n_59940), .C(queue[41]), .Z(n_1766
		));
	notech_nand3 i_120533725(.A(n_3086), .B(n_3082), .C(queue[49]), .Z(n_1753
		));
	notech_and4 i_4125007(.A(n_2511), .B(n_2510), .C(n_2505), .D(n_2509), .Z
		(squeue_40101049));
	notech_nand3 i_118733743(.A(n_59669), .B(n_59940), .C(queue[40]), .Z(n_1750
		));
	notech_or2 i_117433756(.A(n_59945), .B(n_17355), .Z(n_1737));
	notech_and4 i_4025006(.A(n_2497), .B(n_2496), .C(n_2491), .D(n_2495), .Z
		(squeue_39101050));
	notech_nand3 i_115633774(.A(n_59669), .B(n_59940), .C(queue[39]), .Z(n_1734
		));
	notech_or2 i_114333787(.A(n_59996), .B(n_17338), .Z(n_1721));
	notech_and4 i_3925005(.A(n_2483), .B(n_2482), .C(n_2477), .D(n_2481), .Z
		(squeue_38101051));
	notech_nand3 i_112533805(.A(n_59669), .B(n_59940), .C(queue[38]), .Z(n_1718
		));
	notech_or2 i_111233818(.A(n_59996), .B(n_17337), .Z(n_1705));
	notech_and4 i_3725003(.A(n_2469), .B(n_2468), .C(n_2463), .D(n_2467), .Z
		(squeue_36101052));
	notech_nand3 i_109433836(.A(n_59669), .B(n_59940), .C(queue[36]), .Z(n_1702
		));
	notech_nand3 i_108133849(.A(n_3086), .B(n_3082), .C(queue[44]), .Z(n_1689
		));
	notech_and4 i_3625002(.A(n_2455), .B(n_2454), .C(n_2449), .D(n_2453), .Z
		(squeue_35101053));
	notech_nand3 i_106333867(.A(n_59669), .B(n_59940), .C(queue[35]), .Z(n_1686
		));
	notech_nand3 i_105033880(.A(n_3086), .B(n_3082), .C(queue[43]), .Z(n_1673
		));
	notech_and4 i_3525001(.A(n_2441), .B(n_2440), .C(n_2435), .D(n_2439), .Z
		(squeue_34101054));
	notech_nand3 i_103233898(.A(n_59669), .B(n_59940), .C(queue[34]), .Z(n_1670
		));
	notech_nand3 i_101933911(.A(n_3086), .B(n_3082), .C(queue[42]), .Z(n_1657
		));
	notech_and4 i_3425000(.A(n_2427), .B(n_2426), .C(n_2421), .D(n_2425), .Z
		(squeue_33101055));
	notech_nand3 i_100133929(.A(n_59669), .B(n_59940), .C(queue[33]), .Z(n_1654
		));
	notech_nand3 i_98833942(.A(n_3086), .B(n_3082), .C(queue[41]), .Z(n_1641
		));
	notech_and4 i_3324999(.A(n_2413), .B(n_2412), .C(n_2407), .D(n_2411), .Z
		(squeue_32101056));
	notech_nand3 i_97033960(.A(n_59669), .B(n_59940), .C(queue[32]), .Z(n_1638
		));
	notech_nand3 i_95733973(.A(n_3086), .B(n_3082), .C(queue[40]), .Z(n_1625
		));
	notech_and4 i_3224998(.A(n_2399), .B(n_2398), .C(n_2393), .D(n_2397), .Z
		(squeue_31101057));
	notech_xor2 i_4535424(.A(fault_wptr[0]), .B(fault_wptr[1]), .Z(n_99957531
		));
	notech_and2 i_3635432(.A(n_17301), .B(n_17300), .Z(n_100257534));
	notech_or2 i_28435189(.A(n_100457536), .B(n_309459575), .Z(n_100357535)
		);
	notech_ao4 i_3435434(.A(n_61359), .B(n_312559606), .C(n_101057542), .D(n_101157543
		), .Z(n_100457536));
	notech_or4 i_28135192(.A(n_61153), .B(n_309459575), .C(n_17294), .D(n_100257534
		), .Z(n_100657538));
	notech_nao3 i_28235191(.A(n_14128702), .B(pg_fault), .C(n_309459575), .Z
		(n_100757539));
	notech_nao3 i_46535008(.A(n_8288), .B(n_14128702), .C(pg_fault), .Z(n_101057542
		));
	notech_nand2 i_46335010(.A(n_34592), .B(n_17872), .Z(n_101157543));
	notech_nao3 i_7271(.A(n_63814), .B(n_130357803), .C(tagV[1]), .Z(n_8288)
		);
	notech_nand2 i_1434908(.A(n_34592), .B(n_17292), .Z(n_8291));
	notech_ao4 i_4634880(.A(n_130657804), .B(n_8291), .C(n_312559606), .D(n_61359
		), .Z(n_101657548));
	notech_nand3 i_6634960(.A(n_61567), .B(n_8293), .C(n_309659577), .Z(n_7794
		));
	notech_ao3 i_4934877(.A(n_17294), .B(n_61398), .C(n_309459575), .Z(n_101957551
		));
	notech_nao3 i_65526(.A(n_7794), .B(n_309559576), .C(n_101957551), .Z(\nbus_12122[0] 
		));
	notech_ao4 i_21628603(.A(n_61359), .B(n_17820), .C(n_56561), .D(n_17873)
		, .Z(n_36671));
	notech_or4 i_174033190(.A(n_62854), .B(n_61430), .C(n_61398), .D(n_17874
		), .Z(n_102257554));
	notech_nand2 i_12828515(.A(n_130957807), .B(n_102257554), .Z(n_36143));
	notech_or4 i_174433186(.A(n_62854), .B(n_61430), .C(n_61398), .D(n_17875
		), .Z(n_102457556));
	notech_nand2 i_12728514(.A(n_131257808), .B(n_102457556), .Z(n_36137));
	notech_or4 i_174833182(.A(n_62854), .B(n_61430), .C(n_61398), .D(n_17876
		), .Z(n_102657558));
	notech_nand2 i_12628513(.A(n_131357809), .B(n_102657558), .Z(n_36131));
	notech_or4 i_175233178(.A(n_62854), .B(n_61430), .C(n_61398), .D(n_17877
		), .Z(n_102957560));
	notech_nand2 i_12528512(.A(n_131657810), .B(n_102957560), .Z(n_36125));
	notech_or4 i_175633174(.A(n_62854), .B(n_61431), .C(n_61398), .D(n_17878
		), .Z(n_103357562));
	notech_nand2 i_12428511(.A(n_131757811), .B(n_103357562), .Z(n_36119));
	notech_or4 i_176033170(.A(n_62858), .B(n_61431), .C(n_61399), .D(n_17879
		), .Z(n_103957564));
	notech_nand2 i_12328510(.A(n_131957812), .B(n_103957564), .Z(n_36113));
	notech_or4 i_176433166(.A(n_62858), .B(n_61430), .C(n_61399), .D(n_17880
		), .Z(n_104157566));
	notech_nand2 i_12228509(.A(n_132057813), .B(n_104157566), .Z(n_36107));
	notech_or4 i_176833162(.A(n_62858), .B(n_61430), .C(n_61398), .D(n_17881
		), .Z(n_104357568));
	notech_nand2 i_12128508(.A(n_132257814), .B(n_104357568), .Z(n_36101));
	notech_or4 i_177233158(.A(n_62858), .B(n_61430), .C(n_61398), .D(n_17882
		), .Z(n_104657570));
	notech_nand2 i_12028507(.A(n_132357815), .B(n_104657570), .Z(n_36095));
	notech_or4 i_177633154(.A(n_62858), .B(n_61430), .C(n_61398), .D(n_17883
		), .Z(n_104857572));
	notech_nand2 i_11928506(.A(n_132457816), .B(n_104857572), .Z(n_36089));
	notech_or4 i_178033150(.A(n_62858), .B(n_61430), .C(n_61398), .D(n_17884
		), .Z(n_105357574));
	notech_nand2 i_11828505(.A(n_132557817), .B(n_105357574), .Z(n_36083));
	notech_or4 i_178433146(.A(n_62858), .B(n_61426), .C(n_61398), .D(n_17885
		), .Z(n_105557576));
	notech_nand2 i_11728504(.A(n_132657818), .B(n_105557576), .Z(n_36077));
	notech_or4 i_179233138(.A(n_62858), .B(n_61426), .C(n_61394), .D(n_17886
		), .Z(n_105757578));
	notech_nand2 i_11528502(.A(n_132757819), .B(n_105757578), .Z(n_36065));
	notech_or4 i_179633134(.A(n_62852), .B(n_61426), .C(n_61394), .D(n_17887
		), .Z(n_105957580));
	notech_nand2 i_11428501(.A(n_132857820), .B(n_105957580), .Z(n_36059));
	notech_or4 i_180033130(.A(n_62852), .B(n_61426), .C(n_61394), .D(n_17888
		), .Z(n_106157582));
	notech_nand2 i_11328500(.A(n_132957821), .B(n_106157582), .Z(n_36053));
	notech_or4 i_180433126(.A(n_62852), .B(n_61426), .C(n_61394), .D(n_17889
		), .Z(n_106357584));
	notech_nand2 i_11228499(.A(n_133057822), .B(n_106357584), .Z(n_36047));
	notech_or4 i_180833122(.A(n_62852), .B(n_61426), .C(n_61394), .D(n_17890
		), .Z(n_106557586));
	notech_nand2 i_11128498(.A(n_133157823), .B(n_106557586), .Z(n_36041));
	notech_or4 i_181233118(.A(n_62852), .B(n_61426), .C(n_61394), .D(n_17891
		), .Z(n_106757588));
	notech_nand2 i_11028497(.A(n_133257824), .B(n_106757588), .Z(n_36035));
	notech_or4 i_181633114(.A(n_62852), .B(n_61426), .C(n_61394), .D(n_17892
		), .Z(n_106957590));
	notech_nand2 i_10928496(.A(n_133357825), .B(n_106957590), .Z(n_36029));
	notech_or4 i_182033110(.A(n_62852), .B(n_61430), .C(n_61394), .D(n_17893
		), .Z(n_107157592));
	notech_nand2 i_10828495(.A(n_133457826), .B(n_107157592), .Z(n_36023));
	notech_or4 i_182433106(.A(n_62852), .B(n_61426), .C(n_61398), .D(n_17894
		), .Z(n_107357594));
	notech_nand2 i_10728494(.A(n_133557827), .B(n_107357594), .Z(n_36017));
	notech_or4 i_182833102(.A(n_62852), .B(n_61430), .C(n_61394), .D(n_17895
		), .Z(n_107557596));
	notech_nand2 i_10628493(.A(n_133657828), .B(n_107557596), .Z(n_36011));
	notech_or4 i_183233098(.A(n_62854), .B(n_61430), .C(n_61398), .D(n_17896
		), .Z(n_107757598));
	notech_nand2 i_10528492(.A(n_133757829), .B(n_107757598), .Z(n_36005));
	notech_or4 i_183633094(.A(n_62854), .B(n_61426), .C(n_61398), .D(n_17897
		), .Z(n_107957600));
	notech_nand2 i_10428491(.A(n_133857830), .B(n_107957600), .Z(n_35999));
	notech_or4 i_184033090(.A(n_62854), .B(n_61426), .C(n_61394), .D(n_17898
		), .Z(n_108157602));
	notech_nand2 i_10328490(.A(n_133957831), .B(n_108157602), .Z(n_35993));
	notech_or4 i_184433086(.A(n_62854), .B(n_61426), .C(n_61394), .D(n_17899
		), .Z(n_108357604));
	notech_nand2 i_10228489(.A(n_134057832), .B(n_108357604), .Z(n_35987));
	notech_or4 i_184933081(.A(n_62852), .B(n_61426), .C(n_61394), .D(n_17900
		), .Z(n_108657607));
	notech_nand2 i_10128488(.A(n_134157833), .B(n_108657607), .Z(n_35981));
	notech_or4 i_185333077(.A(n_62852), .B(n_61431), .C(n_61394), .D(n_17901
		), .Z(n_108857609));
	notech_nand2 i_10028487(.A(n_134257834), .B(n_108857609), .Z(n_35975));
	notech_or4 i_185833072(.A(n_62854), .B(n_61433), .C(n_61399), .D(n_17902
		), .Z(n_109157612));
	notech_nand2 i_9928486(.A(n_134357835), .B(n_109157612), .Z(n_35969));
	notech_or4 i_186233068(.A(n_62852), .B(n_61433), .C(n_61401), .D(n_17903
		), .Z(n_109357614));
	notech_nand2 i_9828485(.A(n_134457836), .B(n_109357614), .Z(n_35963));
	notech_or4 i_186733063(.A(n_62861), .B(n_61433), .C(n_61401), .D(n_17904
		), .Z(n_109657617));
	notech_nand2 i_9728484(.A(n_134557837), .B(n_109657617), .Z(n_35957));
	notech_or4 i_187133059(.A(n_62861), .B(n_61433), .C(n_61401), .D(n_17905
		), .Z(n_109857619));
	notech_nand2 i_9628483(.A(n_134657838), .B(n_109857619), .Z(n_35951));
	notech_or4 i_187633054(.A(n_62861), .B(n_61433), .C(n_61401), .D(n_17906
		), .Z(n_110157622));
	notech_nand2 i_9528482(.A(n_134757839), .B(n_110157622), .Z(n_35945));
	notech_or4 i_188133049(.A(n_62861), .B(n_61433), .C(n_61401), .D(n_17907
		), .Z(n_110457625));
	notech_nand2 i_9428481(.A(n_134857840), .B(n_110457625), .Z(n_35939));
	notech_or4 i_188533045(.A(n_62859), .B(n_61433), .C(n_61401), .D(n_17908
		), .Z(n_110657627));
	notech_nand2 i_9328480(.A(n_134957841), .B(n_110657627), .Z(n_35933));
	notech_or4 i_189033040(.A(n_62859), .B(n_61433), .C(n_61401), .D(n_17909
		), .Z(n_110957630));
	notech_nand2 i_9228479(.A(n_135057842), .B(n_110957630), .Z(n_35927));
	notech_or4 i_190033030(.A(n_62861), .B(n_61433), .C(n_61401), .D(n_17910
		), .Z(n_111257633));
	notech_nand2 i_9028477(.A(n_135157843), .B(n_111257633), .Z(n_35915));
	notech_or4 i_190533025(.A(n_62859), .B(n_61433), .C(n_61401), .D(n_17911
		), .Z(n_111557636));
	notech_nand2 i_8928476(.A(n_135257844), .B(n_111557636), .Z(n_35909));
	notech_or4 i_191033020(.A(n_62861), .B(n_61433), .C(n_61401), .D(n_17873
		), .Z(n_112257639));
	notech_nand2 i_8828475(.A(n_135357845), .B(n_112257639), .Z(n_35903));
	notech_or4 i_191533015(.A(n_62861), .B(n_61433), .C(n_61401), .D(n_17912
		), .Z(n_112457641));
	notech_nand2 i_8728474(.A(n_135457846), .B(n_112457641), .Z(n_35897));
	notech_or4 i_192033010(.A(n_62861), .B(n_61433), .C(n_61401), .D(n_17913
		), .Z(n_112757643));
	notech_nand2 i_8628473(.A(n_135557847), .B(n_112757643), .Z(n_35891));
	notech_or4 i_192433006(.A(n_62861), .B(n_61433), .C(n_61401), .D(n_17914
		), .Z(n_112957645));
	notech_nand2 i_8528472(.A(n_135657848), .B(n_112957645), .Z(n_35885));
	notech_or4 i_192833002(.A(n_62861), .B(n_61433), .C(n_61401), .D(n_17915
		), .Z(n_113157647));
	notech_nand2 i_8428471(.A(n_135757849), .B(n_113157647), .Z(n_35879));
	notech_or4 i_193232998(.A(n_62861), .B(n_61433), .C(n_61401), .D(n_17916
		), .Z(n_113357649));
	notech_nand2 i_8328470(.A(n_135857850), .B(n_113357649), .Z(n_35873));
	notech_or4 i_193632994(.A(n_62861), .B(n_61433), .C(n_61401), .D(n_17917
		), .Z(n_113657651));
	notech_nand2 i_8228469(.A(n_135957851), .B(n_113657651), .Z(n_35867));
	notech_or4 i_194032990(.A(n_62861), .B(n_61431), .C(n_61401), .D(n_17918
		), .Z(n_113857653));
	notech_nand2 i_8128468(.A(n_136057852), .B(n_113857653), .Z(n_35861));
	notech_or4 i_194432986(.A(n_62861), .B(n_61431), .C(n_61399), .D(n_17919
		), .Z(n_114357655));
	notech_nand2 i_8028467(.A(n_136157853), .B(n_114357655), .Z(n_35855));
	notech_or4 i_194832982(.A(n_62858), .B(n_61431), .C(n_61399), .D(n_17920
		), .Z(n_114557657));
	notech_nand2 i_7928466(.A(n_136257854), .B(n_114557657), .Z(n_35849));
	notech_or4 i_195232978(.A(n_62858), .B(n_61431), .C(n_61399), .D(n_17921
		), .Z(n_114757659));
	notech_nand2 i_7828465(.A(n_136357855), .B(n_114757659), .Z(n_35843));
	notech_or4 i_195632974(.A(n_62859), .B(n_61431), .C(n_61399), .D(n_17922
		), .Z(n_114957661));
	notech_nand2 i_7728464(.A(n_136457856), .B(n_114957661), .Z(n_35837));
	notech_or4 i_196032970(.A(n_62859), .B(n_61431), .C(n_61399), .D(n_17923
		), .Z(n_115157663));
	notech_nand2 i_7628463(.A(n_136557857), .B(n_115157663), .Z(n_35831));
	notech_or4 i_196432966(.A(n_62858), .B(n_61431), .C(n_61399), .D(n_17924
		), .Z(n_115357665));
	notech_nand2 i_7528462(.A(n_136657858), .B(n_115357665), .Z(n_35825));
	notech_or4 i_196832962(.A(n_62858), .B(n_61431), .C(n_61399), .D(n_17925
		), .Z(n_115557667));
	notech_nand2 i_7428461(.A(n_136757859), .B(n_115557667), .Z(n_35819));
	notech_or4 i_197232958(.A(n_62858), .B(n_61431), .C(n_61399), .D(n_17926
		), .Z(n_115757669));
	notech_nand2 i_7328460(.A(n_136857860), .B(n_115757669), .Z(n_35813));
	notech_or4 i_197632954(.A(n_62858), .B(n_61431), .C(n_61399), .D(n_17927
		), .Z(n_115957671));
	notech_nand2 i_7228459(.A(n_136957861), .B(n_115957671), .Z(n_35807));
	notech_or4 i_198032950(.A(n_62859), .B(n_61433), .C(n_61399), .D(n_17928
		), .Z(n_116157673));
	notech_nand2 i_7128458(.A(n_137057862), .B(n_116157673), .Z(n_35801));
	notech_or4 i_198432946(.A(n_62859), .B(n_61431), .C(n_61401), .D(n_17929
		), .Z(n_116357675));
	notech_nand2 i_7028457(.A(n_137157863), .B(n_116357675), .Z(n_35795));
	notech_or4 i_198832942(.A(n_62859), .B(n_61431), .C(n_61399), .D(n_17930
		), .Z(n_116557677));
	notech_nand2 i_6928456(.A(n_137257864), .B(n_116557677), .Z(n_35789));
	notech_or4 i_199232938(.A(n_62859), .B(n_61431), .C(n_61399), .D(n_17931
		), .Z(n_116757679));
	notech_nand2 i_6828455(.A(n_137357865), .B(n_116757679), .Z(n_35783));
	notech_or4 i_199632934(.A(n_62859), .B(n_61431), .C(n_61399), .D(n_17932
		), .Z(n_116957681));
	notech_nand2 i_6728454(.A(n_137457866), .B(n_116957681), .Z(n_35777));
	notech_or4 i_200032930(.A(n_62859), .B(n_61431), .C(n_61399), .D(n_17933
		), .Z(n_117157683));
	notech_nand2 i_6628453(.A(n_137557867), .B(n_117157683), .Z(n_35771));
	notech_or4 i_200432926(.A(n_62859), .B(n_61426), .C(n_61399), .D(n_17934
		), .Z(n_117357685));
	notech_nand2 i_6528452(.A(n_137657868), .B(n_117357685), .Z(n_35765));
	notech_or4 i_200832922(.A(n_62859), .B(n_61419), .C(n_61394), .D(n_17935
		), .Z(n_117557687));
	notech_nand2 i_6428451(.A(n_137757869), .B(n_117557687), .Z(n_35759));
	notech_or4 i_201232918(.A(n_62859), .B(n_61419), .C(n_61388), .D(n_17936
		), .Z(n_117757689));
	notech_nand2 i_6328450(.A(n_137857870), .B(n_117757689), .Z(n_35753));
	notech_or4 i_201632914(.A(code_req), .B(n_61419), .C(n_61388), .D(n_17937
		), .Z(n_117957691));
	notech_nand2 i_6228449(.A(n_137957871), .B(n_117957691), .Z(n_35747));
	notech_or4 i_202032910(.A(code_req), .B(n_61419), .C(n_61388), .D(n_17938
		), .Z(n_118157693));
	notech_nand2 i_6128448(.A(n_138057872), .B(n_118157693), .Z(n_35741));
	notech_or4 i_202432906(.A(n_62846), .B(n_61419), .C(n_61388), .D(n_17939
		), .Z(n_118357695));
	notech_nand2 i_6028447(.A(n_138157873), .B(n_118357695), .Z(n_35735));
	notech_or4 i_202832902(.A(n_62846), .B(n_61419), .C(n_61388), .D(n_17940
		), .Z(n_118557697));
	notech_nand2 i_5928446(.A(n_138257874), .B(n_118557697), .Z(n_35729));
	notech_or4 i_203232898(.A(code_req), .B(n_61419), .C(n_61386), .D(n_17941
		), .Z(n_118757699));
	notech_nand2 i_5828445(.A(n_138357875), .B(n_118757699), .Z(n_35723));
	notech_or4 i_203632894(.A(code_req), .B(n_61419), .C(n_61388), .D(n_17942
		), .Z(n_118957701));
	notech_nand2 i_5728444(.A(n_138457876), .B(n_118957701), .Z(n_35717));
	notech_or4 i_204032890(.A(code_req), .B(n_61421), .C(n_61388), .D(n_17943
		), .Z(n_119157703));
	notech_nand2 i_5628443(.A(n_138557877), .B(n_119157703), .Z(n_35711));
	notech_or4 i_204432886(.A(code_req), .B(n_61421), .C(n_61388), .D(n_17944
		), .Z(n_119357705));
	notech_nand2 i_5528442(.A(n_138657878), .B(n_119357705), .Z(n_35705));
	notech_or4 i_204832882(.A(n_62846), .B(n_61421), .C(n_61388), .D(n_17945
		), .Z(n_119557707));
	notech_nand2 i_5428441(.A(n_138757879), .B(n_119557707), .Z(n_35699));
	notech_or4 i_205232878(.A(n_62846), .B(n_61421), .C(n_61388), .D(n_17946
		), .Z(n_119757709));
	notech_nand2 i_5328440(.A(n_138857880), .B(n_119757709), .Z(n_35693));
	notech_or4 i_205632874(.A(n_62846), .B(n_61419), .C(n_61388), .D(n_17947
		), .Z(n_119957711));
	notech_nand2 i_5228439(.A(n_138957881), .B(n_119957711), .Z(n_35687));
	notech_or4 i_206032870(.A(n_62846), .B(n_61419), .C(n_61388), .D(n_17948
		), .Z(n_120157713));
	notech_nand2 i_5128438(.A(n_139057882), .B(n_120157713), .Z(n_35681));
	notech_or4 i_206432866(.A(n_62846), .B(n_61421), .C(n_61388), .D(n_17949
		), .Z(n_120357715));
	notech_nand2 i_5028437(.A(n_139157883), .B(n_120357715), .Z(n_35675));
	notech_or4 i_206832862(.A(n_62846), .B(n_61421), .C(n_61388), .D(n_17950
		), .Z(n_120557717));
	notech_nand2 i_4928436(.A(n_139257884), .B(n_120557717), .Z(n_35669));
	notech_or4 i_207232858(.A(n_62846), .B(n_61419), .C(n_61388), .D(n_17951
		), .Z(n_120757719));
	notech_nand2 i_4828435(.A(n_139357885), .B(n_120757719), .Z(n_35663));
	notech_or4 i_207632854(.A(n_62846), .B(n_61418), .C(n_61386), .D(n_17952
		), .Z(n_120957721));
	notech_nand2 i_4728434(.A(n_139457886), .B(n_120957721), .Z(n_35657));
	notech_or4 i_208032850(.A(code_req), .B(n_61418), .C(n_61386), .D(n_17953
		), .Z(n_121157723));
	notech_nand2 i_4628433(.A(n_139557887), .B(n_121157723), .Z(n_35651));
	notech_or4 i_208432846(.A(n_62841), .B(n_61418), .C(n_61386), .D(n_17954
		), .Z(n_121357725));
	notech_nand2 i_4528432(.A(n_139657888), .B(n_121357725), .Z(n_35645));
	notech_or4 i_208832842(.A(n_62841), .B(n_61418), .C(n_61386), .D(n_17955
		), .Z(n_121557727));
	notech_nand2 i_4428431(.A(n_139757889), .B(n_121557727), .Z(n_35639));
	notech_or4 i_209232838(.A(n_62841), .B(n_61418), .C(n_61386), .D(n_17956
		), .Z(n_121757729));
	notech_nand2 i_4328430(.A(n_139857890), .B(n_121757729), .Z(n_35633));
	notech_or4 i_209632834(.A(n_62841), .B(n_61418), .C(n_61386), .D(n_17957
		), .Z(n_121957731));
	notech_nand2 i_4228429(.A(n_139957891), .B(n_121957731), .Z(n_35627));
	notech_or4 i_210032830(.A(code_req), .B(n_61418), .C(n_61386), .D(n_17958
		), .Z(n_122157733));
	notech_nand2 i_4128428(.A(n_140057892), .B(n_122157733), .Z(n_35621));
	notech_or4 i_210432826(.A(code_req), .B(n_61418), .C(n_61386), .D(n_17959
		), .Z(n_122357735));
	notech_nand2 i_4028427(.A(n_140157893), .B(n_122357735), .Z(n_35615));
	notech_or4 i_210832822(.A(n_62841), .B(n_61419), .C(n_61386), .D(n_17960
		), .Z(n_122557737));
	notech_nand2 i_3928426(.A(n_140257894), .B(n_122557737), .Z(n_35609));
	notech_or4 i_211732818(.A(n_62841), .B(n_61419), .C(n_61386), .D(n_17961
		), .Z(n_122757739));
	notech_nand2 i_3828425(.A(n_140357895), .B(n_122757739), .Z(n_35603));
	notech_or4 i_212232814(.A(code_req), .B(n_61419), .C(n_61386), .D(n_17962
		), .Z(n_122957741));
	notech_nand2 i_3728424(.A(n_140457896), .B(n_122957741), .Z(n_35597));
	notech_or4 i_212632810(.A(code_req), .B(n_61419), .C(n_61386), .D(n_17963
		), .Z(n_123157743));
	notech_nand2 i_3628423(.A(n_140557897), .B(n_123157743), .Z(n_35591));
	notech_or4 i_213032806(.A(code_req), .B(n_61419), .C(n_61386), .D(n_17964
		), .Z(n_123757745));
	notech_nand2 i_3528422(.A(n_140657898), .B(n_123757745), .Z(n_35585));
	notech_or4 i_213432802(.A(code_req), .B(n_61418), .C(n_61386), .D(n_17965
		), .Z(n_123957747));
	notech_nand2 i_3428421(.A(n_140757899), .B(n_123957747), .Z(n_35579));
	notech_or4 i_213832798(.A(code_req), .B(n_61419), .C(n_61386), .D(n_17966
		), .Z(n_124157749));
	notech_nand2 i_3328420(.A(n_140857900), .B(n_124157749), .Z(n_35573));
	notech_or4 i_214232794(.A(n_62841), .B(n_61419), .C(n_61386), .D(n_17967
		), .Z(n_124357751));
	notech_nand2 i_3228419(.A(n_140957901), .B(n_124357751), .Z(n_35567));
	notech_or4 i_214632790(.A(code_req), .B(n_61421), .C(n_61386), .D(n_17968
		), .Z(n_124557753));
	notech_nand2 i_3128418(.A(n_141057902), .B(n_124557753), .Z(n_35561));
	notech_or4 i_215032786(.A(code_req), .B(n_61424), .C(n_61388), .D(n_17969
		), .Z(n_124757755));
	notech_nand2 i_3028417(.A(n_141157903), .B(n_124757755), .Z(n_35555));
	notech_or4 i_215432782(.A(n_62846), .B(n_61424), .C(n_61392), .D(n_17970
		), .Z(n_124957757));
	notech_nand2 i_2928416(.A(n_141257904), .B(n_124957757), .Z(n_35549));
	notech_or4 i_216232774(.A(n_62849), .B(n_61424), .C(n_61392), .D(n_17971
		), .Z(n_125157759));
	notech_nand2 i_2728414(.A(n_141357905), .B(n_125157759), .Z(n_35537));
	notech_or4 i_216632770(.A(n_62849), .B(n_61424), .C(n_61392), .D(n_17972
		), .Z(n_125357761));
	notech_nand2 i_2628413(.A(n_141457906), .B(n_125357761), .Z(n_35531));
	notech_or4 i_217032766(.A(n_62849), .B(n_61424), .C(n_61392), .D(n_17973
		), .Z(n_125557763));
	notech_nand2 i_2528412(.A(n_141557907), .B(n_125557763), .Z(n_35525));
	notech_or4 i_217432762(.A(n_62849), .B(n_61424), .C(n_61392), .D(n_17974
		), .Z(n_125757765));
	notech_nand2 i_2428411(.A(n_141657908), .B(n_125757765), .Z(n_35519));
	notech_or4 i_217832758(.A(n_62849), .B(n_61424), .C(n_61392), .D(n_17975
		), .Z(n_125957767));
	notech_nand2 i_2328410(.A(n_141757909), .B(n_125957767), .Z(n_35513));
	notech_or4 i_218232754(.A(n_62849), .B(n_61424), .C(n_61392), .D(n_17976
		), .Z(n_126157769));
	notech_nand2 i_2228409(.A(n_141857910), .B(n_126157769), .Z(n_35507));
	notech_or4 i_218632750(.A(n_62849), .B(n_61426), .C(n_61392), .D(n_17977
		), .Z(n_126357771));
	notech_nand2 i_2128408(.A(n_141957911), .B(n_126357771), .Z(n_35501));
	notech_or4 i_219832738(.A(n_62849), .B(n_61426), .C(n_61394), .D(n_17978
		), .Z(n_126557773));
	notech_nand2 i_1828405(.A(n_142057912), .B(n_126557773), .Z(n_35483));
	notech_or4 i_220232734(.A(n_62849), .B(n_61426), .C(n_61394), .D(n_17979
		), .Z(n_126757775));
	notech_nand2 i_1728404(.A(n_142157913), .B(n_126757775), .Z(n_35477));
	notech_or4 i_220632730(.A(n_62849), .B(n_61426), .C(n_61394), .D(n_17980
		), .Z(n_126957777));
	notech_nand2 i_1628403(.A(n_142257914), .B(n_126957777), .Z(n_35471));
	notech_or4 i_221032726(.A(n_62852), .B(n_61424), .C(n_61394), .D(n_17981
		), .Z(n_127157779));
	notech_nand2 i_1528402(.A(n_142357915), .B(n_127157779), .Z(n_35465));
	notech_or4 i_222632710(.A(n_62852), .B(n_61424), .C(n_61392), .D(n_17982
		), .Z(n_127357781));
	notech_nand2 i_1128398(.A(n_142457916), .B(n_127357781), .Z(n_35441));
	notech_or4 i_223032706(.A(n_62849), .B(n_61424), .C(n_61392), .D(n_17983
		), .Z(n_127557783));
	notech_nand2 i_1028397(.A(n_142557917), .B(n_127557783), .Z(n_35435));
	notech_or4 i_223432702(.A(n_62849), .B(n_61424), .C(n_61392), .D(n_17984
		), .Z(n_127757785));
	notech_nand2 i_928396(.A(n_142657918), .B(n_127757785), .Z(n_35429));
	notech_or4 i_223832698(.A(n_62849), .B(n_61424), .C(n_61392), .D(n_17985
		), .Z(n_127957787));
	notech_nand2 i_828395(.A(n_142757919), .B(n_127957787), .Z(n_35423));
	notech_or4 i_224232694(.A(n_62849), .B(n_61421), .C(n_61392), .D(n_17986
		), .Z(n_128157789));
	notech_nand2 i_728394(.A(n_142857920), .B(n_128157789), .Z(n_35417));
	notech_or4 i_224632690(.A(n_62847), .B(n_61421), .C(n_61390), .D(n_17987
		), .Z(n_128357791));
	notech_nand2 i_628393(.A(n_142957921), .B(n_128357791), .Z(n_35411));
	notech_or4 i_225032686(.A(n_62847), .B(n_61421), .C(n_61390), .D(n_17988
		), .Z(n_128557793));
	notech_nand2 i_528392(.A(n_143057922), .B(n_128557793), .Z(n_35405));
	notech_or4 i_226232674(.A(n_62847), .B(n_61421), .C(n_61390), .D(n_17989
		), .Z(n_128857795));
	notech_nand2 i_228389(.A(n_143157923), .B(n_128857795), .Z(n_35387));
	notech_or4 i_226632670(.A(n_62847), .B(n_61421), .C(n_61390), .D(n_17990
		), .Z(n_129357797));
	notech_nand2 i_128388(.A(n_143257924), .B(n_129357797), .Z(n_35381));
	notech_or2 i_1634906(.A(n_61567), .B(n_17293), .Z(n_14278717));
	notech_nor2 i_1734905(.A(n_62847), .B(n_61421), .Z(n_14238713));
	notech_and4 i_4434882(.A(tagV[2]), .B(n_36941), .C(n_17680), .D(n_17681)
		, .Z(n_130357803));
	notech_ao3 i_4234924(.A(n_17301), .B(n_61153), .C(n_62846), .Z(n_14128702
		));
	notech_or4 i_1934903(.A(n_62846), .B(pg_fault), .C(n_61421), .D(n_61388)
		, .Z(n_130657804));
	notech_and2 i_3434889(.A(n_61567), .B(n_8293), .Z(n_130757805));
	notech_ao4 i_174233188(.A(n_61359), .B(n_17860), .C(n_61153), .D(n_17675
		), .Z(n_130957807));
	notech_ao4 i_174633184(.A(n_61329), .B(n_17859), .C(n_61153), .D(n_17673
		), .Z(n_131257808));
	notech_ao4 i_175033180(.A(n_61329), .B(n_17858), .C(n_61153), .D(n_17671
		), .Z(n_131357809));
	notech_ao4 i_175433176(.A(n_61329), .B(n_17857), .C(n_61157), .D(n_17669
		), .Z(n_131657810));
	notech_ao4 i_175833172(.A(n_61329), .B(n_17856), .C(n_61157), .D(n_17667
		), .Z(n_131757811));
	notech_ao4 i_176233168(.A(n_61329), .B(n_17855), .C(n_61157), .D(n_17665
		), .Z(n_131957812));
	notech_ao4 i_176633164(.A(n_61359), .B(n_17854), .C(n_61157), .D(n_17663
		), .Z(n_132057813));
	notech_ao4 i_177033160(.A(n_61329), .B(n_17853), .C(n_61157), .D(n_17661
		), .Z(n_132257814));
	notech_ao4 i_177433156(.A(n_61329), .B(n_17852), .C(n_61157), .D(n_17659
		), .Z(n_132357815));
	notech_ao4 i_177833152(.A(n_61363), .B(n_17851), .C(n_61157), .D(n_17657
		), .Z(n_132457816));
	notech_ao4 i_178233148(.A(n_61363), .B(n_17850), .C(n_61157), .D(n_17655
		), .Z(n_132557817));
	notech_ao4 i_178633144(.A(n_61363), .B(n_17849), .C(n_61151), .D(n_17653
		), .Z(n_132657818));
	notech_ao4 i_179433136(.A(n_61363), .B(n_17847), .C(n_61151), .D(n_17649
		), .Z(n_132757819));
	notech_ao4 i_179833132(.A(n_61363), .B(n_17846), .C(n_61151), .D(n_17647
		), .Z(n_132857820));
	notech_ao4 i_180233128(.A(n_61363), .B(n_17845), .C(n_61151), .D(n_17645
		), .Z(n_132957821));
	notech_ao4 i_180633124(.A(n_61363), .B(n_17844), .C(n_61151), .D(n_17643
		), .Z(n_133057822));
	notech_ao4 i_181033120(.A(n_61363), .B(n_17843), .C(n_61151), .D(n_17641
		), .Z(n_133157823));
	notech_ao4 i_181433116(.A(n_61359), .B(n_17842), .C(n_61151), .D(n_17639
		), .Z(n_133257824));
	notech_ao4 i_181833112(.A(n_61359), .B(n_17841), .C(n_61151), .D(n_17637
		), .Z(n_133357825));
	notech_ao4 i_182233108(.A(n_61359), .B(n_17840), .C(n_61151), .D(n_17635
		), .Z(n_133457826));
	notech_ao4 i_182633104(.A(n_61359), .B(n_17839), .C(n_61153), .D(n_17633
		), .Z(n_133557827));
	notech_ao4 i_183033100(.A(n_61363), .B(n_17838), .C(n_61153), .D(n_17631
		), .Z(n_133657828));
	notech_ao4 i_183433096(.A(n_61363), .B(n_17837), .C(n_61153), .D(n_17629
		), .Z(n_133757829));
	notech_ao4 i_183833092(.A(n_61359), .B(n_17836), .C(n_61153), .D(n_17627
		), .Z(n_133857830));
	notech_ao4 i_184233088(.A(n_61359), .B(n_17835), .C(n_61151), .D(n_17625
		), .Z(n_133957831));
	notech_ao4 i_184733083(.A(n_61151), .B(n_17623), .C(n_61349), .D(n_17834
		), .Z(n_134057832));
	notech_ao4 i_185133079(.A(n_61349), .B(n_17833), .C(n_61153), .D(n_17621
		), .Z(n_134157833));
	notech_ao4 i_185633074(.A(n_61151), .B(n_17619), .C(n_61344), .D(n_17832
		), .Z(n_134257834));
	notech_ao4 i_186033070(.A(n_61349), .B(n_17831), .C(n_61160), .D(n_17617
		), .Z(n_134357835));
	notech_ao4 i_186533065(.A(n_61160), .B(n_17615), .C(n_61349), .D(n_17830
		), .Z(n_134457836));
	notech_ao4 i_186933061(.A(n_61349), .B(n_17829), .C(n_61160), .D(n_17613
		), .Z(n_134557837));
	notech_ao4 i_187433056(.A(n_61160), .B(n_17611), .C(n_61349), .D(n_17828
		), .Z(n_134657838));
	notech_ao4 i_187933051(.A(n_61158), .B(n_17609), .C(n_61349), .D(n_17827
		), .Z(n_134757839));
	notech_ao4 i_188333047(.A(n_61344), .B(n_17826), .C(n_61158), .D(n_17607
		), .Z(n_134857840));
	notech_ao4 i_188833042(.A(n_61160), .B(n_17605), .C(n_61344), .D(n_17825
		), .Z(n_134957841));
	notech_ao4 i_189333037(.A(n_61158), .B(n_17603), .C(n_61344), .D(n_17824
		), .Z(n_135057842));
	notech_ao4 i_190333027(.A(n_61160), .B(n_17599), .C(n_61344), .D(n_17822
		), .Z(n_135157843));
	notech_ao4 i_190833022(.A(n_61160), .B(n_17597), .C(n_61344), .D(n_17821
		), .Z(n_135257844));
	notech_ao4 i_191333017(.A(n_61160), .B(n_17595), .C(n_61344), .D(n_17820
		), .Z(n_135357845));
	notech_ao4 i_191833012(.A(n_61160), .B(n_17593), .C(n_61344), .D(n_17819
		), .Z(n_135457846));
	notech_ao4 i_192233008(.A(n_61344), .B(n_17818), .C(n_61160), .D(n_17591
		), .Z(n_135557847));
	notech_ao4 i_192633004(.A(n_61329), .B(n_17817), .C(n_61160), .D(n_17589
		), .Z(n_135657848));
	notech_ao4 i_193033000(.A(n_61329), .B(n_17816), .C(n_61160), .D(n_17587
		), .Z(n_135757849));
	notech_ao4 i_193432996(.A(n_61329), .B(n_17815), .C(n_61160), .D(n_17585
		), .Z(n_135857850));
	notech_ao4 i_193832992(.A(n_61329), .B(n_17814), .C(n_61160), .D(n_17583
		), .Z(n_135957851));
	notech_ao4 i_194232988(.A(n_61329), .B(n_17813), .C(n_61157), .D(n_17581
		), .Z(n_136057852));
	notech_ao4 i_194632984(.A(n_61329), .B(n_17812), .C(n_61157), .D(n_17579
		), .Z(n_136157853));
	notech_ao4 i_195032980(.A(n_61329), .B(n_17811), .C(n_61158), .D(n_17577
		), .Z(n_136257854));
	notech_ao4 i_195432976(.A(n_61329), .B(n_17810), .C(n_61158), .D(n_17575
		), .Z(n_136357855));
	notech_ao4 i_195832972(.A(n_61349), .B(n_17809), .C(n_61157), .D(n_17573
		), .Z(n_136457856));
	notech_ao4 i_196232968(.A(n_61349), .B(n_17808), .C(n_61157), .D(n_17571
		), .Z(n_136557857));
	notech_ao4 i_196632964(.A(n_61349), .B(n_17807), .C(n_61157), .D(n_17569
		), .Z(n_136657858));
	notech_ao4 i_197032960(.A(n_61349), .B(n_17806), .C(n_61157), .D(n_17567
		), .Z(n_136757859));
	notech_ao4 i_197432956(.A(n_61349), .B(n_17805), .C(n_61158), .D(n_17565
		), .Z(n_136857860));
	notech_ao4 i_197832952(.A(n_61349), .B(n_17804), .C(n_61158), .D(n_17563
		), .Z(n_136957861));
	notech_ao4 i_198232948(.A(n_61349), .B(n_17803), .C(n_61158), .D(n_17561
		), .Z(n_137057862));
	notech_ao4 i_198632944(.A(n_61349), .B(n_17802), .C(n_61158), .D(n_17559
		), .Z(n_137157863));
	notech_ao4 i_199032940(.A(n_61363), .B(n_17801), .C(n_61158), .D(n_17557
		), .Z(n_137257864));
	notech_ao4 i_199432936(.A(n_61377), .B(n_17800), .C(n_61158), .D(n_17555
		), .Z(n_137357865));
	notech_ao4 i_199832932(.A(n_61377), .B(n_17799), .C(n_61158), .D(n_17553
		), .Z(n_137457866));
	notech_ao4 i_200232928(.A(n_61377), .B(n_17798), .C(n_61158), .D(n_17551
		), .Z(n_137557867));
	notech_ao4 i_200632924(.A(n_61377), .B(n_17797), .C(n_61158), .D(n_17549
		), .Z(n_137657868));
	notech_ao4 i_201032920(.A(n_61377), .B(n_17796), .C(n_61151), .D(n_17547
		), .Z(n_137757869));
	notech_ao4 i_201432916(.A(n_61377), .B(n_17795), .C(n_61151), .D(n_17545
		), .Z(n_137857870));
	notech_ao4 i_201832912(.A(n_61377), .B(n_17794), .C(n_61145), .D(n_17543
		), .Z(n_137957871));
	notech_ao4 i_202232908(.A(n_61377), .B(n_17793), .C(n_61151), .D(n_17541
		), .Z(n_138057872));
	notech_ao4 i_202632904(.A(n_61377), .B(n_17792), .C(n_61151), .D(n_17539
		), .Z(n_138157873));
	notech_ao4 i_203032900(.A(n_61377), .B(n_17791), .C(n_61153), .D(n_17537
		), .Z(n_138257874));
	notech_ao4 i_203432896(.A(n_61372), .B(n_17790), .C(n_61151), .D(n_17535
		), .Z(n_138357875));
	notech_ao4 i_203832892(.A(n_61372), .B(n_17789), .C(n_61151), .D(n_17533
		), .Z(n_138457876));
	notech_ao4 i_204232888(.A(n_61377), .B(n_17788), .C(n_61145), .D(n_17531
		), .Z(n_138557877));
	notech_ao4 i_204632884(.A(n_61377), .B(n_17787), .C(n_61145), .D(n_17529
		), .Z(n_138657878));
	notech_ao4 i_205032880(.A(n_61377), .B(n_17786), .C(n_61145), .D(n_17527
		), .Z(n_138757879));
	notech_ao4 i_205432876(.A(n_61377), .B(n_17785), .C(n_61145), .D(n_17525
		), .Z(n_138857880));
	notech_ao4 i_205832872(.A(n_14228712), .B(n_17784), .C(n_61145), .D(n_17523
		), .Z(n_138957881));
	notech_ao4 i_206232868(.A(n_14228712), .B(n_17783), .C(n_61145), .D(n_17521
		), .Z(n_139057882));
	notech_ao4 i_206632864(.A(n_14228712), .B(n_17782), .C(n_61145), .D(n_17519
		), .Z(n_139157883));
	notech_ao4 i_207032860(.A(n_14228712), .B(n_17781), .C(n_61145), .D(n_17517
		), .Z(n_139257884));
	notech_ao4 i_207432856(.A(n_14228712), .B(n_17780), .C(n_61145), .D(n_17515
		), .Z(n_139357885));
	notech_ao4 i_207832852(.A(n_14228712), .B(n_17779), .C(n_61158), .D(n_17513
		), .Z(n_139457886));
	notech_ao4 i_208232848(.A(n_14228712), .B(n_17778), .C(n_61158), .D(n_17511
		), .Z(n_139557887));
	notech_ao4 i_208632844(.A(n_14228712), .B(n_17777), .C(n_61160), .D(n_17509
		), .Z(n_139657888));
	notech_ao4 i_209032840(.A(n_14228712), .B(n_17776), .C(n_61160), .D(n_17507
		), .Z(n_139757889));
	notech_ao4 i_209432836(.A(n_14228712), .B(n_17775), .C(n_61158), .D(n_17505
		), .Z(n_139857890));
	notech_ao4 i_209832832(.A(n_61377), .B(n_17774), .C(n_61158), .D(n_17503
		), .Z(n_139957891));
	notech_ao4 i_210232828(.A(n_14228712), .B(n_17773), .C(n_61158), .D(n_17501
		), .Z(n_140057892));
	notech_ao4 i_210632824(.A(n_14228712), .B(n_17772), .C(n_61158), .D(n_17499
		), .Z(n_140157893));
	notech_ao4 i_211032820(.A(n_14228712), .B(n_17771), .C(n_61160), .D(n_17497
		), .Z(n_140257894));
	notech_ao4 i_212032816(.A(n_14228712), .B(n_17770), .C(n_61153), .D(n_17495
		), .Z(n_140357895));
	notech_ao4 i_212432812(.A(n_14228712), .B(n_17769), .C(n_61153), .D(n_17493
		), .Z(n_140457896));
	notech_ao4 i_212832808(.A(n_61368), .B(n_17768), .C(n_61153), .D(n_17491
		), .Z(n_140557897));
	notech_ao4 i_213232804(.A(n_61368), .B(n_17767), .C(n_61153), .D(n_17489
		), .Z(n_140657898));
	notech_ao4 i_213632800(.A(n_61368), .B(n_17766), .C(n_61160), .D(n_17487
		), .Z(n_140757899));
	notech_ao4 i_214032796(.A(n_61368), .B(n_17765), .C(n_61160), .D(n_17485
		), .Z(n_140857900));
	notech_ao4 i_214432792(.A(n_61368), .B(n_17764), .C(n_61153), .D(n_17483
		), .Z(n_140957901));
	notech_ao4 i_214832788(.A(n_61368), .B(n_17763), .C(n_61160), .D(n_17481
		), .Z(n_141057902));
	notech_ao4 i_215232784(.A(n_61368), .B(n_17762), .C(n_61148), .D(n_17479
		), .Z(n_141157903));
	notech_ao4 i_215632780(.A(n_61368), .B(n_17761), .C(n_61148), .D(n_17477
		), .Z(n_141257904));
	notech_ao4 i_216432772(.A(n_61363), .B(n_17759), .C(n_61148), .D(n_17473
		), .Z(n_141357905));
	notech_ao4 i_216832768(.A(n_61363), .B(n_17758), .C(n_61148), .D(n_17471
		), .Z(n_141457906));
	notech_ao4 i_217232764(.A(n_61363), .B(n_17757), .C(n_61148), .D(n_17469
		), .Z(n_141557907));
	notech_ao4 i_217632760(.A(n_61363), .B(n_17756), .C(n_61146), .D(n_17467
		), .Z(n_141657908));
	notech_ao4 i_218032756(.A(n_61368), .B(n_17755), .C(n_61148), .D(n_17465
		), .Z(n_141757909));
	notech_ao4 i_218432752(.A(n_61368), .B(n_17754), .C(n_61148), .D(n_17463
		), .Z(n_141857910));
	notech_ao4 i_218832748(.A(n_61368), .B(n_17753), .C(n_61148), .D(n_17461
		), .Z(n_141957911));
	notech_ao4 i_220032736(.A(n_61368), .B(n_17750), .C(n_61148), .D(n_17455
		), .Z(n_142057912));
	notech_ao4 i_220432732(.A(n_61372), .B(n_17749), .C(n_61148), .D(n_17453
		), .Z(n_142157913));
	notech_ao4 i_220832728(.A(n_61372), .B(n_17748), .C(n_61151), .D(n_17451
		), .Z(n_142257914));
	notech_ao4 i_221232724(.A(n_61372), .B(n_17747), .C(n_61151), .D(n_17449
		), .Z(n_142357915));
	notech_ao4 i_222832708(.A(n_61372), .B(n_17743), .C(n_61148), .D(n_17441
		), .Z(n_142457916));
	notech_ao4 i_223232704(.A(n_61372), .B(n_17742), .C(n_61148), .D(n_17439
		), .Z(n_142557917));
	notech_ao4 i_223632700(.A(n_61372), .B(n_17741), .C(n_61148), .D(n_17437
		), .Z(n_142657918));
	notech_ao4 i_224032696(.A(n_61372), .B(n_17740), .C(n_61148), .D(n_17435
		), .Z(n_142757919));
	notech_ao4 i_224432692(.A(n_61372), .B(n_17739), .C(n_61146), .D(n_17433
		), .Z(n_142857920));
	notech_ao4 i_224832688(.A(n_61368), .B(n_17738), .C(n_61146), .D(n_17431
		), .Z(n_142957921));
	notech_ao4 i_225232684(.A(n_61372), .B(n_17737), .C(n_61146), .D(n_17429
		), .Z(n_143057922));
	notech_ao4 i_226432672(.A(n_61368), .B(n_17734), .C(n_61146), .D(n_17423
		), .Z(n_143157923));
	notech_ao4 i_226832668(.A(n_61368), .B(n_17733), .C(n_61145), .D(n_17421
		), .Z(n_143257924));
	notech_nand3 i_3581539(.A(n_59940), .B(queue[7]), .C(n_59669), .Z(n_143357925
		));
	notech_or2 i_3681554(.A(n_59947), .B(n_17322), .Z(n_144857940));
	notech_nand3 i_824974(.A(n_232558817), .B(n_231858810), .C(n_143357925),
		 .Z(squeue[7]));
	notech_nand3 i_9981555(.A(n_59669), .B(n_59938), .C(queue[29]), .Z(n_144957941
		));
	notech_or2 i_10081570(.A(n_59947), .B(n_17344), .Z(n_146457956));
	notech_nand3 i_3024996(.A(n_233958831), .B(n_233258824), .C(n_144957941)
		, .Z(squeue[29]));
	notech_nand3 i_13081571(.A(n_59669), .B(n_59938), .C(queue[37]), .Z(n_146557957
		));
	notech_or2 i_13181586(.A(n_59947), .B(n_17352), .Z(n_148057972));
	notech_nand3 i_3825004(.A(n_235358845), .B(n_234658838), .C(n_146557957)
		, .Z(squeue[37]));
	notech_nand3 i_19281587(.A(n_59669), .B(n_59938), .C(queue[55]), .Z(n_148157973
		));
	notech_or2 i_19381602(.A(n_59947), .B(n_17370), .Z(n_149657988));
	notech_nand3 i_5625022(.A(n_236758859), .B(n_236058852), .C(n_148157973)
		, .Z(squeue[55]));
	notech_nand3 i_22381603(.A(n_59667), .B(n_59938), .C(queue[56]), .Z(n_149757989
		));
	notech_or2 i_22481618(.A(n_59947), .B(n_17371), .Z(n_151258004));
	notech_nand3 i_5725023(.A(n_238158873), .B(n_237458866), .C(n_149757989)
		, .Z(squeue[56]));
	notech_nand3 i_25481619(.A(n_59667), .B(n_59938), .C(queue[57]), .Z(n_151358005
		));
	notech_or2 i_25581634(.A(n_59947), .B(n_17372), .Z(n_152858020));
	notech_nand3 i_5825024(.A(n_239558887), .B(n_238858880), .C(n_151358005)
		, .Z(squeue[57]));
	notech_nand3 i_28581635(.A(n_59667), .B(n_59938), .C(queue[58]), .Z(n_152958021
		));
	notech_or2 i_28681650(.A(n_59947), .B(n_17373), .Z(n_154458036));
	notech_nand3 i_5925025(.A(n_240958901), .B(n_240258894), .C(n_152958021)
		, .Z(squeue[58]));
	notech_nand3 i_31681651(.A(n_59667), .B(n_59938), .C(queue[59]), .Z(n_154558037
		));
	notech_or2 i_31781666(.A(n_59947), .B(n_17374), .Z(n_156058052));
	notech_nand3 i_6025026(.A(n_242358915), .B(n_241658908), .C(n_154558037)
		, .Z(squeue[59]));
	notech_nand3 i_37881667(.A(n_59667), .B(n_59938), .C(queue[61]), .Z(n_156158053
		));
	notech_or2 i_37981682(.A(n_59944), .B(n_17376), .Z(n_157658068));
	notech_nand3 i_6225028(.A(n_243758929), .B(n_243058922), .C(n_156158053)
		, .Z(squeue[61]));
	notech_nand3 i_44081683(.A(n_59667), .B(n_59938), .C(queue[63]), .Z(n_157758069
		));
	notech_or2 i_44181698(.A(n_59944), .B(n_17378), .Z(n_159258084));
	notech_nand3 i_6425030(.A(n_245158943), .B(n_244458936), .C(n_157758069)
		, .Z(squeue[63]));
	notech_nand3 i_50281699(.A(n_59667), .B(n_59938), .C(queue[66]), .Z(n_159358085
		));
	notech_or2 i_50381714(.A(n_59944), .B(n_17381), .Z(n_160858100));
	notech_nand3 i_6725033(.A(n_246558957), .B(n_245858950), .C(n_159358085)
		, .Z(squeue[66]));
	notech_nand3 i_53381715(.A(n_59667), .B(n_59940), .C(queue[67]), .Z(n_160958101
		));
	notech_or2 i_53481730(.A(n_59944), .B(n_17382), .Z(n_162458116));
	notech_nand3 i_6825034(.A(n_247958971), .B(n_247258964), .C(n_160958101)
		, .Z(squeue[67]));
	notech_nand3 i_59581731(.A(n_59667), .B(n_59938), .C(queue[69]), .Z(n_162558117
		));
	notech_or2 i_59681746(.A(n_59944), .B(n_17384), .Z(n_164058132));
	notech_nand3 i_7025036(.A(n_249358985), .B(n_248658978), .C(n_162558117)
		, .Z(squeue[69]));
	notech_nand3 i_65781747(.A(n_59667), .B(n_59938), .C(queue[71]), .Z(n_164158133
		));
	notech_or2 i_65881762(.A(n_59944), .B(n_17386), .Z(n_165658148));
	notech_nand3 i_7225038(.A(n_250758999), .B(n_250058992), .C(n_164158133)
		, .Z(squeue[71]));
	notech_nand3 i_68881763(.A(n_59667), .B(n_59938), .C(queue[72]), .Z(n_165758149
		));
	notech_or2 i_68981778(.A(n_59944), .B(n_17387), .Z(n_167258164));
	notech_nand3 i_7325039(.A(n_252159013), .B(n_251459006), .C(n_165758149)
		, .Z(squeue[72]));
	notech_nand3 i_71981779(.A(n_59667), .B(n_59938), .C(queue[73]), .Z(n_167358165
		));
	notech_or2 i_72081794(.A(n_59944), .B(n_17388), .Z(n_168858180));
	notech_nand3 i_7425040(.A(n_253559027), .B(n_252859020), .C(n_167358165)
		, .Z(squeue[73]));
	notech_nand3 i_75081795(.A(n_59667), .B(n_59938), .C(queue[74]), .Z(n_168958181
		));
	notech_or2 i_75181810(.A(n_59945), .B(n_17389), .Z(n_170458196));
	notech_nand3 i_7525041(.A(n_254959041), .B(n_254259034), .C(n_168958181)
		, .Z(squeue[74]));
	notech_nand3 i_84381811(.A(n_59667), .B(n_59926), .C(queue[77]), .Z(n_170558197
		));
	notech_or2 i_84481826(.A(n_59945), .B(n_17392), .Z(n_172058212));
	notech_nand3 i_7825044(.A(n_256359055), .B(n_255659048), .C(n_170558197)
		, .Z(squeue[77]));
	notech_nand3 i_90581827(.A(n_59667), .B(n_59926), .C(queue[79]), .Z(n_172158213
		));
	notech_or2 i_90681842(.A(n_59945), .B(n_17394), .Z(n_173658228));
	notech_nand3 i_8025046(.A(n_257759069), .B(n_257059062), .C(n_172158213)
		, .Z(squeue[79]));
	notech_nand3 i_93681843(.A(n_59667), .B(n_59926), .C(queue[80]), .Z(n_173758229
		));
	notech_or2 i_93781858(.A(n_59945), .B(n_17395), .Z(n_175258244));
	notech_nand3 i_8125047(.A(n_259159083), .B(n_258459076), .C(n_173758229)
		, .Z(squeue[80]));
	notech_nand3 i_96781859(.A(n_59654), .B(n_59926), .C(queue[81]), .Z(n_175358245
		));
	notech_or2 i_96881874(.A(n_59945), .B(n_17396), .Z(n_176858260));
	notech_nand3 i_8225048(.A(n_260559097), .B(n_259859090), .C(n_175358245)
		, .Z(squeue[81]));
	notech_nand3 i_99881875(.A(n_59654), .B(n_59926), .C(queue[82]), .Z(n_176958261
		));
	notech_or2 i_99981890(.A(n_59945), .B(n_17397), .Z(n_178458276));
	notech_nand3 i_8325049(.A(n_261959111), .B(n_261259104), .C(n_176958261)
		, .Z(squeue[82]));
	notech_nand3 i_102981891(.A(n_59654), .B(n_59926), .C(queue[83]), .Z(n_178558277
		));
	notech_or2 i_103081906(.A(n_59945), .B(n_17398), .Z(n_180058292));
	notech_nand3 i_8425050(.A(n_263359125), .B(n_262659118), .C(n_178558277)
		, .Z(squeue[83]));
	notech_nand3 i_109181907(.A(n_59654), .B(n_59926), .C(queue[85]), .Z(n_180158293
		));
	notech_or2 i_109281922(.A(n_59945), .B(n_17400), .Z(n_181658308));
	notech_nand3 i_8625052(.A(n_264759139), .B(n_264059132), .C(n_180158293)
		, .Z(squeue[85]));
	notech_nand3 i_115381923(.A(n_59654), .B(n_59926), .C(queue[87]), .Z(n_181758309
		));
	notech_or2 i_115481938(.A(n_59950), .B(n_17402), .Z(n_183258324));
	notech_nand3 i_8825054(.A(n_266159153), .B(n_265459146), .C(n_181758309)
		, .Z(squeue[87]));
	notech_nand3 i_118481939(.A(n_59654), .B(n_59928), .C(queue[88]), .Z(n_183358325
		));
	notech_or2 i_118581954(.A(n_59950), .B(n_17403), .Z(n_184858340));
	notech_nand3 i_8925055(.A(n_267559167), .B(n_266859160), .C(n_183358325)
		, .Z(squeue[88]));
	notech_nand3 i_121581955(.A(n_59654), .B(n_59928), .C(queue[89]), .Z(n_184958341
		));
	notech_or2 i_121681970(.A(n_59950), .B(n_17404), .Z(n_186458356));
	notech_nand3 i_9025056(.A(n_268959181), .B(n_268259174), .C(n_184958341)
		, .Z(squeue[89]));
	notech_nand3 i_124681971(.A(n_59654), .B(n_59928), .C(queue[90]), .Z(n_186558357
		));
	notech_or2 i_124781986(.A(n_59950), .B(n_17405), .Z(n_188058372));
	notech_nand3 i_9125057(.A(n_270359195), .B(n_269659188), .C(n_186558357)
		, .Z(squeue[90]));
	notech_nand3 i_127781987(.A(n_59654), .B(n_59928), .C(queue[91]), .Z(n_188158373
		));
	notech_or2 i_127882002(.A(n_59950), .B(n_17406), .Z(n_189658388));
	notech_nand3 i_9225058(.A(n_271759209), .B(n_271059202), .C(n_188158373)
		, .Z(squeue[91]));
	notech_nand3 i_133982003(.A(n_59654), .B(n_59928), .C(queue[93]), .Z(n_189758389
		));
	notech_or2 i_134082018(.A(n_59950), .B(n_17408), .Z(n_191258404));
	notech_nand3 i_9425060(.A(n_273159223), .B(n_272459216), .C(n_189758389)
		, .Z(squeue[93]));
	notech_nand3 i_140182019(.A(n_59654), .B(n_59926), .C(queue[95]), .Z(n_191358405
		));
	notech_or2 i_140282034(.A(n_59950), .B(n_17410), .Z(n_192858420));
	notech_nand3 i_9625062(.A(n_274559237), .B(n_273859230), .C(n_191358405)
		, .Z(squeue[95]));
	notech_nand3 i_143282035(.A(n_59654), .B(n_59928), .C(queue[96]), .Z(n_192958421
		));
	notech_or2 i_143382050(.A(n_59950), .B(n_17411), .Z(n_194458436));
	notech_nand3 i_9725063(.A(n_275959251), .B(n_275259244), .C(n_192958421)
		, .Z(squeue[96]));
	notech_nand3 i_146382051(.A(n_59654), .B(n_59928), .C(queue[97]), .Z(n_194558437
		));
	notech_or2 i_146482066(.A(n_59952), .B(n_17412), .Z(n_196058452));
	notech_nand3 i_9825064(.A(n_277359265), .B(n_276659258), .C(n_194558437)
		, .Z(squeue[97]));
	notech_nand3 i_149482067(.A(n_59654), .B(n_59926), .C(queue[98]), .Z(n_196158453
		));
	notech_or2 i_149582082(.A(n_59952), .B(n_17413), .Z(n_197658468));
	notech_nand3 i_9925065(.A(n_278759279), .B(n_278059272), .C(n_196158453)
		, .Z(squeue[98]));
	notech_nand3 i_152582083(.A(n_59654), .B(n_59925), .C(queue[99]), .Z(n_197758469
		));
	notech_or2 i_152682098(.A(n_59952), .B(n_17414), .Z(n_199258484));
	notech_nand3 i_10025066(.A(n_280159293), .B(n_279459286), .C(n_197758469
		), .Z(squeue[99]));
	notech_nand3 i_1587(.A(n_59654), .B(n_59925), .C(queue[101]), .Z(n_199358485
		));
	notech_or2 i_1588(.A(n_59952), .B(n_17416), .Z(n_200858500));
	notech_nand3 i_10225068(.A(n_281559307), .B(n_280859300), .C(n_199358485
		), .Z(squeue[101]));
	notech_nand3 i_1649(.A(n_59652), .B(n_59925), .C(queue[103]), .Z(n_200958501
		));
	notech_or2 i_1650(.A(n_59952), .B(n_17418), .Z(n_202458516));
	notech_nand3 i_10425070(.A(n_282959321), .B(n_282259314), .C(n_200958501
		), .Z(squeue[103]));
	notech_nand3 i_1680(.A(n_59652), .B(n_59925), .C(queue[104]), .Z(n_202558517
		));
	notech_or2 i_1681(.A(n_59950), .B(n_17421), .Z(n_204058532));
	notech_nand3 i_10525071(.A(n_284359335), .B(n_283659328), .C(n_202558517
		), .Z(squeue[104]));
	notech_nand3 i_1711(.A(n_59652), .B(n_59925), .C(queue[105]), .Z(n_204158533
		));
	notech_or2 i_1712(.A(n_59952), .B(n_17423), .Z(n_205658548));
	notech_nand3 i_10625072(.A(n_285759349), .B(n_285059342), .C(n_204158533
		), .Z(squeue[105]));
	notech_nand3 i_1742(.A(n_59652), .B(n_59925), .C(queue[106]), .Z(n_205758549
		));
	notech_or2 i_1743(.A(n_59952), .B(n_17425), .Z(n_207258564));
	notech_nand3 i_10725073(.A(n_287159363), .B(n_286459356), .C(n_205758549
		), .Z(squeue[106]));
	notech_nand3 i_1773(.A(n_59652), .B(n_59925), .C(queue[107]), .Z(n_207358565
		));
	notech_or2 i_1774(.A(n_59947), .B(n_17427), .Z(n_208858580));
	notech_nand3 i_10825074(.A(n_288559377), .B(n_287859370), .C(n_207358565
		), .Z(squeue[107]));
	notech_nand3 i_1835(.A(n_59652), .B(n_59925), .C(queue[109]), .Z(n_208958581
		));
	notech_or2 i_1836(.A(n_59947), .B(n_17431), .Z(n_210458596));
	notech_nand3 i_11025076(.A(n_289959391), .B(n_289259384), .C(n_208958581
		), .Z(squeue[109]));
	notech_nand3 i_1897(.A(n_59652), .B(n_59926), .C(queue[111]), .Z(n_210558597
		));
	notech_or2 i_1898(.A(n_59947), .B(n_17435), .Z(n_212058612));
	notech_nand3 i_11225078(.A(n_291359405), .B(n_290659398), .C(n_210558597
		), .Z(squeue[111]));
	notech_nand3 i_1928(.A(n_59652), .B(n_59926), .C(queue[112]), .Z(n_212158613
		));
	notech_or2 i_1929(.A(n_59947), .B(n_17437), .Z(n_213658628));
	notech_nand3 i_11325079(.A(n_292859419), .B(n_292059412), .C(n_212158613
		), .Z(squeue[112]));
	notech_nand3 i_1959(.A(n_59652), .B(n_59926), .C(queue[113]), .Z(n_213758629
		));
	notech_or2 i_1960(.A(n_59947), .B(n_17439), .Z(n_215258644));
	notech_nand3 i_11425080(.A(n_294559433), .B(n_293559426), .C(n_213758629
		), .Z(squeue[113]));
	notech_nand3 i_1990(.A(n_59652), .B(n_59926), .C(queue[114]), .Z(n_215358645
		));
	notech_or2 i_1991(.A(n_59947), .B(n_17441), .Z(n_216858660));
	notech_nand3 i_11525081(.A(n_296359447), .B(n_295559440), .C(n_215358645
		), .Z(squeue[114]));
	notech_nand3 i_2021(.A(n_59652), .B(n_59926), .C(queue[115]), .Z(n_216958661
		));
	notech_or2 i_2022(.A(n_59947), .B(n_17443), .Z(n_218458676));
	notech_nand3 i_11625082(.A(n_297859461), .B(n_297159454), .C(n_216958661
		), .Z(squeue[115]));
	notech_nand3 i_2083(.A(n_59652), .B(n_59926), .C(queue[117]), .Z(n_218558677
		));
	notech_or2 i_2084(.A(n_59947), .B(n_17447), .Z(n_220058692));
	notech_nand3 i_11825084(.A(n_299459475), .B(n_298759468), .C(n_218558677
		), .Z(squeue[117]));
	notech_nand3 i_2145(.A(n_59652), .B(n_59926), .C(queue[119]), .Z(n_220158693
		));
	notech_or2 i_2146(.A(n_59950), .B(n_17451), .Z(n_221658708));
	notech_nand3 i_12025086(.A(n_300859489), .B(n_300159482), .C(n_220158693
		), .Z(squeue[119]));
	notech_nand3 i_2176(.A(n_59652), .B(n_59926), .C(queue[120]), .Z(n_221758709
		));
	notech_or2 i_2177(.A(n_59950), .B(n_17453), .Z(n_223258724));
	notech_nand3 i_12125087(.A(n_302259503), .B(n_301559496), .C(n_221758709
		), .Z(squeue[120]));
	notech_nand3 i_2207(.A(n_59652), .B(n_59928), .C(queue[121]), .Z(n_223358725
		));
	notech_or2 i_2208(.A(n_59950), .B(n_17455), .Z(n_224858740));
	notech_nand3 i_12225088(.A(n_303659517), .B(n_302959510), .C(n_223358725
		), .Z(squeue[121]));
	notech_nand3 i_2238(.A(n_59652), .B(n_59931), .C(queue[122]), .Z(n_224958741
		));
	notech_or2 i_2239(.A(n_59950), .B(n_17457), .Z(n_226458756));
	notech_nand3 i_12325089(.A(n_305059531), .B(n_304359524), .C(n_224958741
		), .Z(squeue[122]));
	notech_nand3 i_2269(.A(n_59659), .B(n_59931), .C(queue[123]), .Z(n_226558757
		));
	notech_or2 i_2270(.A(n_59950), .B(n_17459), .Z(n_228058772));
	notech_nand3 i_12425090(.A(n_306459545), .B(n_305759538), .C(n_226558757
		), .Z(squeue[123]));
	notech_nand3 i_2331(.A(n_59659), .B(n_59931), .C(queue[125]), .Z(n_228158773
		));
	notech_or2 i_2332(.A(n_59950), .B(n_17463), .Z(n_229658788));
	notech_nand3 i_12625092(.A(n_307859559), .B(n_307159552), .C(n_228158773
		), .Z(squeue[125]));
	notech_nand3 i_2393(.A(n_59659), .B(n_59931), .C(queue[127]), .Z(n_229758789
		));
	notech_or2 i_2394(.A(n_59950), .B(n_17467), .Z(n_231258804));
	notech_nand3 i_12825094(.A(n_309259573), .B(n_308559566), .C(n_229758789
		), .Z(squeue[127]));
	notech_ao4 i_3782099(.A(n_60029), .B(n_17330), .C(n_60013), .D(n_17346),
		 .Z(n_231358805));
	notech_ao4 i_3882101(.A(n_59966), .B(n_17314), .C(n_17418), .D(n_59685),
		 .Z(n_231558807));
	notech_ao4 i_3982102(.A(n_17402), .B(n_59717), .C(n_17410), .D(n_59701),
		 .Z(n_231658808));
	notech_and4 i_4882104(.A(n_231658808), .B(n_231558807), .C(n_231358805),
		 .D(n_144857940), .Z(n_231858810));
	notech_ao4 i_4082105(.A(n_17386), .B(n_59749), .C(n_17394), .D(n_59733),
		 .Z(n_231958811));
	notech_ao4 i_4182106(.A(n_17370), .B(n_60045), .C(n_17378), .D(n_59765),
		 .Z(n_232058812));
	notech_ao4 i_4282108(.A(n_17354), .B(n_60077), .C(n_60061), .D(n_17362),
		 .Z(n_232258814));
	notech_ao4 i_4382109(.A(n_59996), .B(n_17306), .C(n_60093), .D(n_17338),
		 .Z(n_232358815));
	notech_and4 i_4982111(.A(n_232358815), .B(n_232258814), .C(n_232058812),
		 .D(n_231958811), .Z(n_232558817));
	notech_ao4 i_10182113(.A(n_60029), .B(n_17352), .C(n_60013), .D(n_17368)
		, .Z(n_232758819));
	notech_ao4 i_10282115(.A(n_59966), .B(n_17336), .C(n_59685), .D(n_17463)
		, .Z(n_232958821));
	notech_ao4 i_10382116(.A(n_59717), .B(n_17431), .C(n_59701), .D(n_17447)
		, .Z(n_233058822));
	notech_and4 i_11282118(.A(n_233058822), .B(n_232958821), .C(n_232758819)
		, .D(n_146457956), .Z(n_233258824));
	notech_ao4 i_10482119(.A(n_59749), .B(n_17408), .C(n_59733), .D(n_17416)
		, .Z(n_233358825));
	notech_ao4 i_10582120(.A(n_60045), .B(n_17392), .C(n_59765), .D(n_17400)
		, .Z(n_233458826));
	notech_ao4 i_10682122(.A(n_60077), .B(n_17376), .C(n_60061), .D(n_17384)
		, .Z(n_233658828));
	notech_ao4 i_10782123(.A(n_59996), .B(n_17328), .C(n_60093), .D(n_17360)
		, .Z(n_233758829));
	notech_and4 i_11382125(.A(n_233758829), .B(n_233658828), .C(n_233458826)
		, .D(n_233358825), .Z(n_233958831));
	notech_ao4 i_13282127(.A(n_60029), .B(n_17360), .C(n_60013), .D(n_17376)
		, .Z(n_234158833));
	notech_ao4 i_13382129(.A(n_59966), .B(n_17344), .C(n_59685), .D(n_17479)
		, .Z(n_234358835));
	notech_ao4 i_13482130(.A(n_59717), .B(n_17447), .C(n_59701), .D(n_17463)
		, .Z(n_234458836));
	notech_and4 i_14382132(.A(n_234458836), .B(n_234358835), .C(n_234158833)
		, .D(n_148057972), .Z(n_234658838));
	notech_ao4 i_13582133(.A(n_59749), .B(n_17416), .C(n_59733), .D(n_17431)
		, .Z(n_234758839));
	notech_ao4 i_13682134(.A(n_60045), .B(n_17400), .C(n_59765), .D(n_17408)
		, .Z(n_234858840));
	notech_ao4 i_13782136(.A(n_60077), .B(n_17384), .C(n_60061), .D(n_17392)
		, .Z(n_235058842));
	notech_ao4 i_13882137(.A(n_59996), .B(n_17336), .C(n_60093), .D(n_17368)
		, .Z(n_235158843));
	notech_and4 i_14482139(.A(n_235158843), .B(n_235058842), .C(n_234858840)
		, .D(n_234758839), .Z(n_235358845));
	notech_ao4 i_19482141(.A(n_60029), .B(n_17378), .C(n_60013), .D(n_17394)
		, .Z(n_235558847));
	notech_ao4 i_19582143(.A(n_59966), .B(n_17362), .C(n_59685), .D(n_17515)
		, .Z(n_235758849));
	notech_ao4 i_19682144(.A(n_59717), .B(n_17483), .C(n_59701), .D(n_17499)
		, .Z(n_235858850));
	notech_and4 i_20582146(.A(n_235858850), .B(n_235758849), .C(n_235558847)
		, .D(n_149657988), .Z(n_236058852));
	notech_ao4 i_19782147(.A(n_59749), .B(n_17451), .C(n_59733), .D(n_17467)
		, .Z(n_236158853));
	notech_ao4 i_19882148(.A(n_60045), .B(n_17418), .C(n_59765), .D(n_17435)
		, .Z(n_236258854));
	notech_ao4 i_19982150(.A(n_60077), .B(n_17402), .C(n_60061), .D(n_17410)
		, .Z(n_236458856));
	notech_ao4 i_20082151(.A(n_59994), .B(n_17354), .C(n_60093), .D(n_17386)
		, .Z(n_236558857));
	notech_and4 i_20682153(.A(n_236558857), .B(n_236458856), .C(n_236258854)
		, .D(n_236158853), .Z(n_236758859));
	notech_ao4 i_22582155(.A(n_60029), .B(n_17379), .C(n_60013), .D(n_17395)
		, .Z(n_236958861));
	notech_ao4 i_22682157(.A(n_59966), .B(n_17363), .C(n_59685), .D(n_17517)
		, .Z(n_237158863));
	notech_ao4 i_22782158(.A(n_59717), .B(n_17485), .C(n_59701), .D(n_17501)
		, .Z(n_237258864));
	notech_and4 i_23682160(.A(n_237258864), .B(n_237158863), .C(n_236958861)
		, .D(n_151258004), .Z(n_237458866));
	notech_ao4 i_22882161(.A(n_59749), .B(n_17453), .C(n_59733), .D(n_17469)
		, .Z(n_237558867));
	notech_ao4 i_22982162(.A(n_60045), .B(n_17421), .C(n_59765), .D(n_17437)
		, .Z(n_237658868));
	notech_ao4 i_23082164(.A(n_60077), .B(n_17403), .C(n_60061), .D(n_17411)
		, .Z(n_237858870));
	notech_ao4 i_23182165(.A(n_59996), .B(n_17355), .C(n_60093), .D(n_17387)
		, .Z(n_237958871));
	notech_and4 i_23782167(.A(n_237958871), .B(n_237858870), .C(n_237658868)
		, .D(n_237558867), .Z(n_238158873));
	notech_ao4 i_25682169(.A(n_60029), .B(n_17380), .C(n_60013), .D(n_17396)
		, .Z(n_238358875));
	notech_ao4 i_25735709(.A(n_59966), .B(n_17364), .C(n_59685), .D(n_17519)
		, .Z(n_238558877));
	notech_ao4 i_25882171(.A(n_59717), .B(n_17487), .C(n_59701), .D(n_17503)
		, .Z(n_238658878));
	notech_and4 i_26782173(.A(n_238658878), .B(n_238558877), .C(n_238358875)
		, .D(n_152858020), .Z(n_238858880));
	notech_ao4 i_25982174(.A(n_59749), .B(n_17455), .C(n_59733), .D(n_17471)
		, .Z(n_238958881));
	notech_ao4 i_26082175(.A(n_60045), .B(n_17423), .C(n_59765), .D(n_17439)
		, .Z(n_239058882));
	notech_ao4 i_26182177(.A(n_60077), .B(n_17404), .C(n_60061), .D(n_17412)
		, .Z(n_239258884));
	notech_ao4 i_26282178(.A(n_59994), .B(n_17356), .C(n_60093), .D(n_17388)
		, .Z(n_239358885));
	notech_and4 i_26882180(.A(n_239358885), .B(n_239258884), .C(n_239058882)
		, .D(n_238958881), .Z(n_239558887));
	notech_ao4 i_28782182(.A(n_60029), .B(n_17381), .C(n_60013), .D(n_17397)
		, .Z(n_239758889));
	notech_ao4 i_28882184(.A(n_59966), .B(n_17365), .C(n_59685), .D(n_17521)
		, .Z(n_239958891));
	notech_ao4 i_28982185(.A(n_59717), .B(n_17489), .C(n_59701), .D(n_17505)
		, .Z(n_240058892));
	notech_and4 i_29882187(.A(n_240058892), .B(n_239958891), .C(n_239758889)
		, .D(n_154458036), .Z(n_240258894));
	notech_ao4 i_29082188(.A(n_59749), .B(n_17457), .C(n_59733), .D(n_17473)
		, .Z(n_240358895));
	notech_ao4 i_29182189(.A(n_60045), .B(n_17425), .C(n_59765), .D(n_17441)
		, .Z(n_240458896));
	notech_ao4 i_29282191(.A(n_60077), .B(n_17405), .C(n_60061), .D(n_17413)
		, .Z(n_240658898));
	notech_ao4 i_29382192(.A(n_59994), .B(n_17357), .C(n_60093), .D(n_17389)
		, .Z(n_240758899));
	notech_and4 i_29982194(.A(n_240758899), .B(n_240658898), .C(n_240458896)
		, .D(n_240358895), .Z(n_240958901));
	notech_ao4 i_31882196(.A(n_60027), .B(n_17382), .C(n_60011), .D(n_17398)
		, .Z(n_241158903));
	notech_ao4 i_31982198(.A(n_59966), .B(n_17366), .C(n_59683), .D(n_17523)
		, .Z(n_241358905));
	notech_ao4 i_32082199(.A(n_59715), .B(n_17491), .C(n_59699), .D(n_17507)
		, .Z(n_241458906));
	notech_and4 i_32982201(.A(n_241458906), .B(n_241358905), .C(n_241158903)
		, .D(n_156058052), .Z(n_241658908));
	notech_ao4 i_32182202(.A(n_59747), .B(n_17459), .C(n_59731), .D(n_17475)
		, .Z(n_241758909));
	notech_ao4 i_32282203(.A(n_60043), .B(n_17427), .C(n_59763), .D(n_17443)
		, .Z(n_241858910));
	notech_ao4 i_32382205(.A(n_60075), .B(n_17406), .C(n_60059), .D(n_17414)
		, .Z(n_242058912));
	notech_ao4 i_32482206(.A(n_59994), .B(n_17358), .C(n_60091), .D(n_17390)
		, .Z(n_242158913));
	notech_and4 i_33082208(.A(n_242158913), .B(n_242058912), .C(n_241858910)
		, .D(n_241758909), .Z(n_242358915));
	notech_ao4 i_38082210(.A(n_60027), .B(n_17384), .C(n_60011), .D(n_17400)
		, .Z(n_242558917));
	notech_ao4 i_38182212(.A(n_59963), .B(n_17368), .C(n_59683), .D(n_17527)
		, .Z(n_242758919));
	notech_ao4 i_38282213(.A(n_59715), .B(n_17495), .C(n_59699), .D(n_17511)
		, .Z(n_242858920));
	notech_and4 i_39182215(.A(n_242858920), .B(n_242758919), .C(n_242558917)
		, .D(n_157658068), .Z(n_243058922));
	notech_ao4 i_38382216(.A(n_59747), .B(n_17463), .C(n_59731), .D(n_17479)
		, .Z(n_243158923));
	notech_ao4 i_38482217(.A(n_60043), .B(n_17431), .C(n_59763), .D(n_17447)
		, .Z(n_243258924));
	notech_ao4 i_38582219(.A(n_60075), .B(n_17408), .C(n_60059), .D(n_17416)
		, .Z(n_243458926));
	notech_ao4 i_38682220(.A(n_59996), .B(n_17360), .C(n_60091), .D(n_17392)
		, .Z(n_243558927));
	notech_and4 i_39282222(.A(n_243558927), .B(n_243458926), .C(n_243258924)
		, .D(n_243158923), .Z(n_243758929));
	notech_ao4 i_44282224(.A(n_60027), .B(n_17386), .C(n_60011), .D(n_17402)
		, .Z(n_243958931));
	notech_ao4 i_44382226(.A(n_59963), .B(n_17370), .C(n_59683), .D(n_17531)
		, .Z(n_244158933));
	notech_ao4 i_44482227(.A(n_59715), .B(n_17499), .C(n_59699), .D(n_17515)
		, .Z(n_244258934));
	notech_and4 i_45382229(.A(n_244258934), .B(n_244158933), .C(n_243958931)
		, .D(n_159258084), .Z(n_244458936));
	notech_ao4 i_44582230(.A(n_59747), .B(n_17467), .C(n_59731), .D(n_17483)
		, .Z(n_244558937));
	notech_ao4 i_44682231(.A(n_60043), .B(n_17435), .C(n_59763), .D(n_17451)
		, .Z(n_244658938));
	notech_ao4 i_44782233(.A(n_60075), .B(n_17410), .C(n_60059), .D(n_17418)
		, .Z(n_244858940));
	notech_ao4 i_44882234(.A(n_59996), .B(n_17362), .C(n_60091), .D(n_17394)
		, .Z(n_244958941));
	notech_and4 i_45482236(.A(n_244958941), .B(n_244858940), .C(n_244658938)
		, .D(n_244558937), .Z(n_245158943));
	notech_ao4 i_50482238(.A(n_60027), .B(n_17389), .C(n_60011), .D(n_17405)
		, .Z(n_245358945));
	notech_ao4 i_50582240(.A(n_59963), .B(n_17373), .C(n_59683), .D(n_17537)
		, .Z(n_245558947));
	notech_ao4 i_50682241(.A(n_59715), .B(n_17505), .C(n_59699), .D(n_17521)
		, .Z(n_245658948));
	notech_and4 i_51582243(.A(n_245658948), .B(n_245558947), .C(n_245358945)
		, .D(n_160858100), .Z(n_245858950));
	notech_ao4 i_50782244(.A(n_59747), .B(n_17473), .C(n_59731), .D(n_17489)
		, .Z(n_245958951));
	notech_ao4 i_50882245(.A(n_60043), .B(n_17441), .C(n_59763), .D(n_17457)
		, .Z(n_246058952));
	notech_ao4 i_50982247(.A(n_60075), .B(n_17413), .C(n_60059), .D(n_17425)
		, .Z(n_246258954));
	notech_ao4 i_51082248(.A(n_59996), .B(n_17365), .C(n_60091), .D(n_17397)
		, .Z(n_246358955));
	notech_and4 i_51682250(.A(n_246358955), .B(n_246258954), .C(n_246058952)
		, .D(n_245958951), .Z(n_246558957));
	notech_ao4 i_53582252(.A(n_60027), .B(n_17390), .C(n_60011), .D(n_17406)
		, .Z(n_246758959));
	notech_ao4 i_53682254(.A(n_59963), .B(n_17374), .C(n_59683), .D(n_17539)
		, .Z(n_246958961));
	notech_ao4 i_53782255(.A(n_59715), .B(n_17507), .C(n_59699), .D(n_17523)
		, .Z(n_247058962));
	notech_and4 i_54682257(.A(n_247058962), .B(n_246958961), .C(n_246758959)
		, .D(n_162458116), .Z(n_247258964));
	notech_ao4 i_53882258(.A(n_59747), .B(n_17475), .C(n_59731), .D(n_17491)
		, .Z(n_247358965));
	notech_ao4 i_53982259(.A(n_60043), .B(n_17443), .C(n_59763), .D(n_17459)
		, .Z(n_247458966));
	notech_ao4 i_54082261(.A(n_60075), .B(n_17414), .C(n_60059), .D(n_17427)
		, .Z(n_247658968));
	notech_ao4 i_54182262(.A(n_59996), .B(n_17366), .C(n_60091), .D(n_17398)
		, .Z(n_247758969));
	notech_and4 i_54782264(.A(n_247758969), .B(n_247658968), .C(n_247458966)
		, .D(n_247358965), .Z(n_247958971));
	notech_ao4 i_59782266(.A(n_60029), .B(n_17392), .C(n_60013), .D(n_17408)
		, .Z(n_248158973));
	notech_ao4 i_59882268(.A(n_59963), .B(n_17376), .C(n_59685), .D(n_17543)
		, .Z(n_248358975));
	notech_ao4 i_59982269(.A(n_59717), .B(n_17511), .C(n_59701), .D(n_17527)
		, .Z(n_248458976));
	notech_and4 i_60882271(.A(n_248458976), .B(n_248358975), .C(n_248158973)
		, .D(n_164058132), .Z(n_248658978));
	notech_ao4 i_60082272(.A(n_59749), .B(n_17479), .C(n_59733), .D(n_17495)
		, .Z(n_248758979));
	notech_ao4 i_60182273(.A(n_60045), .B(n_17447), .C(n_59765), .D(n_17463)
		, .Z(n_248858980));
	notech_ao4 i_60282275(.A(n_60077), .B(n_17416), .C(n_60061), .D(n_17431)
		, .Z(n_249058982));
	notech_ao4 i_60382276(.A(n_59996), .B(n_17368), .C(n_60093), .D(n_17400)
		, .Z(n_249158983));
	notech_and4 i_60982278(.A(n_249158983), .B(n_249058982), .C(n_248858980)
		, .D(n_248758979), .Z(n_249358985));
	notech_ao4 i_65982280(.A(n_60029), .B(n_17394), .C(n_60013), .D(n_17410)
		, .Z(n_249558987));
	notech_ao4 i_66082282(.A(n_59963), .B(n_17378), .C(n_59685), .D(n_17547)
		, .Z(n_249758989));
	notech_ao4 i_66182283(.A(n_59717), .B(n_17515), .C(n_59701), .D(n_17531)
		, .Z(n_249858990));
	notech_and4 i_67082285(.A(n_249858990), .B(n_249758989), .C(n_249558987)
		, .D(n_165658148), .Z(n_250058992));
	notech_ao4 i_66282286(.A(n_59749), .B(n_17483), .C(n_59733), .D(n_17499)
		, .Z(n_250158993));
	notech_ao4 i_66382287(.A(n_60045), .B(n_17451), .C(n_59765), .D(n_17467)
		, .Z(n_250258994));
	notech_ao4 i_66482289(.A(n_60077), .B(n_17418), .C(n_60061), .D(n_17435)
		, .Z(n_250458996));
	notech_ao4 i_66582290(.A(n_59996), .B(n_17370), .C(n_60093), .D(n_17402)
		, .Z(n_250558997));
	notech_and4 i_67182292(.A(n_250558997), .B(n_250458996), .C(n_250258994)
		, .D(n_250158993), .Z(n_250758999));
	notech_ao4 i_69082294(.A(n_60029), .B(n_17395), .C(n_60013), .D(n_17411)
		, .Z(n_250959001));
	notech_ao4 i_69182296(.A(n_59963), .B(n_17379), .C(n_59685), .D(n_17549)
		, .Z(n_251159003));
	notech_ao4 i_69282297(.A(n_59717), .B(n_17517), .C(n_59701), .D(n_17533)
		, .Z(n_251259004));
	notech_and4 i_70182299(.A(n_251259004), .B(n_251159003), .C(n_250959001)
		, .D(n_167258164), .Z(n_251459006));
	notech_ao4 i_69382300(.A(n_59749), .B(n_17485), .C(n_59733), .D(n_17501)
		, .Z(n_251559007));
	notech_ao4 i_69482301(.A(n_60045), .B(n_17453), .C(n_59765), .D(n_17469)
		, .Z(n_251659008));
	notech_ao4 i_69582303(.A(n_60077), .B(n_17421), .C(n_60061), .D(n_17437)
		, .Z(n_251859010));
	notech_ao4 i_69682304(.A(n_59982), .B(n_17371), .C(n_60093), .D(n_17403)
		, .Z(n_251959011));
	notech_and4 i_70282306(.A(n_251959011), .B(n_251859010), .C(n_251659008)
		, .D(n_251559007), .Z(n_252159013));
	notech_ao4 i_72182308(.A(n_60029), .B(n_17396), .C(n_60013), .D(n_17412)
		, .Z(n_252359015));
	notech_ao4 i_72282310(.A(n_59963), .B(n_17380), .C(n_59685), .D(n_17551)
		, .Z(n_252559017));
	notech_ao4 i_72382311(.A(n_59717), .B(n_17519), .C(n_59701), .D(n_17535)
		, .Z(n_252659018));
	notech_and4 i_73282313(.A(n_252659018), .B(n_252559017), .C(n_252359015)
		, .D(n_168858180), .Z(n_252859020));
	notech_ao4 i_72482314(.A(n_59749), .B(n_17487), .C(n_59733), .D(n_17503)
		, .Z(n_252959021));
	notech_ao4 i_72582315(.A(n_60045), .B(n_17455), .C(n_59765), .D(n_17471)
		, .Z(n_253059022));
	notech_ao4 i_72682317(.A(n_60077), .B(n_17423), .C(n_60061), .D(n_17439)
		, .Z(n_253259024));
	notech_ao4 i_72782318(.A(n_59982), .B(n_17372), .C(n_60093), .D(n_17404)
		, .Z(n_253359025));
	notech_and4 i_73382320(.A(n_253359025), .B(n_253259024), .C(n_253059022)
		, .D(n_252959021), .Z(n_253559027));
	notech_ao4 i_75282322(.A(n_60017), .B(n_17397), .C(n_60001), .D(n_17413)
		, .Z(n_253759029));
	notech_ao4 i_75382324(.A(n_59964), .B(n_17381), .C(n_59673), .D(n_17553)
		, .Z(n_253959031));
	notech_ao4 i_75482325(.A(n_59705), .B(n_17521), .C(n_59689), .D(n_17537)
		, .Z(n_254059032));
	notech_and4 i_76382327(.A(n_254059032), .B(n_253959031), .C(n_253759029)
		, .D(n_170458196), .Z(n_254259034));
	notech_ao4 i_75582328(.A(n_59737), .B(n_17489), .C(n_59721), .D(n_17505)
		, .Z(n_254359035));
	notech_ao4 i_75682329(.A(n_60033), .B(n_17457), .C(n_59753), .D(n_17473)
		, .Z(n_254459036));
	notech_ao4 i_75782331(.A(n_60065), .B(n_17425), .C(n_60049), .D(n_17441)
		, .Z(n_254659038));
	notech_ao4 i_75882332(.A(n_59982), .B(n_17373), .C(n_60081), .D(n_17405)
		, .Z(n_254759039));
	notech_and4 i_76482334(.A(n_254759039), .B(n_254659038), .C(n_254459036)
		, .D(n_254359035), .Z(n_254959041));
	notech_ao4 i_84582336(.A(n_60017), .B(n_17400), .C(n_60001), .D(n_17416)
		, .Z(n_255159043));
	notech_ao4 i_84682338(.A(n_59964), .B(n_17384), .C(n_59673), .D(n_17559)
		, .Z(n_255359045));
	notech_ao4 i_84782339(.A(n_59705), .B(n_17527), .C(n_59689), .D(n_17543)
		, .Z(n_255459046));
	notech_and4 i_85682341(.A(n_255459046), .B(n_255359045), .C(n_255159043)
		, .D(n_172058212), .Z(n_255659048));
	notech_ao4 i_84882342(.A(n_59737), .B(n_17495), .C(n_59721), .D(n_17511)
		, .Z(n_255759049));
	notech_ao4 i_84982343(.A(n_60033), .B(n_17463), .C(n_59753), .D(n_17479)
		, .Z(n_255859050));
	notech_ao4 i_85082345(.A(n_60065), .B(n_17431), .C(n_60049), .D(n_17447)
		, .Z(n_256059052));
	notech_ao4 i_85182346(.A(n_59982), .B(n_17376), .C(n_60081), .D(n_17408)
		, .Z(n_256159053));
	notech_and4 i_85782348(.A(n_256159053), .B(n_256059052), .C(n_255859050)
		, .D(n_255759049), .Z(n_256359055));
	notech_ao4 i_90782350(.A(n_60017), .B(n_17402), .C(n_60001), .D(n_17418)
		, .Z(n_256559057));
	notech_ao4 i_90882352(.A(n_59964), .B(n_17386), .C(n_59673), .D(n_17563)
		, .Z(n_256759059));
	notech_ao4 i_90982353(.A(n_59705), .B(n_17531), .C(n_59689), .D(n_17547)
		, .Z(n_256859060));
	notech_and4 i_91882355(.A(n_256859060), .B(n_256759059), .C(n_256559057)
		, .D(n_173658228), .Z(n_257059062));
	notech_ao4 i_91082356(.A(n_59737), .B(n_17499), .C(n_59721), .D(n_17515)
		, .Z(n_257159063));
	notech_ao4 i_91182357(.A(n_60033), .B(n_17467), .C(n_59753), .D(n_17483)
		, .Z(n_257259064));
	notech_ao4 i_91282359(.A(n_60065), .B(n_17435), .C(n_60049), .D(n_17451)
		, .Z(n_257459066));
	notech_ao4 i_91382360(.A(n_59982), .B(n_17378), .C(n_60081), .D(n_17410)
		, .Z(n_257559067));
	notech_and4 i_91982362(.A(n_257559067), .B(n_257459066), .C(n_257259064)
		, .D(n_257159063), .Z(n_257759069));
	notech_ao4 i_93882364(.A(n_60017), .B(n_17403), .C(n_60001), .D(n_17421)
		, .Z(n_257959071));
	notech_ao4 i_93982366(.A(n_59964), .B(n_17387), .C(n_59673), .D(n_17565)
		, .Z(n_258159073));
	notech_ao4 i_94082367(.A(n_59705), .B(n_17533), .C(n_59689), .D(n_17549)
		, .Z(n_258259074));
	notech_and4 i_94982369(.A(n_258259074), .B(n_258159073), .C(n_257959071)
		, .D(n_175258244), .Z(n_258459076));
	notech_ao4 i_94182370(.A(n_59737), .B(n_17501), .C(n_59721), .D(n_17517)
		, .Z(n_258559077));
	notech_ao4 i_94282371(.A(n_60033), .B(n_17469), .C(n_59753), .D(n_17485)
		, .Z(n_258659078));
	notech_ao4 i_94382373(.A(n_60065), .B(n_17437), .C(n_60049), .D(n_17453)
		, .Z(n_258859080));
	notech_ao4 i_94482374(.A(n_59982), .B(n_17379), .C(n_60081), .D(n_17411)
		, .Z(n_258959081));
	notech_and4 i_95082376(.A(n_258959081), .B(n_258859080), .C(n_258659078)
		, .D(n_258559077), .Z(n_259159083));
	notech_ao4 i_96982378(.A(n_60017), .B(n_17404), .C(n_60001), .D(n_17423)
		, .Z(n_259359085));
	notech_ao4 i_97082380(.A(n_59964), .B(n_17388), .C(n_59673), .D(n_17567)
		, .Z(n_259559087));
	notech_ao4 i_97182381(.A(n_59705), .B(n_17535), .C(n_59689), .D(n_17551)
		, .Z(n_259659088));
	notech_and4 i_98082383(.A(n_259659088), .B(n_259559087), .C(n_259359085)
		, .D(n_176858260), .Z(n_259859090));
	notech_ao4 i_97282384(.A(n_59737), .B(n_17503), .C(n_59721), .D(n_17519)
		, .Z(n_259959091));
	notech_ao4 i_97382385(.A(n_60033), .B(n_17471), .C(n_59753), .D(n_17487)
		, .Z(n_260059092));
	notech_ao4 i_97482387(.A(n_60065), .B(n_17439), .C(n_60049), .D(n_17455)
		, .Z(n_260259094));
	notech_ao4 i_97582388(.A(n_59988), .B(n_17380), .C(n_60081), .D(n_17412)
		, .Z(n_260359095));
	notech_and4 i_98182390(.A(n_260359095), .B(n_260259094), .C(n_260059092)
		, .D(n_259959091), .Z(n_260559097));
	notech_ao4 i_100082392(.A(n_60017), .B(n_17405), .C(n_60001), .D(n_17425
		), .Z(n_260759099));
	notech_ao4 i_100182394(.A(n_59964), .B(n_17389), .C(n_59673), .D(n_17569
		), .Z(n_260959101));
	notech_ao4 i_100282395(.A(n_59705), .B(n_17537), .C(n_59689), .D(n_17553
		), .Z(n_261059102));
	notech_and4 i_101182397(.A(n_261059102), .B(n_260959101), .C(n_260759099
		), .D(n_178458276), .Z(n_261259104));
	notech_ao4 i_100382398(.A(n_59737), .B(n_17505), .C(n_59721), .D(n_17521
		), .Z(n_261359105));
	notech_ao4 i_100482399(.A(n_60033), .B(n_17473), .C(n_59753), .D(n_17489
		), .Z(n_261459106));
	notech_ao4 i_100582401(.A(n_60065), .B(n_17441), .C(n_60049), .D(n_17457
		), .Z(n_261659108));
	notech_ao4 i_100682402(.A(n_59988), .B(n_17381), .C(n_60081), .D(n_17413
		), .Z(n_261759109));
	notech_and4 i_101282404(.A(n_261759109), .B(n_261659108), .C(n_261459106
		), .D(n_261359105), .Z(n_261959111));
	notech_ao4 i_103182406(.A(n_60027), .B(n_17406), .C(n_60011), .D(n_17427
		), .Z(n_262159113));
	notech_ao4 i_103282408(.A(n_59964), .B(n_17390), .C(n_59683), .D(n_17571
		), .Z(n_262359115));
	notech_ao4 i_103382409(.A(n_59715), .B(n_17539), .C(n_59699), .D(n_17555
		), .Z(n_262459116));
	notech_and4 i_104282411(.A(n_262459116), .B(n_262359115), .C(n_262159113
		), .D(n_180058292), .Z(n_262659118));
	notech_ao4 i_103482412(.A(n_59747), .B(n_17507), .C(n_59731), .D(n_17523
		), .Z(n_262759119));
	notech_ao4 i_103582413(.A(n_60043), .B(n_17475), .C(n_59763), .D(n_17491
		), .Z(n_262859120));
	notech_ao4 i_103682415(.A(n_60075), .B(n_17443), .C(n_60059), .D(n_17459
		), .Z(n_263059122));
	notech_ao4 i_103782416(.A(n_59988), .B(n_17382), .C(n_60091), .D(n_17414
		), .Z(n_263159123));
	notech_and4 i_104382418(.A(n_263159123), .B(n_263059122), .C(n_262859120
		), .D(n_262759119), .Z(n_263359125));
	notech_ao4 i_109382420(.A(n_60017), .B(n_17408), .C(n_60001), .D(n_17431
		), .Z(n_263559127));
	notech_ao4 i_109482422(.A(n_59964), .B(n_17392), .C(n_59673), .D(n_17575
		), .Z(n_263759129));
	notech_ao4 i_109582423(.A(n_59705), .B(n_17543), .C(n_59689), .D(n_17559
		), .Z(n_263859130));
	notech_and4 i_110482425(.A(n_263859130), .B(n_263759129), .C(n_263559127
		), .D(n_181658308), .Z(n_264059132));
	notech_ao4 i_109682426(.A(n_59737), .B(n_17511), .C(n_59721), .D(n_17527
		), .Z(n_264159133));
	notech_ao4 i_109782427(.A(n_60033), .B(n_17479), .C(n_59753), .D(n_17495
		), .Z(n_264259134));
	notech_ao4 i_109882429(.A(n_60065), .B(n_17447), .C(n_60049), .D(n_17463
		), .Z(n_264459136));
	notech_ao4 i_109982430(.A(n_59982), .B(n_17384), .C(n_60081), .D(n_17416
		), .Z(n_264559137));
	notech_and4 i_110582432(.A(n_264559137), .B(n_264459136), .C(n_264259134
		), .D(n_264159133), .Z(n_264759139));
	notech_ao4 i_115582434(.A(n_60017), .B(n_17410), .C(n_60001), .D(n_17435
		), .Z(n_264959141));
	notech_ao4 i_115682436(.A(n_59969), .B(n_17394), .C(n_59673), .D(n_17579
		), .Z(n_265159143));
	notech_ao4 i_115782437(.A(n_59705), .B(n_17547), .C(n_59689), .D(n_17563
		), .Z(n_265259144));
	notech_and4 i_116682439(.A(n_265259144), .B(n_265159143), .C(n_264959141
		), .D(n_183258324), .Z(n_265459146));
	notech_ao4 i_115882440(.A(n_59737), .B(n_17515), .C(n_59721), .D(n_17531
		), .Z(n_265559147));
	notech_ao4 i_115982441(.A(n_60033), .B(n_17483), .C(n_59753), .D(n_17499
		), .Z(n_265659148));
	notech_ao4 i_116082443(.A(n_60065), .B(n_17451), .C(n_60049), .D(n_17467
		), .Z(n_265859150));
	notech_ao4 i_116182444(.A(n_59988), .B(n_17386), .C(n_60081), .D(n_17418
		), .Z(n_265959151));
	notech_and4 i_116782446(.A(n_265959151), .B(n_265859150), .C(n_265659148
		), .D(n_265559147), .Z(n_266159153));
	notech_ao4 i_118682448(.A(n_60017), .B(n_17411), .C(n_60001), .D(n_17437
		), .Z(n_266359155));
	notech_ao4 i_118782450(.A(n_59969), .B(n_17395), .C(n_59673), .D(n_17581
		), .Z(n_266559157));
	notech_ao4 i_118882451(.A(n_59705), .B(n_17549), .C(n_59689), .D(n_17565
		), .Z(n_266659158));
	notech_and4 i_119782453(.A(n_266659158), .B(n_266559157), .C(n_266359155
		), .D(n_184858340), .Z(n_266859160));
	notech_ao4 i_118982454(.A(n_59737), .B(n_17517), .C(n_59721), .D(n_17533
		), .Z(n_266959161));
	notech_ao4 i_119082455(.A(n_60033), .B(n_17485), .C(n_59753), .D(n_17501
		), .Z(n_267059162));
	notech_ao4 i_119182457(.A(n_60065), .B(n_17453), .C(n_60049), .D(n_17469
		), .Z(n_267259164));
	notech_ao4 i_119282458(.A(n_59982), .B(n_17387), .C(n_60081), .D(n_17421
		), .Z(n_267359165));
	notech_and4 i_119882460(.A(n_267359165), .B(n_267259164), .C(n_267059162
		), .D(n_266959161), .Z(n_267559167));
	notech_ao4 i_121782462(.A(n_60017), .B(n_17412), .C(n_60001), .D(n_17439
		), .Z(n_267759169));
	notech_ao4 i_121882464(.A(n_59969), .B(n_17396), .C(n_59673), .D(n_17583
		), .Z(n_267959171));
	notech_ao4 i_121982465(.A(n_59705), .B(n_17551), .C(n_59689), .D(n_17567
		), .Z(n_268059172));
	notech_and4 i_122882467(.A(n_268059172), .B(n_267959171), .C(n_267759169
		), .D(n_186458356), .Z(n_268259174));
	notech_ao4 i_122082468(.A(n_59737), .B(n_17519), .C(n_59721), .D(n_17535
		), .Z(n_268359175));
	notech_ao4 i_122182469(.A(n_60033), .B(n_17487), .C(n_59753), .D(n_17503
		), .Z(n_268459176));
	notech_ao4 i_122282471(.A(n_60065), .B(n_17455), .C(n_60049), .D(n_17471
		), .Z(n_268659178));
	notech_ao4 i_122382472(.A(n_59982), .B(n_17388), .C(n_60081), .D(n_17423
		), .Z(n_268759179));
	notech_and4 i_122982474(.A(n_268759179), .B(n_268659178), .C(n_268459176
		), .D(n_268359175), .Z(n_268959181));
	notech_ao4 i_124882476(.A(n_60017), .B(n_17413), .C(n_60001), .D(n_17441
		), .Z(n_269159183));
	notech_ao4 i_124982478(.A(n_59969), .B(n_17397), .C(n_59673), .D(n_17585
		), .Z(n_269359185));
	notech_ao4 i_125082479(.A(n_59705), .B(n_17553), .C(n_59689), .D(n_17569
		), .Z(n_269459186));
	notech_and4 i_125982481(.A(n_269459186), .B(n_269359185), .C(n_269159183
		), .D(n_188058372), .Z(n_269659188));
	notech_ao4 i_125182482(.A(n_59737), .B(n_17521), .C(n_59721), .D(n_17537
		), .Z(n_269759189));
	notech_ao4 i_125282483(.A(n_60033), .B(n_17489), .C(n_59753), .D(n_17505
		), .Z(n_269859190));
	notech_ao4 i_125382485(.A(n_60065), .B(n_17457), .C(n_60049), .D(n_17473
		), .Z(n_270059192));
	notech_ao4 i_125482486(.A(n_59982), .B(n_17389), .C(n_60081), .D(n_17425
		), .Z(n_270159193));
	notech_and4 i_126082488(.A(n_270159193), .B(n_270059192), .C(n_269859190
		), .D(n_269759189), .Z(n_270359195));
	notech_ao4 i_127982490(.A(n_60017), .B(n_17414), .C(n_60001), .D(n_17443
		), .Z(n_270559197));
	notech_ao4 i_128082492(.A(n_59969), .B(n_17398), .C(n_59673), .D(n_17587
		), .Z(n_270759199));
	notech_ao4 i_128182493(.A(n_59705), .B(n_17555), .C(n_59689), .D(n_17571
		), .Z(n_270859200));
	notech_and4 i_129082495(.A(n_270859200), .B(n_270759199), .C(n_270559197
		), .D(n_189658388), .Z(n_271059202));
	notech_ao4 i_128282496(.A(n_59737), .B(n_17523), .C(n_59721), .D(n_17539
		), .Z(n_271159203));
	notech_ao4 i_128382497(.A(n_60033), .B(n_17491), .C(n_59753), .D(n_17507
		), .Z(n_271259204));
	notech_ao4 i_128482499(.A(n_60065), .B(n_17459), .C(n_60049), .D(n_17475
		), .Z(n_271459206));
	notech_ao4 i_128582500(.A(n_59982), .B(n_17390), .C(n_60081), .D(n_17427
		), .Z(n_271559207));
	notech_and4 i_129182502(.A(n_271559207), .B(n_271459206), .C(n_271259204
		), .D(n_271159203), .Z(n_271759209));
	notech_ao4 i_134182504(.A(n_60017), .B(n_17416), .C(n_60001), .D(n_17447
		), .Z(n_271959211));
	notech_ao4 i_134282506(.A(n_59969), .B(n_17400), .C(n_59673), .D(n_17591
		), .Z(n_272159213));
	notech_ao4 i_134382507(.A(n_59705), .B(n_17559), .C(n_59689), .D(n_17575
		), .Z(n_272259214));
	notech_and4 i_135282509(.A(n_272259214), .B(n_272159213), .C(n_271959211
		), .D(n_191258404), .Z(n_272459216));
	notech_ao4 i_134482510(.A(n_59737), .B(n_17527), .C(n_59721), .D(n_17543
		), .Z(n_272559217));
	notech_ao4 i_134582511(.A(n_60033), .B(n_17495), .C(n_59753), .D(n_17511
		), .Z(n_272659218));
	notech_ao4 i_134682513(.A(n_60065), .B(n_17463), .C(n_60049), .D(n_17479
		), .Z(n_272859220));
	notech_ao4 i_134782514(.A(n_59982), .B(n_17392), .C(n_60081), .D(n_17431
		), .Z(n_272959221));
	notech_and4 i_135382516(.A(n_272959221), .B(n_272859220), .C(n_272659218
		), .D(n_272559217), .Z(n_273159223));
	notech_ao4 i_140382518(.A(n_60017), .B(n_17418), .C(n_60001), .D(n_17451
		), .Z(n_273359225));
	notech_ao4 i_140482520(.A(n_59969), .B(n_17402), .C(n_59673), .D(n_17595
		), .Z(n_273559227));
	notech_ao4 i_140582521(.A(n_59705), .B(n_17563), .C(n_59689), .D(n_17579
		), .Z(n_273659228));
	notech_and4 i_141482523(.A(n_273659228), .B(n_273559227), .C(n_273359225
		), .D(n_192858420), .Z(n_273859230));
	notech_ao4 i_140682524(.A(n_59737), .B(n_17531), .C(n_59721), .D(n_17547
		), .Z(n_273959231));
	notech_ao4 i_140782525(.A(n_60033), .B(n_17499), .C(n_59753), .D(n_17515
		), .Z(n_274059232));
	notech_ao4 i_140882527(.A(n_60065), .B(n_17467), .C(n_60049), .D(n_17483
		), .Z(n_274259234));
	notech_ao4 i_140982528(.A(n_59982), .B(n_17394), .C(n_60081), .D(n_17435
		), .Z(n_274359235));
	notech_and4 i_141582530(.A(n_274359235), .B(n_274259234), .C(n_274059232
		), .D(n_273959231), .Z(n_274559237));
	notech_ao4 i_143482532(.A(n_60017), .B(n_17421), .C(n_60001), .D(n_17453
		), .Z(n_274759239));
	notech_ao4 i_143582534(.A(n_59969), .B(n_17403), .C(n_59673), .D(n_17597
		), .Z(n_274959241));
	notech_ao4 i_143682535(.A(n_59705), .B(n_17565), .C(n_59689), .D(n_17581
		), .Z(n_275059242));
	notech_and4 i_144582537(.A(n_275059242), .B(n_274959241), .C(n_274759239
		), .D(n_194458436), .Z(n_275259244));
	notech_ao4 i_143782538(.A(n_59737), .B(n_17533), .C(n_59721), .D(n_17549
		), .Z(n_275359245));
	notech_ao4 i_143882539(.A(n_60033), .B(n_17501), .C(n_59753), .D(n_17517
		), .Z(n_275459246));
	notech_ao4 i_143982541(.A(n_60065), .B(n_17469), .C(n_60049), .D(n_17485
		), .Z(n_275659248));
	notech_ao4 i_144082542(.A(n_59982), .B(n_17395), .C(n_60081), .D(n_17437
		), .Z(n_275759249));
	notech_and4 i_144682544(.A(n_275759249), .B(n_275659248), .C(n_275459246
		), .D(n_275359245), .Z(n_275959251));
	notech_ao4 i_146582546(.A(n_60017), .B(n_17423), .C(n_60001), .D(n_17455
		), .Z(n_276159253));
	notech_ao4 i_146682548(.A(n_59971), .B(n_17404), .C(n_59673), .D(n_17599
		), .Z(n_276359255));
	notech_ao4 i_146782549(.A(n_59705), .B(n_17567), .C(n_59689), .D(n_17583
		), .Z(n_276459256));
	notech_and4 i_147682551(.A(n_276459256), .B(n_276359255), .C(n_276159253
		), .D(n_196058452), .Z(n_276659258));
	notech_ao4 i_146882552(.A(n_59737), .B(n_17535), .C(n_59721), .D(n_17551
		), .Z(n_276759259));
	notech_ao4 i_146982553(.A(n_60033), .B(n_17503), .C(n_59753), .D(n_17519
		), .Z(n_276859260));
	notech_ao4 i_147082555(.A(n_60065), .B(n_17471), .C(n_60049), .D(n_17487
		), .Z(n_277059262));
	notech_ao4 i_147182556(.A(n_59982), .B(n_17396), .C(n_60081), .D(n_17439
		), .Z(n_277159263));
	notech_and4 i_147782558(.A(n_277159263), .B(n_277059262), .C(n_276859260
		), .D(n_276759259), .Z(n_277359265));
	notech_ao4 i_149682560(.A(n_60017), .B(n_17425), .C(n_60001), .D(n_17457
		), .Z(n_277559267));
	notech_ao4 i_149782562(.A(n_59971), .B(n_17405), .C(n_59673), .D(n_17601
		), .Z(n_277759269));
	notech_ao4 i_149882563(.A(n_59705), .B(n_17569), .C(n_59689), .D(n_17585
		), .Z(n_277859270));
	notech_and4 i_150782565(.A(n_277859270), .B(n_277759269), .C(n_277559267
		), .D(n_197658468), .Z(n_278059272));
	notech_ao4 i_149982566(.A(n_59737), .B(n_17537), .C(n_59721), .D(n_17553
		), .Z(n_278159273));
	notech_ao4 i_150082567(.A(n_60033), .B(n_17505), .C(n_59753), .D(n_17521
		), .Z(n_278259274));
	notech_ao4 i_150182569(.A(n_60065), .B(n_17473), .C(n_60049), .D(n_17489
		), .Z(n_278459276));
	notech_ao4 i_150282570(.A(n_59982), .B(n_17397), .C(n_60081), .D(n_17441
		), .Z(n_278559277));
	notech_and4 i_150882572(.A(n_278559277), .B(n_278459276), .C(n_278259274
		), .D(n_278159273), .Z(n_278759279));
	notech_ao4 i_152782574(.A(n_60017), .B(n_17427), .C(n_60001), .D(n_17459
		), .Z(n_278959281));
	notech_ao4 i_152882575(.A(n_59971), .B(n_17406), .C(n_59673), .D(n_17603
		), .Z(n_279159283));
	notech_ao4 i_152982576(.A(n_59705), .B(n_17571), .C(n_59689), .D(n_17587
		), .Z(n_279259284));
	notech_and4 i_1538(.A(n_279259284), .B(n_279159283), .C(n_278959281), .D
		(n_199258484), .Z(n_279459286));
	notech_ao4 i_153082577(.A(n_59737), .B(n_17539), .C(n_59721), .D(n_17555
		), .Z(n_279559287));
	notech_ao4 i_153182578(.A(n_60033), .B(n_17507), .C(n_59753), .D(n_17523
		), .Z(n_279659288));
	notech_ao4 i_153282579(.A(n_60065), .B(n_17475), .C(n_60049), .D(n_17491
		), .Z(n_279859290));
	notech_ao4 i_153382580(.A(n_59982), .B(n_17398), .C(n_60081), .D(n_17443
		), .Z(n_279959291));
	notech_and4 i_1539(.A(n_279959291), .B(n_279859290), .C(n_279659288), .D
		(n_279559287), .Z(n_280159293));
	notech_ao4 i_1589(.A(n_60027), .B(n_17431), .C(n_60011), .D(n_17463), .Z
		(n_280359295));
	notech_ao4 i_1590(.A(n_59971), .B(n_17408), .C(n_59683), .D(n_17607), .Z
		(n_280559297));
	notech_ao4 i_1591(.A(n_59715), .B(n_17575), .C(n_59699), .D(n_17591), .Z
		(n_280659298));
	notech_and4 i_1600(.A(n_280659298), .B(n_280559297), .C(n_280359295), .D
		(n_200858500), .Z(n_280859300));
	notech_ao4 i_1592(.A(n_59747), .B(n_17543), .C(n_59731), .D(n_17559), .Z
		(n_280959301));
	notech_ao4 i_1593(.A(n_60043), .B(n_17511), .C(n_59763), .D(n_17527), .Z
		(n_281059302));
	notech_ao4 i_1594(.A(n_60075), .B(n_17479), .C(n_60059), .D(n_17495), .Z
		(n_281259304));
	notech_ao4 i_1595(.A(n_59982), .B(n_17400), .C(n_60091), .D(n_17447), .Z
		(n_281359305));
	notech_and4 i_1601(.A(n_281359305), .B(n_281259304), .C(n_281059302), .D
		(n_280959301), .Z(n_281559307));
	notech_ao4 i_1651(.A(n_60023), .B(n_17435), .C(n_60007), .D(n_17467), .Z
		(n_281759309));
	notech_ao4 i_1652(.A(n_59971), .B(n_17410), .C(n_59679), .D(n_17611), .Z
		(n_281959311));
	notech_ao4 i_1653(.A(n_59711), .B(n_17579), .C(n_59695), .D(n_17595), .Z
		(n_282059312));
	notech_and4 i_1662(.A(n_282059312), .B(n_281959311), .C(n_281759309), .D
		(n_202458516), .Z(n_282259314));
	notech_ao4 i_1654(.A(n_59743), .B(n_17547), .C(n_59727), .D(n_17563), .Z
		(n_282359315));
	notech_ao4 i_1655(.A(n_60039), .B(n_17515), .C(n_59759), .D(n_17531), .Z
		(n_282459316));
	notech_ao4 i_1656(.A(n_60071), .B(n_17483), .C(n_60055), .D(n_17499), .Z
		(n_282659318));
	notech_ao4 i_1657(.A(n_59988), .B(n_17402), .C(n_60087), .D(n_17451), .Z
		(n_282759319));
	notech_and4 i_1663(.A(n_282759319), .B(n_282659318), .C(n_282459316), .D
		(n_282359315), .Z(n_282959321));
	notech_ao4 i_1682(.A(n_60023), .B(n_17437), .C(n_60007), .D(n_17469), .Z
		(n_283159323));
	notech_ao4 i_1683(.A(n_59969), .B(n_17411), .C(n_59679), .D(n_17613), .Z
		(n_283359325));
	notech_ao4 i_1684(.A(n_59711), .B(n_17581), .C(n_59695), .D(n_17597), .Z
		(n_283459326));
	notech_and4 i_1693(.A(n_283459326), .B(n_283359325), .C(n_283159323), .D
		(n_204058532), .Z(n_283659328));
	notech_ao4 i_1685(.A(n_59743), .B(n_17549), .C(n_59727), .D(n_17565), .Z
		(n_283759329));
	notech_ao4 i_1686(.A(n_60039), .B(n_17517), .C(n_59759), .D(n_17533), .Z
		(n_283859330));
	notech_ao4 i_1687(.A(n_60071), .B(n_17485), .C(n_60055), .D(n_17501), .Z
		(n_284059332));
	notech_ao4 i_1688(.A(n_59989), .B(n_17403), .C(n_60087), .D(n_17453), .Z
		(n_284159333));
	notech_and4 i_1694(.A(n_284159333), .B(n_284059332), .C(n_283859330), .D
		(n_283759329), .Z(n_284359335));
	notech_ao4 i_1713(.A(n_60023), .B(n_17439), .C(n_60007), .D(n_17471), .Z
		(n_284559337));
	notech_ao4 i_1714(.A(n_59971), .B(n_17412), .C(n_59679), .D(n_17615), .Z
		(n_284759339));
	notech_ao4 i_1715(.A(n_59711), .B(n_17583), .C(n_59695), .D(n_17599), .Z
		(n_284859340));
	notech_and4 i_1724(.A(n_284859340), .B(n_284759339), .C(n_284559337), .D
		(n_205658548), .Z(n_285059342));
	notech_ao4 i_1716(.A(n_59743), .B(n_17551), .C(n_59727), .D(n_17567), .Z
		(n_285159343));
	notech_ao4 i_1717(.A(n_60039), .B(n_17519), .C(n_59759), .D(n_17535), .Z
		(n_285259344));
	notech_ao4 i_1718(.A(n_60071), .B(n_17487), .C(n_60055), .D(n_17503), .Z
		(n_285459346));
	notech_ao4 i_1719(.A(n_59989), .B(n_17404), .C(n_60087), .D(n_17455), .Z
		(n_285559347));
	notech_and4 i_1725(.A(n_285559347), .B(n_285459346), .C(n_285259344), .D
		(n_285159343), .Z(n_285759349));
	notech_ao4 i_1744(.A(n_60023), .B(n_17441), .C(n_60007), .D(n_17473), .Z
		(n_285959351));
	notech_ao4 i_1745(.A(n_59971), .B(n_17413), .C(n_59679), .D(n_17617), .Z
		(n_286159353));
	notech_ao4 i_1746(.A(n_59711), .B(n_17585), .C(n_59695), .D(n_17601), .Z
		(n_286259354));
	notech_and4 i_1755(.A(n_286259354), .B(n_286159353), .C(n_285959351), .D
		(n_207258564), .Z(n_286459356));
	notech_ao4 i_1747(.A(n_59743), .B(n_17553), .C(n_59727), .D(n_17569), .Z
		(n_286559357));
	notech_ao4 i_1748(.A(n_60039), .B(n_17521), .C(n_59759), .D(n_17537), .Z
		(n_286659358));
	notech_ao4 i_1749(.A(n_60071), .B(n_17489), .C(n_60055), .D(n_17505), .Z
		(n_286859360));
	notech_ao4 i_1750(.A(n_59989), .B(n_17405), .C(n_60087), .D(n_17457), .Z
		(n_286959361));
	notech_and4 i_1756(.A(n_286959361), .B(n_286859360), .C(n_286659358), .D
		(n_286559357), .Z(n_287159363));
	notech_ao4 i_1775(.A(n_60023), .B(n_17443), .C(n_60007), .D(n_17475), .Z
		(n_287359365));
	notech_ao4 i_1776(.A(n_59966), .B(n_17414), .C(n_59679), .D(n_17619), .Z
		(n_287559367));
	notech_ao4 i_1777(.A(n_59711), .B(n_17587), .C(n_59695), .D(n_17603), .Z
		(n_287659368));
	notech_and4 i_1786(.A(n_287659368), .B(n_287559367), .C(n_287359365), .D
		(n_208858580), .Z(n_287859370));
	notech_ao4 i_1778(.A(n_59743), .B(n_17555), .C(n_59727), .D(n_17571), .Z
		(n_287959371));
	notech_ao4 i_1779(.A(n_60039), .B(n_17523), .C(n_59759), .D(n_17539), .Z
		(n_288059372));
	notech_ao4 i_1780(.A(n_60071), .B(n_17491), .C(n_60055), .D(n_17507), .Z
		(n_288259374));
	notech_ao4 i_1781(.A(n_59988), .B(n_17406), .C(n_60087), .D(n_17459), .Z
		(n_288359375));
	notech_and4 i_1787(.A(n_288359375), .B(n_288259374), .C(n_288059372), .D
		(n_287959371), .Z(n_288559377));
	notech_ao4 i_1837(.A(n_60023), .B(n_17447), .C(n_60007), .D(n_17479), .Z
		(n_288759379));
	notech_ao4 i_1838(.A(n_59966), .B(n_17416), .C(n_59679), .D(n_17623), .Z
		(n_288959381));
	notech_ao4 i_1839(.A(n_59711), .B(n_17591), .C(n_59695), .D(n_17607), .Z
		(n_289059382));
	notech_and4 i_1848(.A(n_289059382), .B(n_288959381), .C(n_288759379), .D
		(n_210458596), .Z(n_289259384));
	notech_ao4 i_1840(.A(n_59743), .B(n_17559), .C(n_59727), .D(n_17575), .Z
		(n_289359385));
	notech_ao4 i_1841(.A(n_60039), .B(n_17527), .C(n_59759), .D(n_17543), .Z
		(n_289459386));
	notech_ao4 i_1842(.A(n_60071), .B(n_17495), .C(n_60055), .D(n_17511), .Z
		(n_289659388));
	notech_ao4 i_1843(.A(n_59988), .B(n_17408), .C(n_60087), .D(n_17463), .Z
		(n_289759389));
	notech_and4 i_1849(.A(n_289759389), .B(n_289659388), .C(n_289459386), .D
		(n_289359385), .Z(n_289959391));
	notech_ao4 i_1899(.A(n_60023), .B(n_17451), .C(n_60007), .D(n_17483), .Z
		(n_290159393));
	notech_ao4 i_1900(.A(n_59966), .B(n_17418), .C(n_59679), .D(n_17627), .Z
		(n_290359395));
	notech_ao4 i_1901(.A(n_59711), .B(n_17595), .C(n_59695), .D(n_17611), .Z
		(n_290459396));
	notech_and4 i_1910(.A(n_290459396), .B(n_290359395), .C(n_290159393), .D
		(n_212058612), .Z(n_290659398));
	notech_ao4 i_1902(.A(n_59743), .B(n_17563), .C(n_59727), .D(n_17579), .Z
		(n_290759399));
	notech_ao4 i_1903(.A(n_60039), .B(n_17531), .C(n_59759), .D(n_17547), .Z
		(n_290859400));
	notech_ao4 i_1904(.A(n_60071), .B(n_17499), .C(n_60055), .D(n_17515), .Z
		(n_291059402));
	notech_ao4 i_1905(.A(n_59989), .B(n_17410), .C(n_60087), .D(n_17467), .Z
		(n_291159403));
	notech_and4 i_1911(.A(n_291159403), .B(n_291059402), .C(n_290859400), .D
		(n_290759399), .Z(n_291359405));
	notech_ao4 i_1930(.A(n_60023), .B(n_17453), .C(n_60007), .D(n_17485), .Z
		(n_291559407));
	notech_ao4 i_1931(.A(n_59966), .B(n_17421), .C(n_59679), .D(n_17629), .Z
		(n_291759409));
	notech_ao4 i_1932(.A(n_59711), .B(n_17597), .C(n_59695), .D(n_17613), .Z
		(n_291859410));
	notech_and4 i_1941(.A(n_291859410), .B(n_291759409), .C(n_291559407), .D
		(n_213658628), .Z(n_292059412));
	notech_ao4 i_1933(.A(n_59743), .B(n_17565), .C(n_59727), .D(n_17581), .Z
		(n_292159413));
	notech_ao4 i_1934(.A(n_60039), .B(n_17533), .C(n_59759), .D(n_17549), .Z
		(n_292259414));
	notech_ao4 i_1935(.A(n_60071), .B(n_17501), .C(n_60055), .D(n_17517), .Z
		(n_292459416));
	notech_ao4 i_1936(.A(n_59989), .B(n_17411), .C(n_60087), .D(n_17469), .Z
		(n_292559417));
	notech_and4 i_1942(.A(n_292559417), .B(n_292459416), .C(n_292259414), .D
		(n_292159413), .Z(n_292859419));
	notech_ao4 i_1961(.A(n_60023), .B(n_17455), .C(n_60007), .D(n_17487), .Z
		(n_293059421));
	notech_ao4 i_1962(.A(n_59966), .B(n_17423), .C(n_59679), .D(n_17631), .Z
		(n_293259423));
	notech_ao4 i_1963(.A(n_59711), .B(n_17599), .C(n_59695), .D(n_17615), .Z
		(n_293359424));
	notech_and4 i_1972(.A(n_293359424), .B(n_293259423), .C(n_293059421), .D
		(n_215258644), .Z(n_293559426));
	notech_ao4 i_1964(.A(n_59743), .B(n_17567), .C(n_59727), .D(n_17583), .Z
		(n_293759427));
	notech_ao4 i_1965(.A(n_60039), .B(n_17535), .C(n_59759), .D(n_17551), .Z
		(n_293859428));
	notech_ao4 i_1966(.A(n_60071), .B(n_17503), .C(n_60055), .D(n_17519), .Z
		(n_294159430));
	notech_ao4 i_1967(.A(n_59989), .B(n_17412), .C(n_60087), .D(n_17471), .Z
		(n_294259431));
	notech_and4 i_1973(.A(n_294259431), .B(n_294159430), .C(n_293859428), .D
		(n_293759427), .Z(n_294559433));
	notech_ao4 i_1992(.A(n_60029), .B(n_17457), .C(n_60013), .D(n_17489), .Z
		(n_294859435));
	notech_ao4 i_1993(.A(n_59966), .B(n_17425), .C(n_59685), .D(n_17633), .Z
		(n_295159437));
	notech_ao4 i_1994(.A(n_59717), .B(n_17601), .C(n_59701), .D(n_17617), .Z
		(n_295259438));
	notech_and4 i_2003(.A(n_295259438), .B(n_295159437), .C(n_294859435), .D
		(n_216858660), .Z(n_295559440));
	notech_ao4 i_1995(.A(n_59749), .B(n_17569), .C(n_59733), .D(n_17585), .Z
		(n_295659441));
	notech_ao4 i_1996(.A(n_60045), .B(n_17537), .C(n_59765), .D(n_17553), .Z
		(n_295759442));
	notech_ao4 i_1997(.A(n_60077), .B(n_17505), .C(n_60061), .D(n_17521), .Z
		(n_296059444));
	notech_ao4 i_1998(.A(n_59989), .B(n_17413), .C(n_60093), .D(n_17473), .Z
		(n_296159445));
	notech_and4 i_2004(.A(n_296159445), .B(n_296059444), .C(n_295759442), .D
		(n_295659441), .Z(n_296359447));
	notech_ao4 i_2023(.A(n_60027), .B(n_17459), .C(n_60011), .D(n_17491), .Z
		(n_296659449));
	notech_ao4 i_2024(.A(n_59966), .B(n_17427), .C(n_59683), .D(n_17635), .Z
		(n_296859451));
	notech_ao4 i_2025(.A(n_59715), .B(n_17603), .C(n_59699), .D(n_17619), .Z
		(n_296959452));
	notech_and4 i_2034(.A(n_296959452), .B(n_296859451), .C(n_296659449), .D
		(n_218458676), .Z(n_297159454));
	notech_ao4 i_2026(.A(n_59747), .B(n_17571), .C(n_59731), .D(n_17587), .Z
		(n_297259455));
	notech_ao4 i_2027(.A(n_60043), .B(n_17539), .C(n_59763), .D(n_17555), .Z
		(n_297359456));
	notech_ao4 i_2028(.A(n_60075), .B(n_17507), .C(n_60059), .D(n_17523), .Z
		(n_297559458));
	notech_ao4 i_2029(.A(n_59989), .B(n_17414), .C(n_60091), .D(n_17475), .Z
		(n_297659459));
	notech_and4 i_2035(.A(n_297659459), .B(n_297559458), .C(n_297359456), .D
		(n_297259455), .Z(n_297859461));
	notech_ao4 i_2085(.A(n_60027), .B(n_17463), .C(n_60011), .D(n_17495), .Z
		(n_298259463));
	notech_ao4 i_2086(.A(n_59966), .B(n_17431), .C(n_59683), .D(n_17639), .Z
		(n_298459465));
	notech_ao4 i_2087(.A(n_59715), .B(n_17607), .C(n_59699), .D(n_17623), .Z
		(n_298559466));
	notech_and4 i_2096(.A(n_298559466), .B(n_298459465), .C(n_298259463), .D
		(n_220058692), .Z(n_298759468));
	notech_ao4 i_2088(.A(n_59747), .B(n_17575), .C(n_59731), .D(n_17591), .Z
		(n_298859469));
	notech_ao4 i_2089(.A(n_60043), .B(n_17543), .C(n_59763), .D(n_17559), .Z
		(n_298959470));
	notech_ao4 i_2090(.A(n_60075), .B(n_17511), .C(n_60059), .D(n_17527), .Z
		(n_299159472));
	notech_ao4 i_2091(.A(n_59989), .B(n_17416), .C(n_60091), .D(n_17479), .Z
		(n_299259473));
	notech_and4 i_2097(.A(n_299259473), .B(n_299159472), .C(n_298959470), .D
		(n_298859469), .Z(n_299459475));
	notech_ao4 i_2147(.A(n_60027), .B(n_17467), .C(n_60011), .D(n_17499), .Z
		(n_299659477));
	notech_ao4 i_2148(.A(n_59969), .B(n_17435), .C(n_59683), .D(n_17643), .Z
		(n_299859479));
	notech_ao4 i_2149(.A(n_59715), .B(n_17611), .C(n_59699), .D(n_17627), .Z
		(n_299959480));
	notech_and4 i_2158(.A(n_299959480), .B(n_299859479), .C(n_299659477), .D
		(n_221658708), .Z(n_300159482));
	notech_ao4 i_2150(.A(n_59747), .B(n_17579), .C(n_59731), .D(n_17595), .Z
		(n_300259483));
	notech_ao4 i_2151(.A(n_60043), .B(n_17547), .C(n_59763), .D(n_17563), .Z
		(n_300359484));
	notech_ao4 i_2152(.A(n_60075), .B(n_17515), .C(n_60059), .D(n_17531), .Z
		(n_300559486));
	notech_ao4 i_2153(.A(n_59988), .B(n_17418), .C(n_60091), .D(n_17483), .Z
		(n_300659487));
	notech_and4 i_2159(.A(n_300659487), .B(n_300559486), .C(n_300359484), .D
		(n_300259483), .Z(n_300859489));
	notech_ao4 i_2178(.A(n_60027), .B(n_17469), .C(n_60011), .D(n_17501), .Z
		(n_301059491));
	notech_ao4 i_2179(.A(n_59969), .B(n_17437), .C(n_59683), .D(n_17645), .Z
		(n_301259493));
	notech_ao4 i_2180(.A(n_59715), .B(n_17613), .C(n_59699), .D(n_17629), .Z
		(n_301359494));
	notech_and4 i_2189(.A(n_301359494), .B(n_301259493), .C(n_301059491), .D
		(n_223258724), .Z(n_301559496));
	notech_ao4 i_2181(.A(n_59747), .B(n_17581), .C(n_59731), .D(n_17597), .Z
		(n_301659497));
	notech_ao4 i_2182(.A(n_60043), .B(n_17549), .C(n_59763), .D(n_17565), .Z
		(n_301759498));
	notech_ao4 i_2183(.A(n_60075), .B(n_17517), .C(n_60059), .D(n_17533), .Z
		(n_301959500));
	notech_ao4 i_2184(.A(n_59988), .B(n_17421), .C(n_60091), .D(n_17485), .Z
		(n_302059501));
	notech_and4 i_2190(.A(n_302059501), .B(n_301959500), .C(n_301759498), .D
		(n_301659497), .Z(n_302259503));
	notech_ao4 i_2209(.A(n_60029), .B(n_17471), .C(n_60013), .D(n_17503), .Z
		(n_302459505));
	notech_ao4 i_2210(.A(n_59969), .B(n_17439), .C(n_59685), .D(n_17647), .Z
		(n_302659507));
	notech_ao4 i_2211(.A(n_59717), .B(n_17615), .C(n_59701), .D(n_17631), .Z
		(n_302759508));
	notech_and4 i_2220(.A(n_302759508), .B(n_302659507), .C(n_302459505), .D
		(n_224858740), .Z(n_302959510));
	notech_ao4 i_2212(.A(n_59749), .B(n_17583), .C(n_59733), .D(n_17599), .Z
		(n_303059511));
	notech_ao4 i_2213(.A(n_60045), .B(n_17551), .C(n_59765), .D(n_17567), .Z
		(n_303159512));
	notech_ao4 i_2214(.A(n_60077), .B(n_17519), .C(n_60061), .D(n_17535), .Z
		(n_303359514));
	notech_ao4 i_2215(.A(n_59988), .B(n_17423), .C(n_60093), .D(n_17487), .Z
		(n_303459515));
	notech_and4 i_2221(.A(n_303459515), .B(n_303359514), .C(n_303159512), .D
		(n_303059511), .Z(n_303659517));
	notech_ao4 i_2240(.A(n_60029), .B(n_17473), .C(n_60013), .D(n_17505), .Z
		(n_303859519));
	notech_ao4 i_2241(.A(n_59969), .B(n_17441), .C(n_59685), .D(n_17649), .Z
		(n_304059521));
	notech_ao4 i_2242(.A(n_59717), .B(n_17617), .C(n_59701), .D(n_17633), .Z
		(n_304159522));
	notech_and4 i_2251(.A(n_304159522), .B(n_304059521), .C(n_303859519), .D
		(n_226458756), .Z(n_304359524));
	notech_ao4 i_2243(.A(n_59749), .B(n_17585), .C(n_59733), .D(n_17601), .Z
		(n_304459525));
	notech_ao4 i_2244(.A(n_60045), .B(n_17553), .C(n_59765), .D(n_17569), .Z
		(n_304559526));
	notech_ao4 i_2245(.A(n_60077), .B(n_17521), .C(n_60061), .D(n_17537), .Z
		(n_304759528));
	notech_ao4 i_2246(.A(n_59988), .B(n_17425), .C(n_60093), .D(n_17489), .Z
		(n_304859529));
	notech_and4 i_2252(.A(n_304859529), .B(n_304759528), .C(n_304559526), .D
		(n_304459525), .Z(n_305059531));
	notech_ao4 i_2271(.A(n_60029), .B(n_17475), .C(n_60013), .D(n_17507), .Z
		(n_305259533));
	notech_ao4 i_2272(.A(n_59969), .B(n_17443), .C(n_59685), .D(n_17651), .Z
		(n_305459535));
	notech_ao4 i_2273(.A(n_59717), .B(n_17619), .C(n_59701), .D(n_17635), .Z
		(n_305559536));
	notech_and4 i_2282(.A(n_305559536), .B(n_305459535), .C(n_305259533), .D
		(n_228058772), .Z(n_305759538));
	notech_ao4 i_2274(.A(n_59749), .B(n_17587), .C(n_59733), .D(n_17603), .Z
		(n_305859539));
	notech_ao4 i_2275(.A(n_60045), .B(n_17555), .C(n_59765), .D(n_17571), .Z
		(n_305959540));
	notech_ao4 i_2276(.A(n_60077), .B(n_17523), .C(n_60061), .D(n_17539), .Z
		(n_306159542));
	notech_ao4 i_2277(.A(n_59988), .B(n_17427), .C(n_60093), .D(n_17491), .Z
		(n_306259543));
	notech_and4 i_2283(.A(n_306259543), .B(n_306159542), .C(n_305959540), .D
		(n_305859539), .Z(n_306459545));
	notech_ao4 i_2333(.A(n_60029), .B(n_17479), .C(n_60013), .D(n_17511), .Z
		(n_306659547));
	notech_ao4 i_2334(.A(n_59969), .B(n_17447), .C(n_59685), .D(n_17655), .Z
		(n_306859549));
	notech_ao4 i_2335(.A(n_59717), .B(n_17623), .C(n_59701), .D(n_17639), .Z
		(n_306959550));
	notech_and4 i_2344(.A(n_306959550), .B(n_306859549), .C(n_306659547), .D
		(n_229658788), .Z(n_307159552));
	notech_ao4 i_2336(.A(n_59749), .B(n_17591), .C(n_59733), .D(n_17607), .Z
		(n_307259553));
	notech_ao4 i_2337(.A(n_60045), .B(n_17559), .C(n_59765), .D(n_17575), .Z
		(n_307359554));
	notech_ao4 i_2338(.A(n_60077), .B(n_17527), .C(n_60061), .D(n_17543), .Z
		(n_307559556));
	notech_ao4 i_2339(.A(n_59988), .B(n_17431), .C(n_60093), .D(n_17495), .Z
		(n_307659557));
	notech_and4 i_2345(.A(n_307659557), .B(n_307559556), .C(n_307359554), .D
		(n_307259553), .Z(n_307859559));
	notech_ao4 i_2395(.A(n_60029), .B(n_17483), .C(n_60013), .D(n_17515), .Z
		(n_308059561));
	notech_ao4 i_2396(.A(n_59969), .B(n_17451), .C(n_59685), .D(n_17659), .Z
		(n_308259563));
	notech_ao4 i_2397(.A(n_59717), .B(n_17627), .C(n_59701), .D(n_17643), .Z
		(n_308359564));
	notech_and4 i_2406(.A(n_308359564), .B(n_308259563), .C(n_308059561), .D
		(n_231258804), .Z(n_308559566));
	notech_ao4 i_2398(.A(n_59749), .B(n_17595), .C(n_59733), .D(n_17611), .Z
		(n_308659567));
	notech_ao4 i_2399(.A(n_60045), .B(n_17563), .C(n_59765), .D(n_17579), .Z
		(n_308759568));
	notech_ao4 i_2400(.A(n_60077), .B(n_17531), .C(n_60061), .D(n_17547), .Z
		(n_308959570));
	notech_ao4 i_2401(.A(n_59988), .B(n_17435), .C(n_60093), .D(n_17499), .Z
		(n_309059571));
	notech_and4 i_2407(.A(n_309059571), .B(n_308959570), .C(n_308759568), .D
		(n_308659567), .Z(n_309259573));
	notech_nand3 i_65510(.A(n_100357535), .B(n_8293), .C(n_7794), .Z(n_36936
		));
	notech_nand3 i_93933991(.A(n_59659), .B(n_59931), .C(queue[31]), .Z(n_1622
		));
	notech_and4 i_64623(.A(n_309559576), .B(n_7794), .C(n_100657538), .D(n_100757539
		), .Z(\nbus_12116[0] ));
	notech_nor2 i_6835700(.A(fault_wptr[0]), .B(fault_wptr[1]), .Z(n_7792)
		);
	notech_ao4 i_222675(.A(n_17301), .B(n_8293), .C(n_99957531), .D(n_14278717
		), .Z(n_34958));
	notech_nao3 i_7266(.A(pg_fault), .B(n_17298), .C(n_61438), .Z(n_8293));
	notech_nao3 i_2634897(.A(n_8293), .B(n_309659577), .C(n_61567), .Z(n_309459575
		));
	notech_or4 i_6534926(.A(n_61567), .B(n_17293), .C(n_17297), .D(n_61145),
		 .Z(n_7795));
	notech_or2 i_7134929(.A(n_101657548), .B(n_309459575), .Z(n_309559576)
		);
	notech_nand2 i_211934961(.A(n_7792), .B(fault_wptr_en), .Z(n_309659577)
		);
	notech_nor2 i_3734958(.A(n_14128702), .B(n_61388), .Z(n_309759578));
	notech_nand2 i_5051(.A(n_17862), .B(n_17861), .Z(n_312459605));
	notech_or4 i_3834923(.A(nbus_12105[5]), .B(nbus_12105[4]), .C(nbus_12105
		[6]), .D(n_14238713), .Z(n_14228712));
	notech_nand2 i_211634922(.A(code_ack), .B(n_62847), .Z(n_312559606));
	notech_nao3 i_7269(.A(n_17862), .B(n_17861), .C(nbus_12105[6]), .Z(n_14258715
		));
	notech_or2 i_92634004(.A(n_59988), .B(n_17330), .Z(n_1609));
	notech_and4 i_3124997(.A(n_2385), .B(n_2384), .C(n_2379), .D(n_2383), .Z
		(squeue_30101058));
	notech_nand3 i_90834022(.A(n_59659), .B(n_59931), .C(queue[30]), .Z(n_1606
		));
	notech_or2 i_89534035(.A(n_59988), .B(n_17329), .Z(n_1593));
	notech_and4 i_2924995(.A(n_2371), .B(n_2370), .C(n_2365), .D(n_2369), .Z
		(squeue_28101059));
	notech_nand3 i_87734053(.A(n_59659), .B(n_59931), .C(queue[28]), .Z(n_1590
		));
	notech_nand3 i_4235426(.A(code_ack), .B(n_62846), .C(n_8288), .Z(n_8359690
		));
	notech_ao3 i_22935244(.A(n_61390), .B(n_17861), .C(n_61567), .Z(n_26059867
		));
	notech_ao4 i_4435425(.A(n_61563), .B(n_61390), .C(n_51860125), .D(n_17861
		), .Z(n_26359870));
	notech_xor2 i_3935429(.A(addrshft[4]), .B(n_46960076), .Z(n_26759874));
	notech_and2 i_27835195(.A(purge_cnt[10]), .B(purge), .Z(n_29559902));
	notech_or4 i_28035193(.A(n_61145), .B(n_309459575), .C(n_17294), .D(n_7792
		), .Z(n_29759904));
	notech_or4 i_3535433(.A(useq_ptr[3]), .B(useq_ptr[2]), .C(useq_ptr[1]), 
		.D(useq_ptr[0]), .Z(n_29859905));
	notech_and2 i_5020(.A(addr_0[0]), .B(n_17991), .Z(n_29959906));
	notech_and2 i_5022(.A(addr_0[1]), .B(n_17991), .Z(n_30059907));
	notech_and2 i_5023(.A(addr_0[2]), .B(n_17991), .Z(n_30159908));
	notech_and2 i_5024(.A(addr_0[3]), .B(n_17991), .Z(n_30259909));
	notech_and2 i_5026(.A(n_34600), .B(n_47060077), .Z(n_30359910));
	notech_and2 i_5027(.A(n_34602), .B(n_47060077), .Z(n_30459911));
	notech_and2 i_5028(.A(n_34604), .B(n_47060077), .Z(n_30559912));
	notech_and2 i_5029(.A(n_34606), .B(n_47060077), .Z(n_30659913));
	notech_and2 i_5030(.A(n_34608), .B(n_47060077), .Z(n_30759914));
	notech_and2 i_5031(.A(n_34610), .B(n_47060077), .Z(n_30859915));
	notech_and2 i_5032(.A(n_34612), .B(n_47060077), .Z(n_30959916));
	notech_and2 i_5033(.A(n_34614), .B(n_47060077), .Z(n_31059917));
	notech_and2 i_5034(.A(n_34616), .B(n_47060077), .Z(n_31159918));
	notech_and2 i_5035(.A(n_34618), .B(n_47060077), .Z(n_31259919));
	notech_and2 i_5036(.A(n_34620), .B(n_47060077), .Z(n_31359920));
	notech_nor2 i_5037(.A(n_61567), .B(wptr[0]), .Z(n_31459921));
	notech_and2 i_5055(.A(n_63814), .B(n_8359690), .Z(codeWEN));
	notech_and2 i_334035461(.A(idata[0]), .B(n_63802), .Z(cacheD[0]));
	notech_and2 i_333935462(.A(idata[1]), .B(n_63802), .Z(cacheD[1]));
	notech_and2 i_333835463(.A(idata[2]), .B(n_63802), .Z(cacheD[2]));
	notech_and2 i_333735464(.A(idata[3]), .B(n_63802), .Z(cacheD[3]));
	notech_and2 i_333635465(.A(idata[4]), .B(n_63802), .Z(cacheD[4]));
	notech_and2 i_333535466(.A(idata[5]), .B(n_63802), .Z(cacheD[5]));
	notech_and2 i_333435467(.A(idata[6]), .B(n_63802), .Z(cacheD[6]));
	notech_and2 i_333335468(.A(idata[7]), .B(n_63802), .Z(cacheD[7]));
	notech_and2 i_333235469(.A(idata[8]), .B(n_63802), .Z(cacheD[8]));
	notech_and2 i_333135470(.A(idata[9]), .B(n_63802), .Z(cacheD[9]));
	notech_and2 i_333035471(.A(idata[10]), .B(n_63802), .Z(cacheD[10]));
	notech_and2 i_332935472(.A(idata[11]), .B(n_63802), .Z(cacheD[11]));
	notech_and2 i_332835473(.A(idata[12]), .B(n_63802), .Z(cacheD[12]));
	notech_and2 i_332735474(.A(idata[13]), .B(n_63802), .Z(cacheD[13]));
	notech_and2 i_332635475(.A(idata[14]), .B(n_63802), .Z(cacheD[14]));
	notech_and2 i_332535476(.A(idata[15]), .B(n_63802), .Z(cacheD[15]));
	notech_and2 i_332435477(.A(idata[16]), .B(n_63810), .Z(cacheD[16]));
	notech_and2 i_332335478(.A(idata[17]), .B(n_63810), .Z(cacheD[17]));
	notech_and2 i_332235479(.A(idata[18]), .B(n_63810), .Z(cacheD[18]));
	notech_and2 i_332135480(.A(idata[19]), .B(n_63810), .Z(cacheD[19]));
	notech_and2 i_332035481(.A(idata[20]), .B(n_63810), .Z(cacheD[20]));
	notech_and2 i_331935482(.A(idata[21]), .B(n_63810), .Z(cacheD[21]));
	notech_and2 i_331835483(.A(idata[22]), .B(n_63810), .Z(cacheD[22]));
	notech_and2 i_331735484(.A(idata[23]), .B(n_63810), .Z(cacheD[23]));
	notech_and2 i_331635485(.A(idata[24]), .B(n_63810), .Z(cacheD[24]));
	notech_and2 i_331535486(.A(idata[25]), .B(n_63810), .Z(cacheD[25]));
	notech_and2 i_331435487(.A(idata[26]), .B(n_63810), .Z(cacheD[26]));
	notech_and2 i_331335488(.A(idata[27]), .B(n_63810), .Z(cacheD[27]));
	notech_and2 i_331235489(.A(idata[28]), .B(n_63810), .Z(cacheD[28]));
	notech_and2 i_331135490(.A(idata[29]), .B(n_63810), .Z(cacheD[29]));
	notech_and2 i_331035491(.A(idata[30]), .B(n_63810), .Z(cacheD[30]));
	notech_and2 i_330935492(.A(idata[31]), .B(n_63810), .Z(cacheD[31]));
	notech_and2 i_330835493(.A(idata[32]), .B(n_63810), .Z(cacheD[32]));
	notech_and2 i_330735494(.A(idata[33]), .B(n_63810), .Z(cacheD[33]));
	notech_and2 i_330635495(.A(idata[34]), .B(n_63810), .Z(cacheD[34]));
	notech_and2 i_330535496(.A(idata[35]), .B(n_63814), .Z(cacheD[35]));
	notech_and2 i_330435497(.A(idata[36]), .B(n_63808), .Z(cacheD[36]));
	notech_and2 i_330335498(.A(idata[37]), .B(n_63808), .Z(cacheD[37]));
	notech_and2 i_330235499(.A(idata[38]), .B(n_63814), .Z(cacheD[38]));
	notech_and2 i_330135500(.A(idata[39]), .B(n_63814), .Z(cacheD[39]));
	notech_and2 i_330035501(.A(idata[40]), .B(n_63814), .Z(cacheD[40]));
	notech_and2 i_329935502(.A(idata[41]), .B(n_63814), .Z(cacheD[41]));
	notech_and2 i_329835503(.A(idata[42]), .B(n_63814), .Z(cacheD[42]));
	notech_and2 i_329735504(.A(idata[43]), .B(n_63814), .Z(cacheD[43]));
	notech_and2 i_329635505(.A(idata[44]), .B(n_63814), .Z(cacheD[44]));
	notech_and2 i_329535506(.A(idata[45]), .B(n_63814), .Z(cacheD[45]));
	notech_and2 i_329435507(.A(idata[46]), .B(n_63814), .Z(cacheD[46]));
	notech_and2 i_329335508(.A(idata[47]), .B(n_63814), .Z(cacheD[47]));
	notech_and2 i_329235509(.A(idata[48]), .B(n_63814), .Z(cacheD[48]));
	notech_and2 i_329135510(.A(idata[49]), .B(n_63814), .Z(cacheD[49]));
	notech_and2 i_329035511(.A(idata[50]), .B(n_63814), .Z(cacheD[50]));
	notech_and2 i_328935512(.A(idata[51]), .B(n_63814), .Z(cacheD[51]));
	notech_and2 i_328835513(.A(idata[52]), .B(n_63814), .Z(cacheD[52]));
	notech_and2 i_328735514(.A(idata[53]), .B(n_63814), .Z(cacheD[53]));
	notech_and2 i_328635515(.A(idata[54]), .B(n_63814), .Z(cacheD[54]));
	notech_and2 i_328535516(.A(idata[55]), .B(n_63808), .Z(cacheD[55]));
	notech_and2 i_328435517(.A(idata[56]), .B(n_63808), .Z(cacheD[56]));
	notech_and2 i_328335518(.A(idata[57]), .B(n_63808), .Z(cacheD[57]));
	notech_and2 i_328235519(.A(idata[58]), .B(n_63808), .Z(cacheD[58]));
	notech_and2 i_328135520(.A(idata[59]), .B(n_63808), .Z(cacheD[59]));
	notech_and2 i_328035521(.A(idata[60]), .B(n_63808), .Z(cacheD[60]));
	notech_and2 i_327935522(.A(idata[61]), .B(n_63808), .Z(cacheD[61]));
	notech_and2 i_327835523(.A(idata[62]), .B(n_63808), .Z(cacheD[62]));
	notech_and2 i_327735524(.A(idata[63]), .B(n_63808), .Z(cacheD[63]));
	notech_and2 i_327635525(.A(idata[64]), .B(n_63808), .Z(cacheD[64]));
	notech_and2 i_327535526(.A(idata[65]), .B(n_63808), .Z(cacheD[65]));
	notech_and2 i_327435527(.A(idata[66]), .B(n_63808), .Z(cacheD[66]));
	notech_and2 i_327335528(.A(idata[67]), .B(n_63808), .Z(cacheD[67]));
	notech_and2 i_327235529(.A(idata[68]), .B(n_63808), .Z(cacheD[68]));
	notech_and2 i_327135530(.A(idata[69]), .B(n_63808), .Z(cacheD[69]));
	notech_and2 i_327035531(.A(idata[70]), .B(n_63802), .Z(cacheD[70]));
	notech_and2 i_326935532(.A(idata[71]), .B(n_63802), .Z(cacheD[71]));
	notech_and2 i_326835533(.A(idata[72]), .B(n_63808), .Z(cacheD[72]));
	notech_and2 i_326735534(.A(idata[73]), .B(n_63812), .Z(cacheD[73]));
	notech_and2 i_326635535(.A(idata[74]), .B(n_63804), .Z(cacheD[74]));
	notech_and2 i_326535536(.A(idata[75]), .B(n_63804), .Z(cacheD[75]));
	notech_and2 i_326435537(.A(idata[76]), .B(n_63804), .Z(cacheD[76]));
	notech_and2 i_326335538(.A(idata[77]), .B(n_63804), .Z(cacheD[77]));
	notech_and2 i_326235539(.A(idata[78]), .B(n_63804), .Z(cacheD[78]));
	notech_and2 i_326135540(.A(idata[79]), .B(n_63804), .Z(cacheD[79]));
	notech_and2 i_326035541(.A(idata[80]), .B(n_63804), .Z(cacheD[80]));
	notech_and2 i_325935542(.A(idata[81]), .B(n_63804), .Z(cacheD[81]));
	notech_and2 i_325835543(.A(idata[82]), .B(n_63804), .Z(cacheD[82]));
	notech_and2 i_325735544(.A(idata[83]), .B(n_63804), .Z(cacheD[83]));
	notech_and2 i_325635545(.A(idata[84]), .B(n_63804), .Z(cacheD[84]));
	notech_and2 i_325535546(.A(idata[85]), .B(n_63804), .Z(cacheD[85]));
	notech_and2 i_325435547(.A(idata[86]), .B(n_63804), .Z(cacheD[86]));
	notech_and2 i_325335548(.A(idata[87]), .B(n_63804), .Z(cacheD[87]));
	notech_and2 i_325235549(.A(idata[88]), .B(n_63804), .Z(cacheD[88]));
	notech_and2 i_325135550(.A(idata[89]), .B(n_63804), .Z(cacheD[89]));
	notech_and2 i_325035551(.A(idata[90]), .B(n_63804), .Z(cacheD[90]));
	notech_and2 i_324935552(.A(idata[91]), .B(n_63812), .Z(cacheD[91]));
	notech_and2 i_324835553(.A(idata[92]), .B(n_63812), .Z(cacheD[92]));
	notech_and2 i_324735554(.A(idata[93]), .B(n_63812), .Z(cacheD[93]));
	notech_and2 i_324635555(.A(idata[94]), .B(n_63812), .Z(cacheD[94]));
	notech_and2 i_324535556(.A(idata[95]), .B(n_63812), .Z(cacheD[95]));
	notech_and2 i_324435557(.A(idata[96]), .B(n_63812), .Z(cacheD[96]));
	notech_and2 i_324335558(.A(idata[97]), .B(n_63812), .Z(cacheD[97]));
	notech_and2 i_324235559(.A(idata[98]), .B(n_63812), .Z(cacheD[98]));
	notech_and2 i_324135560(.A(idata[99]), .B(n_63812), .Z(cacheD[99]));
	notech_and2 i_324035561(.A(idata[100]), .B(n_63812), .Z(cacheD[100]));
	notech_and2 i_323935562(.A(idata[101]), .B(n_63812), .Z(cacheD[101]));
	notech_and2 i_323835563(.A(idata[102]), .B(n_63812), .Z(cacheD[102]));
	notech_and2 i_323735564(.A(idata[103]), .B(n_63812), .Z(cacheD[103]));
	notech_and2 i_323635565(.A(idata[104]), .B(n_63812), .Z(cacheD[104]));
	notech_and2 i_323535566(.A(idata[105]), .B(n_63812), .Z(cacheD[105]));
	notech_and2 i_323435567(.A(idata[106]), .B(n_63812), .Z(cacheD[106]));
	notech_and2 i_323335568(.A(idata[107]), .B(n_63812), .Z(cacheD[107]));
	notech_and2 i_323235569(.A(idata[108]), .B(n_63804), .Z(cacheD[108]));
	notech_and2 i_323135570(.A(idata[109]), .B(n_63812), .Z(cacheD[109]));
	notech_and2 i_323035571(.A(idata[110]), .B(n_63806), .Z(cacheD[110]));
	notech_and2 i_322935572(.A(idata[111]), .B(n_63806), .Z(cacheD[111]));
	notech_and2 i_322835573(.A(idata[112]), .B(n_63806), .Z(cacheD[112]));
	notech_and2 i_322735574(.A(idata[113]), .B(n_63806), .Z(cacheD[113]));
	notech_and2 i_322635575(.A(idata[114]), .B(n_63806), .Z(cacheD[114]));
	notech_and2 i_322535576(.A(idata[115]), .B(n_63806), .Z(cacheD[115]));
	notech_and2 i_322435577(.A(idata[116]), .B(n_63806), .Z(cacheD[116]));
	notech_and2 i_322335578(.A(idata[117]), .B(n_63806), .Z(cacheD[117]));
	notech_and2 i_322235579(.A(idata[118]), .B(n_63806), .Z(cacheD[118]));
	notech_and2 i_322135580(.A(idata[119]), .B(n_63806), .Z(cacheD[119]));
	notech_and2 i_322035581(.A(idata[120]), .B(n_63806), .Z(cacheD[120]));
	notech_and2 i_321935582(.A(idata[121]), .B(n_63806), .Z(cacheD[121]));
	notech_and2 i_321835583(.A(idata[122]), .B(n_63806), .Z(cacheD[122]));
	notech_and2 i_321735584(.A(idata[123]), .B(n_63806), .Z(cacheD[123]));
	notech_and2 i_321635585(.A(idata[124]), .B(n_63806), .Z(cacheD[124]));
	notech_and2 i_321535586(.A(idata[125]), .B(n_63806), .Z(cacheD[125]));
	notech_and2 i_321435587(.A(idata[126]), .B(n_63806), .Z(cacheD[126]));
	notech_and2 i_321335588(.A(idata[127]), .B(n_63806), .Z(cacheD[127]));
	notech_and2 i_321235589(.A(iaddr[14]), .B(n_63806), .Z(cacheD[128]));
	notech_and2 i_321135590(.A(iaddr[15]), .B(cacheD[148]), .Z(cacheD[129])
		);
	notech_and2 i_321035591(.A(iaddr[16]), .B(cacheD[148]), .Z(cacheD[130])
		);
	notech_and2 i_320935592(.A(iaddr[17]), .B(cacheD[148]), .Z(cacheD[131])
		);
	notech_and2 i_320835593(.A(iaddr[18]), .B(cacheD[148]), .Z(cacheD[132])
		);
	notech_and2 i_320735594(.A(iaddr[19]), .B(cacheD[148]), .Z(cacheD[133])
		);
	notech_and2 i_320635595(.A(iaddr[20]), .B(cacheD[148]), .Z(cacheD[134])
		);
	notech_and2 i_320535596(.A(iaddr[21]), .B(cacheD[148]), .Z(cacheD[135])
		);
	notech_and2 i_320435597(.A(iaddr[22]), .B(cacheD[148]), .Z(cacheD[136])
		);
	notech_and2 i_320335598(.A(iaddr[23]), .B(cacheD[148]), .Z(cacheD[137])
		);
	notech_and2 i_320235599(.A(iaddr[24]), .B(cacheD[148]), .Z(cacheD[138])
		);
	notech_and2 i_320135600(.A(iaddr[25]), .B(cacheD[148]), .Z(cacheD[139])
		);
	notech_and2 i_320035601(.A(iaddr[26]), .B(cacheD[148]), .Z(cacheD[140])
		);
	notech_and2 i_319935602(.A(iaddr[27]), .B(cacheD[148]), .Z(cacheD[141])
		);
	notech_and2 i_319835603(.A(iaddr[28]), .B(cacheD[148]), .Z(cacheD[142])
		);
	notech_and2 i_319735604(.A(iaddr[29]), .B(cacheD[148]), .Z(cacheD[143])
		);
	notech_and2 i_319635605(.A(iaddr[30]), .B(cacheD[148]), .Z(cacheD[144])
		);
	notech_and2 i_319535606(.A(iaddr[31]), .B(cacheD[148]), .Z(cacheD[145])
		);
	notech_nao3 i_28335190(.A(n_29859905), .B(n_61145), .C(n_309459575), .Z(n_46260069
		));
	notech_nand2 i_45335020(.A(n_17301), .B(n_17300), .Z(n_46860075));
	notech_or4 i_4035428(.A(addrshft[0]), .B(addrshft[1]), .C(addrshft[3]), 
		.D(addrshft[2]), .Z(n_46960076));
	notech_nor2 i_6235437(.A(n_61438), .B(purge_cnt[10]), .Z(n_47060077));
	notech_mux2 i_127170(.S(n_61567), .A(nbus_12105[0]), .B(pc_in[0]), .Z(n_35323
		));
	notech_mux2 i_222673(.S(n_52060127), .A(n_17296), .B(n_51960126), .Z(n_35229
		));
	notech_ao4 i_122674(.A(fault_wptr[0]), .B(n_14278717), .C(n_8293), .D(n_17300
		), .Z(n_34952));
	notech_mux2 i_2434925(.S(n_61567), .A(addr_0[23]), .B(pc_in[23]), .Z(n_37101
		));
	notech_ao4 i_23028617(.A(n_61372), .B(n_17834), .C(n_56561), .D(n_17899)
		, .Z(n_36755));
	notech_ao4 i_22828615(.A(n_61372), .B(n_17832), .C(n_56561), .D(n_17901)
		, .Z(n_36743));
	notech_ao4 i_22628613(.A(n_61372), .B(n_17830), .C(n_56561), .D(n_17903)
		, .Z(n_36731));
	notech_ao4 i_22428611(.A(n_61372), .B(n_17828), .C(n_56561), .D(n_17905)
		, .Z(n_36719));
	notech_ao4 i_22328610(.A(n_61316), .B(n_17827), .C(n_56561), .D(n_17906)
		, .Z(n_36713));
	notech_ao4 i_22128608(.A(n_61316), .B(n_17825), .C(n_56561), .D(n_17908)
		, .Z(n_36701));
	notech_ao4 i_22028607(.A(n_61316), .B(n_17824), .C(n_56561), .D(n_17909)
		, .Z(n_36695));
	notech_ao4 i_21928606(.A(n_61316), .B(n_17823), .C(n_56561), .D(n_17997)
		, .Z(n_36689));
	notech_ao4 i_21828605(.A(n_61316), .B(n_17822), .C(n_56561), .D(n_17910)
		, .Z(n_36683));
	notech_ao4 i_21728604(.A(n_61316), .B(n_17821), .C(n_56561), .D(n_17911)
		, .Z(n_36677));
	notech_ao4 i_21528602(.A(n_61316), .B(n_17819), .C(n_56561), .D(n_17912)
		, .Z(n_36665));
	notech_or4 i_178833142(.A(n_62847), .B(n_61421), .C(n_61392), .D(n_17996
		), .Z(n_50160108));
	notech_nand2 i_11628503(.A(n_52160128), .B(n_50160108), .Z(n_36071));
	notech_or4 i_189533035(.A(n_62847), .B(n_61424), .C(n_61392), .D(n_17997
		), .Z(n_50460111));
	notech_nand2 i_9128478(.A(n_52260129), .B(n_50460111), .Z(n_35921));
	notech_or4 i_219432742(.A(n_62847), .B(n_61424), .C(n_61392), .D(n_17995
		), .Z(n_50660113));
	notech_nand2 i_1928406(.A(n_52360130), .B(n_50660113), .Z(n_35489));
	notech_or4 i_221432722(.A(n_62847), .B(n_61424), .C(n_61392), .D(n_17994
		), .Z(n_50860115));
	notech_nand2 i_1428401(.A(n_52460131), .B(n_50860115), .Z(n_35459));
	notech_or4 i_221832718(.A(n_62847), .B(n_61424), .C(n_61390), .D(n_17993
		), .Z(n_51060117));
	notech_nand2 i_1328400(.A(n_52560132), .B(n_51060117), .Z(n_35453));
	notech_or4 i_225832678(.A(n_62847), .B(n_61421), .C(n_61390), .D(n_17992
		), .Z(n_51260119));
	notech_nand2 i_328390(.A(n_52660133), .B(n_51260119), .Z(n_35393));
	notech_or2 i_5095(.A(n_61567), .B(n_61146), .Z(n_51860125));
	notech_nor2 i_5096(.A(n_61567), .B(n_61392), .Z(n_51960126));
	notech_xor2 i_2234900(.A(wptr[0]), .B(n_61421), .Z(n_52060127));
	notech_ao4 i_179033140(.A(n_61146), .B(n_17651), .C(n_61316), .D(n_17848
		), .Z(n_52160128));
	notech_ao4 i_189833032(.A(n_61146), .B(n_17601), .C(n_61312), .D(n_17823
		), .Z(n_52260129));
	notech_ao4 i_219632740(.A(n_61312), .B(n_17751), .C(n_61146), .D(n_17457
		), .Z(n_52360130));
	notech_ao4 i_221632720(.A(n_61312), .B(n_17746), .C(n_61146), .D(n_17447
		), .Z(n_52460131));
	notech_ao4 i_222032716(.A(n_61312), .B(n_17745), .C(n_61146), .D(n_17445
		), .Z(n_52560132));
	notech_ao4 i_226032676(.A(n_61316), .B(n_17735), .C(n_61146), .D(n_17425
		), .Z(n_52660133));
	notech_nao3 i_64633(.A(n_7794), .B(n_8293), .C(n_17297), .Z(n_35236));
	notech_nand3 i_64683(.A(n_7794), .B(n_46260069), .C(n_7795), .Z(\nbus_12118[0] 
		));
	notech_nand3 i_64468(.A(n_8293), .B(n_7794), .C(n_29759904), .Z(\nbus_12115[0] 
		));
	notech_mux2 i_64477(.S(n_309659577), .A(n_8293), .B(n_130757805), .Z(n_34969
		));
	notech_or2 i_64638(.A(n_61438), .B(purge), .Z(\nbus_12117[0] ));
	notech_or2 i_65496(.A(n_61438), .B(n_29559902), .Z(n_36919));
	notech_ao4 i_64725(.A(n_61146), .B(n_309459575), .C(n_309559576), .D(n_52860135
		), .Z(\nbus_12119[128] ));
	notech_ao4 i_64724(.A(n_61146), .B(n_309459575), .C(n_309559576), .D(n_46860075
		), .Z(\nbus_12119[0] ));
	notech_mux2 i_135708(.S(purge), .A(iaddr[4]), .B(purge_cnt[0]), .Z(cacheA
		[0]));
	notech_mux2 i_211483(.S(purge), .A(iaddr[5]), .B(purge_cnt[1]), .Z(cacheA
		[1]));
	notech_mux2 i_335707(.S(purge), .A(iaddr[6]), .B(purge_cnt[2]), .Z(cacheA
		[2]));
	notech_mux2 i_435706(.S(purge), .A(iaddr[7]), .B(purge_cnt[3]), .Z(cacheA
		[3]));
	notech_mux2 i_511484(.S(purge), .A(iaddr[8]), .B(purge_cnt[4]), .Z(cacheA
		[4]));
	notech_mux2 i_635705(.S(purge), .A(iaddr[9]), .B(purge_cnt[5]), .Z(cacheA
		[5]));
	notech_mux2 i_735704(.S(purge), .A(iaddr[10]), .B(purge_cnt[6]), .Z(cacheA
		[6]));
	notech_mux2 i_835703(.S(purge), .A(iaddr[11]), .B(purge_cnt[7]), .Z(cacheA
		[7]));
	notech_mux2 i_935702(.S(purge), .A(iaddr[12]), .B(purge_cnt[8]), .Z(cacheA
		[8]));
	notech_mux2 i_1035701(.S(purge), .A(iaddr[13]), .B(purge_cnt[9]), .Z(cacheA
		[9]));
	notech_mux2 i_127158(.S(addrshft[0]), .A(n_3400), .B(n_113256518), .Z(valid_len_0101031
		));
	notech_ao4 i_527162(.A(addrshft[4]), .B(n_3400), .C(n_26759874), .D(n_113256518
		), .Z(valid_len_4101030));
	notech_ao4 i_627175(.A(n_312459605), .B(n_51860125), .C(n_26359870), .D(n_17862
		), .Z(n_35353));
	notech_mux2 i_427173(.S(n_61567), .A(nbus_12105[3]), .B(pc_in[3]), .Z(n_35341
		));
	notech_mux2 i_327172(.S(n_61567), .A(nbus_12105[2]), .B(pc_in[2]), .Z(n_35335
		));
	notech_mux2 i_227171(.S(n_61567), .A(nbus_12105[1]), .B(pc_in[1]), .Z(n_35329
		));
	notech_mux2 i_3235459(.S(n_61567), .A(addr_0[31]), .B(pc_in[31]), .Z(n_37149
		));
	notech_mux2 i_3135458(.S(n_61567), .A(addr_0[30]), .B(pc_in[30]), .Z(n_37143
		));
	notech_mux2 i_3035457(.S(n_61567), .A(addr_0[29]), .B(pc_in[29]), .Z(n_37137
		));
	notech_mux2 i_2935456(.S(n_61567), .A(addr_0[28]), .B(pc_in[28]), .Z(n_37131
		));
	notech_mux2 i_2835455(.S(n_61567), .A(addr_0[27]), .B(pc_in[27]), .Z(n_37125
		));
	notech_mux2 i_2735454(.S(n_61567), .A(addr_0[26]), .B(pc_in[26]), .Z(n_37119
		));
	notech_mux2 i_2635453(.S(n_61563), .A(addr_0[25]), .B(pc_in[25]), .Z(n_37113
		));
	notech_mux2 i_2535452(.S(n_61563), .A(addr_0[24]), .B(pc_in[24]), .Z(n_37107
		));
	notech_mux2 i_2335451(.S(n_61563), .A(addr_0[22]), .B(pc_in[22]), .Z(n_37095
		));
	notech_mux2 i_2235450(.S(n_61563), .A(addr_0[21]), .B(pc_in[21]), .Z(n_37089
		));
	notech_mux2 i_2135449(.S(n_61563), .A(addr_0[20]), .B(pc_in[20]), .Z(n_37083
		));
	notech_mux2 i_2035448(.S(n_61563), .A(addr_0[19]), .B(pc_in[19]), .Z(n_37077
		));
	notech_mux2 i_1935447(.S(n_61559), .A(addr_0[18]), .B(pc_in[18]), .Z(n_37071
		));
	notech_mux2 i_1835446(.S(n_61559), .A(addr_0[17]), .B(pc_in[17]), .Z(n_37065
		));
	notech_mux2 i_1735445(.S(n_61559), .A(addr_0[16]), .B(pc_in[16]), .Z(n_37059
		));
	notech_mux2 i_1635444(.S(n_61563), .A(addr_0[15]), .B(pc_in[15]), .Z(n_37053
		));
	notech_mux2 i_1535443(.S(n_61559), .A(addr_0[14]), .B(pc_in[14]), .Z(n_37047
		));
	notech_mux2 i_1435442(.S(n_61563), .A(addr_0[13]), .B(pc_in[13]), .Z(n_37041
		));
	notech_mux2 i_1335441(.S(n_61563), .A(addr_0[12]), .B(pc_in[12]), .Z(n_37035
		));
	notech_mux2 i_1235440(.S(n_61563), .A(addr_0[11]), .B(pc_in[11]), .Z(n_37029
		));
	notech_mux2 i_1135439(.S(n_61563), .A(addr_0[10]), .B(pc_in[10]), .Z(n_37023
		));
	notech_mux2 i_1022056(.S(n_61563), .A(addr_0[9]), .B(pc_in[9]), .Z(n_37017
		));
	notech_mux2 i_922055(.S(n_61563), .A(addr_0[8]), .B(pc_in[8]), .Z(n_37011
		));
	notech_mux2 i_822054(.S(n_61563), .A(addr_0[7]), .B(pc_in[7]), .Z(n_37005
		));
	notech_mux2 i_722053(.S(n_61563), .A(addr_0[6]), .B(pc_in[6]), .Z(n_36999
		));
	notech_mux2 i_622052(.S(n_61563), .A(addr_0[5]), .B(pc_in[5]), .Z(n_36993
		));
	notech_mux2 i_522051(.S(n_61563), .A(addr_0[4]), .B(pc_in[4]), .Z(n_36987
		));
	notech_ao4 i_25628643(.A(n_56561), .B(n_17874), .C(n_61316), .D(n_17860)
		, .Z(n_36911));
	notech_ao4 i_25528642(.A(n_56561), .B(n_17875), .C(n_61312), .D(n_17859)
		, .Z(n_36905));
	notech_ao4 i_25428641(.A(n_56561), .B(n_17876), .C(n_61316), .D(n_17858)
		, .Z(n_36899));
	notech_ao4 i_25328640(.A(n_56561), .B(n_17877), .C(n_61321), .D(n_17857)
		, .Z(n_36893));
	notech_ao4 i_25228639(.A(n_56559), .B(n_17878), .C(n_61321), .D(n_17856)
		, .Z(n_36887));
	notech_ao4 i_25128638(.A(n_56559), .B(n_17879), .C(n_61321), .D(n_17855)
		, .Z(n_36881));
	notech_ao4 i_25028637(.A(n_56559), .B(n_17880), .C(n_61321), .D(n_17854)
		, .Z(n_36875));
	notech_ao4 i_24928636(.A(n_56559), .B(n_17881), .C(n_61321), .D(n_17853)
		, .Z(n_36869));
	notech_ao4 i_24828635(.A(n_56559), .B(n_17882), .C(n_61321), .D(n_17852)
		, .Z(n_36863));
	notech_ao4 i_24728634(.A(n_56559), .B(n_17883), .C(n_61321), .D(n_17851)
		, .Z(n_36857));
	notech_ao4 i_24628633(.A(n_56559), .B(n_17884), .C(n_61321), .D(n_17850)
		, .Z(n_36851));
	notech_ao4 i_24528632(.A(n_56559), .B(n_17885), .C(n_61321), .D(n_17849)
		, .Z(n_36845));
	notech_ao4 i_24428631(.A(n_61321), .B(n_17848), .C(n_56559), .D(n_17996)
		, .Z(n_36839));
	notech_ao4 i_24328630(.A(n_56559), .B(n_17886), .C(n_61316), .D(n_17847)
		, .Z(n_36833));
	notech_ao4 i_24228629(.A(n_56559), .B(n_17887), .C(n_61316), .D(n_17846)
		, .Z(n_36827));
	notech_ao4 i_24128628(.A(n_56559), .B(n_17888), .C(n_61321), .D(n_17845)
		, .Z(n_36821));
	notech_ao4 i_24028627(.A(n_56559), .B(n_17889), .C(n_61321), .D(n_17844)
		, .Z(n_36815));
	notech_ao4 i_23928626(.A(n_56559), .B(n_17890), .C(n_61321), .D(n_17843)
		, .Z(n_36809));
	notech_ao4 i_23828625(.A(n_56559), .B(n_17891), .C(n_61321), .D(n_17842)
		, .Z(n_36803));
	notech_ao4 i_23728624(.A(n_56559), .B(n_17892), .C(n_61303), .D(n_17841)
		, .Z(n_36797));
	notech_ao4 i_23628623(.A(n_56566), .B(n_17893), .C(n_61303), .D(n_17840)
		, .Z(n_36791));
	notech_ao4 i_23528622(.A(n_56566), .B(n_17894), .C(n_61303), .D(n_17839)
		, .Z(n_36785));
	notech_ao4 i_23428621(.A(n_56566), .B(n_17895), .C(n_61303), .D(n_17838)
		, .Z(n_36779));
	notech_ao4 i_23328620(.A(n_56566), .B(n_17896), .C(n_61307), .D(n_17837)
		, .Z(n_36773));
	notech_ao4 i_23228619(.A(n_56566), .B(n_17897), .C(n_61307), .D(n_17836)
		, .Z(n_36767));
	notech_ao4 i_23128618(.A(n_61303), .B(n_17835), .C(n_56566), .D(n_17898)
		, .Z(n_36761));
	notech_ao4 i_22928616(.A(n_61307), .B(n_17833), .C(n_56566), .D(n_17900)
		, .Z(n_36749));
	notech_ao4 i_22728614(.A(n_61303), .B(n_17831), .C(n_56566), .D(n_17902)
		, .Z(n_36737));
	notech_ao4 i_22528612(.A(n_61303), .B(n_17829), .C(n_56566), .D(n_17904)
		, .Z(n_36725));
	notech_ao4 i_22228609(.A(n_61303), .B(n_17826), .C(n_56566), .D(n_17907)
		, .Z(n_36707));
	notech_ao4 i_21428601(.A(n_61303), .B(n_17818), .C(n_56566), .D(n_17913)
		, .Z(n_36659));
	notech_ao4 i_21328600(.A(n_61303), .B(n_17817), .C(n_56566), .D(n_17914)
		, .Z(n_36653));
	notech_ao4 i_21228599(.A(n_61303), .B(n_17816), .C(n_56566), .D(n_17915)
		, .Z(n_36647));
	notech_ao4 i_21128598(.A(n_61303), .B(n_17815), .C(n_56566), .D(n_17916)
		, .Z(n_36641));
	notech_ao4 i_21028597(.A(n_61303), .B(n_17814), .C(n_56566), .D(n_17917)
		, .Z(n_36635));
	notech_ao4 i_20928596(.A(n_61312), .B(n_17813), .C(n_56566), .D(n_17918)
		, .Z(n_36629));
	notech_ao4 i_20828595(.A(n_61312), .B(n_17812), .C(n_56564), .D(n_17919)
		, .Z(n_36623));
	notech_ao4 i_20728594(.A(n_61307), .B(n_17811), .C(n_56564), .D(n_17920)
		, .Z(n_36617));
	notech_ao4 i_20628593(.A(n_61312), .B(n_17810), .C(n_56564), .D(n_17921)
		, .Z(n_36611));
	notech_ao4 i_20528592(.A(n_61312), .B(n_17809), .C(n_56564), .D(n_17922)
		, .Z(n_36605));
	notech_ao4 i_20428591(.A(n_61312), .B(n_17808), .C(n_56564), .D(n_17923)
		, .Z(n_36599));
	notech_ao4 i_20328590(.A(n_61312), .B(n_17807), .C(n_56564), .D(n_17924)
		, .Z(n_36593));
	notech_ao4 i_20228589(.A(n_61312), .B(n_17806), .C(n_56564), .D(n_17925)
		, .Z(n_36587));
	notech_ao4 i_20128588(.A(n_61307), .B(n_17805), .C(n_56564), .D(n_17926)
		, .Z(n_36581));
	notech_ao4 i_20028587(.A(n_61307), .B(n_17804), .C(n_56564), .D(n_17927)
		, .Z(n_36575));
	notech_ao4 i_19928586(.A(n_61307), .B(n_17803), .C(n_56564), .D(n_17928)
		, .Z(n_36569));
	notech_ao4 i_19828585(.A(n_61307), .B(n_17802), .C(n_56564), .D(n_17929)
		, .Z(n_36563));
	notech_ao4 i_19728584(.A(n_61307), .B(n_17801), .C(n_56564), .D(n_17930)
		, .Z(n_36557));
	notech_ao4 i_19628583(.A(n_61307), .B(n_17800), .C(n_56564), .D(n_17931)
		, .Z(n_36551));
	notech_ao4 i_19528582(.A(n_61307), .B(n_17799), .C(n_56564), .D(n_17932)
		, .Z(n_36545));
	notech_ao4 i_19428581(.A(n_61307), .B(n_17798), .C(n_56564), .D(n_17933)
		, .Z(n_36539));
	notech_ao4 i_19328580(.A(n_61321), .B(n_17797), .C(n_56564), .D(n_17934)
		, .Z(n_36533));
	notech_ao4 i_19228579(.A(n_61335), .B(n_17796), .C(n_56551), .D(n_17935)
		, .Z(n_36527));
	notech_ao4 i_19128578(.A(n_61340), .B(n_17795), .C(n_56551), .D(n_17936)
		, .Z(n_36521));
	notech_ao4 i_19028577(.A(n_61335), .B(n_17794), .C(n_56551), .D(n_17937)
		, .Z(n_36515));
	notech_ao4 i_18928576(.A(n_61335), .B(n_17793), .C(n_56551), .D(n_17938)
		, .Z(n_36509));
	notech_ao4 i_18828575(.A(n_61340), .B(n_17792), .C(n_56551), .D(n_17939)
		, .Z(n_36503));
	notech_ao4 i_18728574(.A(n_61340), .B(n_17791), .C(n_56551), .D(n_17940)
		, .Z(n_36497));
	notech_ao4 i_18628573(.A(n_61340), .B(n_17790), .C(n_56551), .D(n_17941)
		, .Z(n_36491));
	notech_ao4 i_18528572(.A(n_61340), .B(n_17789), .C(n_56551), .D(n_17942)
		, .Z(n_36485));
	notech_ao4 i_18428571(.A(n_61335), .B(n_17788), .C(n_56551), .D(n_17943)
		, .Z(n_36479));
	notech_ao4 i_18328570(.A(n_56551), .B(n_17944), .C(n_61335), .D(n_17787)
		, .Z(n_36473));
	notech_ao4 i_18228569(.A(n_61335), .B(n_17786), .C(n_56551), .D(n_17945)
		, .Z(n_36467));
	notech_ao4 i_18128568(.A(n_61335), .B(n_17785), .C(n_56551), .D(n_17946)
		, .Z(n_36461));
	notech_ao4 i_18028567(.A(n_61335), .B(n_17784), .C(n_56551), .D(n_17947)
		, .Z(n_36455));
	notech_ao4 i_17928566(.A(n_61335), .B(n_17783), .C(n_56551), .D(n_17948)
		, .Z(n_36449));
	notech_ao4 i_17828565(.A(n_61335), .B(n_17782), .C(n_56551), .D(n_17949)
		, .Z(n_36443));
	notech_ao4 i_17728564(.A(n_61335), .B(n_17781), .C(n_56551), .D(n_17950)
		, .Z(n_36437));
	notech_ao4 i_17628563(.A(n_61344), .B(n_17780), .C(n_56549), .D(n_17951)
		, .Z(n_36431));
	notech_ao4 i_17528562(.A(n_61344), .B(n_17779), .C(n_56549), .D(n_17952)
		, .Z(n_36425));
	notech_ao4 i_17428561(.A(n_61340), .B(n_17778), .C(n_56549), .D(n_17953)
		, .Z(n_36419));
	notech_ao4 i_17328560(.A(n_61340), .B(n_17777), .C(n_56549), .D(n_17954)
		, .Z(n_36413));
	notech_ao4 i_17228559(.A(n_61344), .B(n_17776), .C(n_56549), .D(n_17955)
		, .Z(n_36407));
	notech_ao4 i_17128558(.A(n_61344), .B(n_17775), .C(n_56549), .D(n_17956)
		, .Z(n_36401));
	notech_ao4 i_17028557(.A(n_61344), .B(n_17774), .C(n_56549), .D(n_17957)
		, .Z(n_36395));
	notech_ao4 i_16928556(.A(n_61344), .B(n_17773), .C(n_56549), .D(n_17958)
		, .Z(n_36389));
	notech_ao4 i_16828555(.A(n_61340), .B(n_17772), .C(n_56549), .D(n_17959)
		, .Z(n_36383));
	notech_ao4 i_16728554(.A(n_61340), .B(n_17771), .C(n_56549), .D(n_17960)
		, .Z(n_36377));
	notech_ao4 i_16628553(.A(n_61340), .B(n_17770), .C(n_56549), .D(n_17961)
		, .Z(n_36371));
	notech_ao4 i_16528552(.A(n_61340), .B(n_17769), .C(n_56549), .D(n_17962)
		, .Z(n_36365));
	notech_ao4 i_16428551(.A(n_61340), .B(n_17768), .C(n_56549), .D(n_17963)
		, .Z(n_36359));
	notech_ao4 i_16328550(.A(n_61340), .B(n_17767), .C(n_56549), .D(n_17964)
		, .Z(n_36353));
	notech_ao4 i_16228549(.A(n_61340), .B(n_17766), .C(n_56549), .D(n_17965)
		, .Z(n_36347));
	notech_ao4 i_16128548(.A(n_61340), .B(n_17765), .C(n_56549), .D(n_17966)
		, .Z(n_36341));
	notech_ao4 i_16028547(.A(n_61301), .B(n_17764), .C(n_56556), .D(n_17967)
		, .Z(n_36335));
	notech_ao4 i_15928546(.A(n_61301), .B(n_17763), .C(n_56556), .D(n_17968)
		, .Z(n_36329));
	notech_ao4 i_15828545(.A(n_61301), .B(n_17762), .C(n_56556), .D(n_17969)
		, .Z(n_36323));
	notech_ao4 i_15728544(.A(n_61301), .B(n_17761), .C(n_56556), .D(n_17970)
		, .Z(n_36317));
	notech_ao4 i_15628543(.A(n_61331), .B(n_17760), .C(n_56556), .D(n_17868)
		, .Z(n_36311));
	notech_ao4 i_15528542(.A(n_61331), .B(n_17759), .C(n_56556), .D(n_17971)
		, .Z(n_36305));
	notech_ao4 i_15428541(.A(n_61301), .B(n_17758), .C(n_56556), .D(n_17972)
		, .Z(n_36299));
	notech_ao4 i_15328540(.A(n_61331), .B(n_17757), .C(n_56556), .D(n_17973)
		, .Z(n_36293));
	notech_ao4 i_15228539(.A(n_61301), .B(n_17756), .C(n_56556), .D(n_17974)
		, .Z(n_36287));
	notech_ao4 i_15128538(.A(n_61301), .B(n_17755), .C(n_56556), .D(n_17975)
		, .Z(n_36281));
	notech_ao4 i_15028537(.A(n_61301), .B(n_17754), .C(n_56556), .D(n_17976)
		, .Z(n_36275));
	notech_ao4 i_14928536(.A(n_61301), .B(n_17753), .C(n_56556), .D(n_17977)
		, .Z(n_36269));
	notech_ao4 i_14828535(.A(n_61301), .B(n_17752), .C(n_56556), .D(n_17869)
		, .Z(n_36263));
	notech_ao4 i_14728534(.A(n_61301), .B(n_17751), .C(n_56556), .D(n_17995)
		, .Z(n_36257));
	notech_ao4 i_14628533(.A(n_61301), .B(n_17750), .C(n_56556), .D(n_17978)
		, .Z(n_36251));
	notech_ao4 i_14528532(.A(n_61301), .B(n_17749), .C(n_56556), .D(n_17979)
		, .Z(n_36245));
	notech_ao4 i_14428531(.A(n_61331), .B(n_17748), .C(n_56554), .D(n_17980)
		, .Z(n_36239));
	notech_ao4 i_14328530(.A(n_61331), .B(n_17747), .C(n_56554), .D(n_17981)
		, .Z(n_36233));
	notech_ao4 i_14228529(.A(n_61331), .B(n_17746), .C(n_56554), .D(n_17994)
		, .Z(n_36227));
	notech_ao4 i_14128528(.A(n_61331), .B(n_17745), .C(n_56554), .D(n_17993)
		, .Z(n_36221));
	notech_ao4 i_14028527(.A(n_61335), .B(n_17744), .C(n_56554), .D(n_17870)
		, .Z(n_36215));
	notech_ao4 i_13928526(.A(n_61335), .B(n_17743), .C(n_56554), .D(n_17982)
		, .Z(n_36209));
	notech_ao4 i_13828525(.A(n_56554), .B(n_17983), .C(n_61335), .D(n_17742)
		, .Z(n_36203));
	notech_ao4 i_13728524(.A(n_61335), .B(n_17741), .C(n_56554), .D(n_17984)
		, .Z(n_36197));
	notech_ao4 i_13628523(.A(n_61331), .B(n_17740), .C(n_56554), .D(n_17985)
		, .Z(n_36191));
	notech_ao4 i_13528522(.A(n_61331), .B(n_17739), .C(n_56554), .D(n_17986)
		, .Z(n_36185));
	notech_ao4 i_13428521(.A(n_61331), .B(n_17738), .C(n_56554), .D(n_17987)
		, .Z(n_36179));
	notech_ao4 i_13328520(.A(n_61331), .B(n_17737), .C(n_56554), .D(n_17988)
		, .Z(n_36173));
	notech_ao4 i_13228519(.A(n_61331), .B(n_17736), .C(n_56554), .D(n_17871)
		, .Z(n_36167));
	notech_ao4 i_13128518(.A(n_61331), .B(n_17735), .C(n_56554), .D(n_17992)
		, .Z(n_36161));
	notech_ao4 i_13028517(.A(n_61331), .B(n_17734), .C(n_56554), .D(n_17989)
		, .Z(n_36155));
	notech_ao4 i_12928516(.A(n_61331), .B(n_17733), .C(n_56554), .D(n_17990)
		, .Z(n_36149));
	notech_nand3 i_86434066(.A(n_3086), .B(n_60101), .C(queue[36]), .Z(n_1577
		));
	notech_and4 i_2824994(.A(n_2357), .B(n_2356), .C(n_2351), .D(n_2355), .Z
		(squeue_27101060));
	notech_nand3 i_84634084(.A(n_59659), .B(n_59931), .C(queue[27]), .Z(n_1574
		));
	notech_nand3 i_83334097(.A(n_3086), .B(n_60097), .C(queue[35]), .Z(n_1561
		));
	notech_and4 i_2724993(.A(n_2343), .B(n_2342), .C(n_2337), .D(n_2341), .Z
		(squeue_26101061));
	notech_nand3 i_81534115(.A(n_59659), .B(n_59933), .C(queue[26]), .Z(n_1558
		));
	notech_nand3 i_80234128(.A(n_61405), .B(n_60097), .C(queue[34]), .Z(n_1545
		));
	notech_and4 i_2624992(.A(n_2329), .B(n_2328), .C(n_2323), .D(n_2327), .Z
		(squeue_25101062));
	notech_nand3 i_78434146(.A(n_59659), .B(n_59933), .C(queue[25]), .Z(n_1542
		));
	notech_nand3 i_77134159(.A(n_61405), .B(n_60097), .C(queue[33]), .Z(n_1529
		));
	notech_and4 i_2524991(.A(n_2315), .B(n_2314), .C(n_2309), .D(n_2313), .Z
		(squeue_24101063));
	notech_nand3 i_75334177(.A(n_59659), .B(n_59933), .C(queue[24]), .Z(n_1526
		));
	notech_nand3 i_74034190(.A(n_61405), .B(n_60101), .C(queue[32]), .Z(n_1513
		));
	notech_and4 i_2424990(.A(n_2301), .B(n_2300), .C(n_2295), .D(n_2299), .Z
		(squeue_23101064));
	notech_nand3 i_72234208(.A(n_59659), .B(n_59933), .C(queue[23]), .Z(n_1510
		));
	notech_or2 i_70934221(.A(n_59988), .B(n_17322), .Z(n_1497));
	notech_and4 i_2324989(.A(n_2287), .B(n_2286), .C(n_2281), .D(n_2285), .Z
		(squeue_22101065));
	notech_nand3 i_69134239(.A(n_59659), .B(n_59931), .C(queue[22]), .Z(n_1494
		));
	notech_nand3 i_67834252(.A(n_61409), .B(n_60097), .C(queue[30]), .Z(n_1481
		));
	notech_and4 i_2224988(.A(n_2273), .B(n_2272), .C(n_2267), .D(n_2271), .Z
		(squeue_21101066));
	notech_nand3 i_66034270(.A(n_59659), .B(n_59931), .C(queue[21]), .Z(n_1478
		));
	notech_nand3 i_64734283(.A(n_61409), .B(n_60097), .C(queue[29]), .Z(n_1465
		));
	notech_and4 i_2124987(.A(n_2259), .B(n_2258), .C(n_2253), .D(n_2257), .Z
		(squeue_20101067));
	notech_nand3 i_62934301(.A(n_59659), .B(n_59933), .C(queue[20]), .Z(n_1462
		));
	notech_nand3 i_61634314(.A(n_61405), .B(n_60097), .C(queue[28]), .Z(n_1449
		));
	notech_and4 i_2024986(.A(n_2245), .B(n_2244), .C(n_2239), .D(n_2243), .Z
		(squeue_19101068));
	notech_nand3 i_59834332(.A(n_59659), .B(n_59931), .C(queue[19]), .Z(n_1446
		));
	notech_nand3 i_58534345(.A(n_61405), .B(n_60097), .C(queue[27]), .Z(n_1433
		));
	notech_and4 i_1924985(.A(n_2231), .B(n_2230), .C(n_2225), .D(n_2229), .Z
		(squeue_18101069));
	notech_nand3 i_56734363(.A(n_59659), .B(n_59931), .C(queue[18]), .Z(n_1430
		));
	notech_nand2 i_8034959(.A(wptr[0]), .B(n_17301), .Z(n_52860135));
	notech_ao3 i_5047(.A(n_17301), .B(n_17291), .C(n_62847), .Z(n_52960136)
		);
	notech_reg fault_wptr_en_reg(.CP(n_63396), .D(n_15349), .CD(n_62700), .Q
		(fault_wptr_en));
	notech_mux2 i_21790(.S(n_35236), .A(fault_wptr_en), .B(n_17293), .Z(n_15349
		));
	notech_reg addrf_reg_0(.CP(n_63396), .D(iaddr[0]), .CD(n_62700), .Q(addrf
		[0]));
	notech_reg addrf_reg_1(.CP(n_63396), .D(iaddr[1]), .CD(n_62700), .Q(addrf
		[1]));
	notech_reg addrf_reg_2(.CP(n_63396), .D(iaddr[2]), .CD(n_62700), .Q(addrf
		[2]));
	notech_reg addrf_reg_3(.CP(n_63396), .D(iaddr[3]), .CD(n_62700), .Q(addrf
		[3]));
	notech_reg addrf_reg_4(.CP(n_63396), .D(iaddr[4]), .CD(n_62701), .Q(addrf
		[4]));
	notech_reg addrf_reg_5(.CP(n_63396), .D(iaddr[5]), .CD(n_62701), .Q(addrf
		[5]));
	notech_reg addrf_reg_6(.CP(n_63396), .D(iaddr[6]), .CD(n_62701), .Q(addrf
		[6]));
	notech_reg addrf_reg_7(.CP(n_63396), .D(iaddr[7]), .CD(n_62700), .Q(addrf
		[7]));
	notech_reg addrf_reg_8(.CP(n_63396), .D(iaddr[8]), .CD(n_62701), .Q(addrf
		[8]));
	notech_reg addrf_reg_9(.CP(n_63396), .D(iaddr[9]), .CD(n_62700), .Q(addrf
		[9]));
	notech_reg addrf_reg_10(.CP(n_63484), .D(iaddr[10]), .CD(n_62700), .Q(addrf
		[10]));
	notech_reg addrf_reg_11(.CP(n_63484), .D(iaddr[11]), .CD(n_62700), .Q(addrf
		[11]));
	notech_reg addrf_reg_12(.CP(n_63484), .D(iaddr[12]), .CD(n_62699), .Q(addrf
		[12]));
	notech_reg addrf_reg_13(.CP(n_63484), .D(iaddr[13]), .CD(n_62699), .Q(addrf
		[13]));
	notech_reg addrf_reg_14(.CP(n_63484), .D(iaddr[14]), .CD(n_62699), .Q(addrf
		[14]));
	notech_reg addrf_reg_15(.CP(n_63484), .D(iaddr[15]), .CD(n_62700), .Q(addrf
		[15]));
	notech_reg addrf_reg_16(.CP(n_63484), .D(iaddr[16]), .CD(n_62700), .Q(addrf
		[16]));
	notech_reg addrf_reg_17(.CP(n_63484), .D(iaddr[17]), .CD(n_62700), .Q(addrf
		[17]));
	notech_reg addrf_reg_18(.CP(n_63484), .D(iaddr[18]), .CD(n_62700), .Q(addrf
		[18]));
	notech_reg addrf_reg_19(.CP(n_63484), .D(iaddr[19]), .CD(n_62700), .Q(addrf
		[19]));
	notech_reg addrf_reg_20(.CP(n_63484), .D(iaddr[20]), .CD(n_62701), .Q(addrf
		[20]));
	notech_reg addrf_reg_21(.CP(n_63484), .D(iaddr[21]), .CD(n_62702), .Q(addrf
		[21]));
	notech_reg addrf_reg_22(.CP(n_63484), .D(iaddr[22]), .CD(n_62702), .Q(addrf
		[22]));
	notech_reg addrf_reg_23(.CP(n_63484), .D(iaddr[23]), .CD(n_62702), .Q(addrf
		[23]));
	notech_reg addrf_reg_24(.CP(n_63484), .D(iaddr[24]), .CD(n_62702), .Q(addrf
		[24]));
	notech_reg addrf_reg_25(.CP(n_63484), .D(iaddr[25]), .CD(n_62702), .Q(addrf
		[25]));
	notech_reg addrf_reg_26(.CP(n_63484), .D(iaddr[26]), .CD(n_62702), .Q(addrf
		[26]));
	notech_reg addrf_reg_27(.CP(n_63484), .D(iaddr[27]), .CD(n_62702), .Q(addrf
		[27]));
	notech_reg addrf_reg_28(.CP(n_63484), .D(iaddr[28]), .CD(n_62702), .Q(addrf
		[28]));
	notech_reg addrf_reg_29(.CP(n_63482), .D(iaddr[29]), .CD(n_62702), .Q(addrf
		[29]));
	notech_reg addrf_reg_30(.CP(n_63482), .D(iaddr[30]), .CD(n_62702), .Q(addrf
		[30]));
	notech_reg addrf_reg_31(.CP(n_63558), .D(iaddr[31]), .CD(n_62702), .Q(addrf
		[31]));
	notech_reg code_req_reg(.CP(n_63558), .D(n_15419), .CD(n_62701), .Q(n_62863
		));
	notech_mux2 i_21926(.S(n_36936), .A(n_62847), .B(n_52960136), .Z(n_15419
		));
	notech_reg addrshft_reg_0(.CP(n_63558), .D(n_15425), .CD(n_62701), .Q(addrshft
		[0]));
	notech_mux2 i_21934(.S(\nbus_12118[0] ), .A(addrshft[0]), .B(n_35323), .Z
		(n_15425));
	notech_reg addrshft_reg_1(.CP(n_63558), .D(n_15431), .CD(n_62701), .Q(addrshft
		[1]));
	notech_mux2 i_21942(.S(\nbus_12118[0] ), .A(addrshft[1]), .B(n_35329), .Z
		(n_15431));
	notech_reg addrshft_reg_2(.CP(n_63558), .D(n_15437), .CD(n_62701), .Q(addrshft
		[2]));
	notech_mux2 i_21950(.S(\nbus_12118[0] ), .A(addrshft[2]), .B(n_35335), .Z
		(n_15437));
	notech_reg addrshft_reg_3(.CP(n_63558), .D(n_15443), .CD(n_62701), .Q(addrshft
		[3]));
	notech_mux2 i_21958(.S(\nbus_12118[0] ), .A(addrshft[3]), .B(n_35341), .Z
		(n_15443));
	notech_reg addrshft_reg_4(.CP(n_63558), .D(n_15449), .CD(n_62701), .Q(addrshft
		[4]));
	notech_mux2 i_21966(.S(\nbus_12118[0] ), .A(addrshft[4]), .B(n_26059867)
		, .Z(n_15449));
	notech_reg addrshft_reg_5(.CP(n_63558), .D(n_15455), .CD(n_62702), .Q(addrshft
		[5]));
	notech_mux2 i_21974(.S(\nbus_12118[0] ), .A(addrshft[5]), .B(n_17299), .Z
		(n_15455));
	notech_reg wptr_reg_0(.CP(n_63558), .D(n_15461), .CD(n_62701), .Q(wptr[0
		]));
	notech_mux2 i_21982(.S(n_17302), .A(wptr[0]), .B(n_31459921), .Z(n_15461
		));
	notech_reg wptr_reg_1(.CP(n_63558), .D(n_15467), .CD(n_62701), .Q(wptr[1
		]));
	notech_mux2 i_21990(.S(n_17302), .A(n_61424), .B(n_35229), .Z(n_15467)
		);
	notech_nand3 i_55434376(.A(n_61405), .B(n_60097), .C(queue[26]), .Z(n_1417
		));
	notech_reg fault_wptr_reg_0(.CP(n_63558), .D(n_15473), .CD(n_62701), .Q(fault_wptr
		[0]));
	notech_mux2 i_21998(.S(\nbus_12115[0] ), .A(fault_wptr[0]), .B(n_17303),
		 .Z(n_15473));
	notech_reg fault_wptr_reg_1(.CP(n_63558), .D(n_15479), .CD(n_62696), .Q(fault_wptr
		[1]));
	notech_mux2 i_22006(.S(\nbus_12115[0] ), .A(fault_wptr[1]), .B(n_17304),
		 .Z(n_15479));
	notech_reg pc_pg_fault_reg(.CP(n_63558), .D(n_15485), .CD(n_62696), .Q(n_61444
		));
	notech_mux2 i_22014(.S(n_34969), .A(n_61438), .B(n_17297), .Z(n_15485)
		);
	notech_and4 i_1824984(.A(n_2217), .B(n_2216), .C(n_2211), .D(n_2215), .Z
		(squeue_17101070));
	notech_reg purge_cnt_reg_0(.CP(n_63558), .D(n_15491), .CD(n_62696), .Q(purge_cnt
		[0]));
	notech_mux2 i_22022(.S(\nbus_12117[0] ), .A(purge_cnt[0]), .B(n_30359910
		), .Z(n_15491));
	notech_nand3 i_53634394(.A(n_59657), .B(n_59928), .C(queue[17]), .Z(n_1414
		));
	notech_reg purge_cnt_reg_1(.CP(n_63558), .D(n_15497), .CD(n_62696), .Q(purge_cnt
		[1]));
	notech_mux2 i_22030(.S(\nbus_12117[0] ), .A(purge_cnt[1]), .B(n_30459911
		), .Z(n_15497));
	notech_reg purge_cnt_reg_2(.CP(n_63558), .D(n_15503), .CD(n_62696), .Q(purge_cnt
		[2]));
	notech_mux2 i_22038(.S(\nbus_12117[0] ), .A(purge_cnt[2]), .B(n_30559912
		), .Z(n_15503));
	notech_reg purge_cnt_reg_3(.CP(n_63558), .D(n_15509), .CD(n_62697), .Q(purge_cnt
		[3]));
	notech_mux2 i_22046(.S(\nbus_12117[0] ), .A(purge_cnt[3]), .B(n_30659913
		), .Z(n_15509));
	notech_reg purge_cnt_reg_4(.CP(n_63558), .D(n_15515), .CD(n_62697), .Q(purge_cnt
		[4]));
	notech_mux2 i_22054(.S(\nbus_12117[0] ), .A(purge_cnt[4]), .B(n_30759914
		), .Z(n_15515));
	notech_reg purge_cnt_reg_5(.CP(n_63482), .D(n_15521), .CD(n_62697), .Q(purge_cnt
		[5]));
	notech_mux2 i_22062(.S(\nbus_12117[0] ), .A(purge_cnt[5]), .B(n_30859915
		), .Z(n_15521));
	notech_reg purge_cnt_reg_6(.CP(n_63482), .D(n_15527), .CD(n_62696), .Q(purge_cnt
		[6]));
	notech_mux2 i_22070(.S(\nbus_12117[0] ), .A(purge_cnt[6]), .B(n_30959916
		), .Z(n_15527));
	notech_reg purge_cnt_reg_7(.CP(n_63482), .D(n_15533), .CD(n_62696), .Q(purge_cnt
		[7]));
	notech_mux2 i_22078(.S(\nbus_12117[0] ), .A(purge_cnt[7]), .B(n_31059917
		), .Z(n_15533));
	notech_reg purge_cnt_reg_8(.CP(n_63482), .D(n_15539), .CD(n_62696), .Q(purge_cnt
		[8]));
	notech_mux2 i_22086(.S(\nbus_12117[0] ), .A(purge_cnt[8]), .B(n_31159918
		), .Z(n_15539));
	notech_reg purge_cnt_reg_9(.CP(n_63482), .D(n_15545), .CD(n_62695), .Q(purge_cnt
		[9]));
	notech_mux2 i_22094(.S(\nbus_12117[0] ), .A(purge_cnt[9]), .B(n_31259919
		), .Z(n_15545));
	notech_reg purge_cnt_reg_10(.CP(n_63482), .D(n_15551), .CD(n_62696), .Q(purge_cnt
		[10]));
	notech_mux2 i_22102(.S(\nbus_12117[0] ), .A(purge_cnt[10]), .B(n_31359920
		), .Z(n_15551));
	notech_reg_set purge_reg(.CP(n_63482), .D(n_15557), .SD(n_62695), .Q(purge
		));
	notech_mux2 i_22110(.S(n_36919), .A(purge), .B(n_61438), .Z(n_15557));
	notech_reg addr_reg_0(.CP(n_63482), .D(n_15563), .CD(n_62695), .Q(iaddr[
		0]));
	notech_mux2 i_22118(.S(\nbus_12122[0] ), .A(iaddr[0]), .B(n_29959906), .Z
		(n_15563));
	notech_reg addr_reg_1(.CP(n_63482), .D(n_15569), .CD(n_62695), .Q(iaddr[
		1]));
	notech_mux2 i_22126(.S(\nbus_12122[0] ), .A(iaddr[1]), .B(n_30059907), .Z
		(n_15569));
	notech_nand3 i_52334407(.A(n_61405), .B(n_60097), .C(queue[25]), .Z(n_1401
		));
	notech_reg addr_reg_2(.CP(n_63558), .D(n_15575), .CD(n_62696), .Q(iaddr[
		2]));
	notech_mux2 i_22134(.S(\nbus_12122[0] ), .A(iaddr[2]), .B(n_30159908), .Z
		(n_15575));
	notech_reg addr_reg_3(.CP(n_63554), .D(n_15581), .CD(n_62696), .Q(iaddr[
		3]));
	notech_mux2 i_22142(.S(\nbus_12122[0] ), .A(iaddr[3]), .B(n_30259909), .Z
		(n_15581));
	notech_reg addr_reg_4(.CP(n_63480), .D(n_15587), .CD(n_62696), .Q(iaddr[
		4]));
	notech_mux2 i_22150(.S(\nbus_12122[0] ), .A(iaddr[4]), .B(n_36987), .Z(n_15587
		));
	notech_and4 i_1724983(.A(n_2203), .B(n_2202), .C(n_2197), .D(n_2201), .Z
		(squeue_16101071));
	notech_reg addr_reg_5(.CP(n_63554), .D(n_15593), .CD(n_62696), .Q(iaddr[
		5]));
	notech_mux2 i_22158(.S(\nbus_12122[0] ), .A(iaddr[5]), .B(n_36993), .Z(n_15593
		));
	notech_nand3 i_50534425(.A(n_59657), .B(n_59928), .C(queue[16]), .Z(n_1398
		));
	notech_reg addr_reg_6(.CP(n_63554), .D(n_15599), .CD(n_62696), .Q(iaddr[
		6]));
	notech_mux2 i_22166(.S(\nbus_12122[0] ), .A(iaddr[6]), .B(n_36999), .Z(n_15599
		));
	notech_reg addr_reg_7(.CP(n_63554), .D(n_15605), .CD(n_62697), .Q(iaddr[
		7]));
	notech_mux2 i_22174(.S(\nbus_12122[0] ), .A(iaddr[7]), .B(n_37005), .Z(n_15605
		));
	notech_reg addr_reg_8(.CP(n_63554), .D(n_15611), .CD(n_62699), .Q(iaddr[
		8]));
	notech_mux2 i_22182(.S(\nbus_12122[0] ), .A(iaddr[8]), .B(n_37011), .Z(n_15611
		));
	notech_reg addr_reg_9(.CP(n_63554), .D(n_15617), .CD(n_62699), .Q(iaddr[
		9]));
	notech_mux2 i_22190(.S(\nbus_12122[0] ), .A(iaddr[9]), .B(n_37017), .Z(n_15617
		));
	notech_reg_set addr_reg_10(.CP(n_63554), .D(n_15623), .SD(n_62699), .Q(iaddr
		[10]));
	notech_mux2 i_22198(.S(\nbus_12122[0] ), .A(iaddr[10]), .B(n_37023), .Z(n_15623
		));
	notech_reg_set addr_reg_11(.CP(n_63554), .D(n_15629), .SD(n_62699), .Q(iaddr
		[11]));
	notech_mux2 i_22206(.S(\nbus_12122[0] ), .A(iaddr[11]), .B(n_37029), .Z(n_15629
		));
	notech_reg_set addr_reg_12(.CP(n_63554), .D(n_15635), .SD(n_62699), .Q(iaddr
		[12]));
	notech_mux2 i_22214(.S(\nbus_12122[0] ), .A(iaddr[12]), .B(n_37035), .Z(n_15635
		));
	notech_reg_set addr_reg_13(.CP(n_63554), .D(n_15641), .SD(n_62699), .Q(iaddr
		[13]));
	notech_mux2 i_22222(.S(\nbus_12122[0] ), .A(iaddr[13]), .B(n_37041), .Z(n_15641
		));
	notech_reg_set addr_reg_14(.CP(n_63554), .D(n_15647), .SD(n_62699), .Q(iaddr
		[14]));
	notech_mux2 i_22230(.S(\nbus_12122[0] ), .A(iaddr[14]), .B(n_37047), .Z(n_15647
		));
	notech_reg_set addr_reg_15(.CP(n_63634), .D(n_15653), .SD(n_62699), .Q(iaddr
		[15]));
	notech_mux2 i_22238(.S(\nbus_12122[0] ), .A(iaddr[15]), .B(n_37053), .Z(n_15653
		));
	notech_reg_set addr_reg_16(.CP(n_63634), .D(n_15659), .SD(n_62699), .Q(iaddr
		[16]));
	notech_mux2 i_22246(.S(n_61290), .A(iaddr[16]), .B(n_37059), .Z(n_15659)
		);
	notech_reg_set addr_reg_17(.CP(n_63634), .D(n_15665), .SD(n_62699), .Q(iaddr
		[17]));
	notech_mux2 i_22254(.S(n_61290), .A(iaddr[17]), .B(n_37065), .Z(n_15665)
		);
	notech_reg_set addr_reg_18(.CP(n_63634), .D(n_15671), .SD(n_62699), .Q(iaddr
		[18]));
	notech_mux2 i_22262(.S(n_61290), .A(iaddr[18]), .B(n_37071), .Z(n_15671)
		);
	notech_or2 i_49234438(.A(n_59969), .B(n_17323), .Z(n_1385));
	notech_reg_set addr_reg_19(.CP(n_63634), .D(n_15677), .SD(n_62697), .Q(iaddr
		[19]));
	notech_mux2 i_22270(.S(n_61290), .A(iaddr[19]), .B(n_37077), .Z(n_15677)
		);
	notech_reg addr_reg_20(.CP(n_63634), .D(n_15683), .CD(n_62697), .Q(iaddr
		[20]));
	notech_mux2 i_22278(.S(n_61290), .A(iaddr[20]), .B(n_37083), .Z(n_15683)
		);
	notech_reg addr_reg_21(.CP(n_63634), .D(n_15689), .CD(n_62697), .Q(iaddr
		[21]));
	notech_mux2 i_22286(.S(n_61290), .A(iaddr[21]), .B(n_37089), .Z(n_15689)
		);
	notech_and4 i_1624982(.A(n_2189), .B(n_2188), .C(n_2183), .D(n_2187), .Z
		(squeue_15101072));
	notech_reg addr_reg_22(.CP(n_63634), .D(n_15695), .CD(n_62697), .Q(iaddr
		[22]));
	notech_mux2 i_22294(.S(n_61290), .A(iaddr[22]), .B(n_37095), .Z(n_15695)
		);
	notech_nand3 i_47434456(.A(n_59657), .B(n_59928), .C(queue[15]), .Z(n_1382
		));
	notech_reg addr_reg_23(.CP(n_63634), .D(n_15701), .CD(n_62697), .Q(iaddr
		[23]));
	notech_mux2 i_22302(.S(n_61290), .A(iaddr[23]), .B(n_37101), .Z(n_15701)
		);
	notech_reg addr_reg_24(.CP(n_63634), .D(n_15707), .CD(n_62697), .Q(iaddr
		[24]));
	notech_mux2 i_22310(.S(n_61290), .A(iaddr[24]), .B(n_37107), .Z(n_15707)
		);
	notech_reg addr_reg_25(.CP(n_63634), .D(n_15713), .CD(n_62697), .Q(iaddr
		[25]));
	notech_mux2 i_22318(.S(n_61290), .A(iaddr[25]), .B(n_37113), .Z(n_15713)
		);
	notech_reg addr_reg_26(.CP(n_63634), .D(n_15719), .CD(n_62697), .Q(iaddr
		[26]));
	notech_mux2 i_22326(.S(n_61290), .A(iaddr[26]), .B(n_37119), .Z(n_15719)
		);
	notech_reg addr_reg_27(.CP(n_63634), .D(n_15725), .CD(n_62697), .Q(iaddr
		[27]));
	notech_mux2 i_22334(.S(n_61290), .A(iaddr[27]), .B(n_37125), .Z(n_15725)
		);
	notech_reg addr_reg_28(.CP(n_63634), .D(n_15731), .CD(n_62697), .Q(iaddr
		[28]));
	notech_mux2 i_22342(.S(n_61290), .A(iaddr[28]), .B(n_37131), .Z(n_15731)
		);
	notech_reg addr_reg_29(.CP(n_63634), .D(n_15737), .CD(n_62707), .Q(iaddr
		[29]));
	notech_mux2 i_22350(.S(n_61290), .A(iaddr[29]), .B(n_37137), .Z(n_15737)
		);
	notech_reg addr_reg_30(.CP(n_63634), .D(n_15743), .CD(n_62708), .Q(iaddr
		[30]));
	notech_mux2 i_22358(.S(n_61290), .A(iaddr[30]), .B(n_37143), .Z(n_15743)
		);
	notech_reg addr_reg_31(.CP(n_63634), .D(n_15749), .CD(n_62707), .Q(iaddr
		[31]));
	notech_mux2 i_22366(.S(n_61290), .A(iaddr[31]), .B(n_37149), .Z(n_15749)
		);
	notech_reg queue_reg_0(.CP(n_63634), .D(n_15755), .CD(n_62707), .Q(queue
		[0]));
	notech_mux2 i_22374(.S(n_56603), .A(queue[0]), .B(n_35381), .Z(n_15755)
		);
	notech_reg queue_reg_1(.CP(n_63554), .D(n_15761), .CD(n_62707), .Q(queue
		[1]));
	notech_mux2 i_22382(.S(n_56603), .A(queue[1]), .B(n_35387), .Z(n_15761)
		);
	notech_reg queue_reg_2(.CP(n_63480), .D(n_15767), .CD(n_62708), .Q(queue
		[2]));
	notech_mux2 i_22390(.S(n_56603), .A(queue[2]), .B(n_35393), .Z(n_15767)
		);
	notech_reg queue_reg_3(.CP(n_63556), .D(n_15773), .CD(n_62708), .Q(queue
		[3]));
	notech_mux2 i_22398(.S(n_56603), .A(queue[3]), .B(n_35399), .Z(n_15773)
		);
	notech_or2 i_46134469(.A(n_59988), .B(n_17314), .Z(n_1369));
	notech_reg queue_reg_4(.CP(n_63556), .D(n_15779), .CD(n_62708), .Q(queue
		[4]));
	notech_mux2 i_22406(.S(n_56603), .A(queue[4]), .B(n_35405), .Z(n_15779)
		);
	notech_reg queue_reg_5(.CP(n_63556), .D(n_15785), .CD(n_62708), .Q(queue
		[5]));
	notech_mux2 i_22414(.S(n_56603), .A(queue[5]), .B(n_35411), .Z(n_15785)
		);
	notech_reg queue_reg_6(.CP(n_63556), .D(n_15791), .CD(n_62708), .Q(queue
		[6]));
	notech_mux2 i_22422(.S(n_56603), .A(queue[6]), .B(n_35417), .Z(n_15791)
		);
	notech_and4 i_1424980(.A(n_2175), .B(n_2174), .C(n_2169), .D(n_2173), .Z
		(squeue_13101073));
	notech_reg queue_reg_7(.CP(n_63556), .D(n_15797), .CD(n_62707), .Q(queue
		[7]));
	notech_mux2 i_22430(.S(n_56603), .A(queue[7]), .B(n_35423), .Z(n_15797)
		);
	notech_nand3 i_44334487(.A(n_59657), .B(n_59928), .C(queue[13]), .Z(n_1366
		));
	notech_reg queue_reg_8(.CP(n_63556), .D(n_15803), .CD(n_62707), .Q(queue
		[8]));
	notech_mux2 i_22438(.S(n_56603), .A(queue[8]), .B(n_35429), .Z(n_15803)
		);
	notech_reg queue_reg_9(.CP(n_63556), .D(n_15809), .CD(n_62707), .Q(queue
		[9]));
	notech_mux2 i_22446(.S(n_56603), .A(queue[9]), .B(n_35435), .Z(n_15809)
		);
	notech_reg queue_reg_10(.CP(n_63556), .D(n_15815), .CD(n_62707), .Q(queue
		[10]));
	notech_mux2 i_22454(.S(n_56603), .A(queue[10]), .B(n_35441), .Z(n_15815)
		);
	notech_reg queue_reg_11(.CP(n_63556), .D(n_15821), .CD(n_62706), .Q(queue
		[11]));
	notech_mux2 i_22462(.S(n_56603), .A(queue[11]), .B(n_35447), .Z(n_15821)
		);
	notech_reg queue_reg_12(.CP(n_63556), .D(n_15827), .CD(n_62707), .Q(queue
		[12]));
	notech_mux2 i_22470(.S(n_56603), .A(queue[12]), .B(n_35453), .Z(n_15827)
		);
	notech_reg queue_reg_13(.CP(n_63556), .D(n_15833), .CD(n_62707), .Q(queue
		[13]));
	notech_mux2 i_22478(.S(n_56603), .A(queue[13]), .B(n_35459), .Z(n_15833)
		);
	notech_reg queue_reg_14(.CP(n_63556), .D(n_15839), .CD(n_62707), .Q(queue
		[14]));
	notech_mux2 i_22486(.S(n_56603), .A(queue[14]), .B(n_35465), .Z(n_15839)
		);
	notech_reg queue_reg_15(.CP(n_63556), .D(n_15845), .CD(n_62707), .Q(queue
		[15]));
	notech_mux2 i_22494(.S(n_56603), .A(queue[15]), .B(n_35471), .Z(n_15845)
		);
	notech_reg queue_reg_16(.CP(n_63556), .D(n_15851), .CD(n_62707), .Q(queue
		[16]));
	notech_mux2 i_22502(.S(n_56601), .A(queue[16]), .B(n_35477), .Z(n_15851)
		);
	notech_reg queue_reg_17(.CP(n_63556), .D(n_15857), .CD(n_62707), .Q(queue
		[17]));
	notech_mux2 i_22510(.S(n_56601), .A(queue[17]), .B(n_35483), .Z(n_15857)
		);
	notech_reg queue_reg_18(.CP(n_63556), .D(n_15863), .CD(n_62708), .Q(queue
		[18]));
	notech_mux2 i_22518(.S(n_56601), .A(queue[18]), .B(n_35489), .Z(n_15863)
		);
	notech_reg queue_reg_19(.CP(n_63556), .D(n_15869), .CD(n_62709), .Q(queue
		[19]));
	notech_mux2 i_22526(.S(n_56601), .A(queue[19]), .B(n_35495), .Z(n_15869)
		);
	notech_reg queue_reg_20(.CP(n_63556), .D(n_15875), .CD(n_62709), .Q(queue
		[20]));
	notech_mux2 i_22534(.S(n_56601), .A(queue[20]), .B(n_35501), .Z(n_15875)
		);
	notech_nand3 i_43034500(.A(n_61405), .B(n_60097), .C(queue[21]), .Z(n_1353
		));
	notech_reg queue_reg_21(.CP(n_63556), .D(n_15881), .CD(n_62709), .Q(queue
		[21]));
	notech_mux2 i_22542(.S(n_56601), .A(queue[21]), .B(n_35507), .Z(n_15881)
		);
	notech_reg queue_reg_22(.CP(n_63480), .D(n_15887), .CD(n_62709), .Q(queue
		[22]));
	notech_mux2 i_22550(.S(n_56601), .A(queue[22]), .B(n_35513), .Z(n_15887)
		);
	notech_reg queue_reg_23(.CP(n_63480), .D(n_15893), .CD(n_62709), .Q(queue
		[23]));
	notech_mux2 i_22558(.S(n_56601), .A(queue[23]), .B(n_35519), .Z(n_15893)
		);
	notech_and4 i_1324979(.A(n_2161), .B(n_2160), .C(n_2155), .D(n_2159), .Z
		(squeue_12101074));
	notech_reg queue_reg_24(.CP(n_63480), .D(n_15899), .CD(n_62709), .Q(queue
		[24]));
	notech_mux2 i_22566(.S(n_56601), .A(queue[24]), .B(n_35525), .Z(n_15899)
		);
	notech_nand3 i_41234518(.A(n_59657), .B(n_59928), .C(queue[12]), .Z(n_1350
		));
	notech_reg queue_reg_25(.CP(n_63480), .D(n_15905), .CD(n_62709), .Q(queue
		[25]));
	notech_mux2 i_22574(.S(n_56601), .A(queue[25]), .B(n_35531), .Z(n_15905)
		);
	notech_reg queue_reg_26(.CP(n_63480), .D(n_15911), .CD(n_62709), .Q(queue
		[26]));
	notech_mux2 i_22582(.S(n_56601), .A(queue[26]), .B(n_35537), .Z(n_15911)
		);
	notech_reg queue_reg_27(.CP(n_63480), .D(n_15917), .CD(n_62709), .Q(queue
		[27]));
	notech_mux2 i_22590(.S(n_56601), .A(queue[27]), .B(n_35543), .Z(n_15917)
		);
	notech_reg queue_reg_28(.CP(n_63480), .D(n_15923), .CD(n_62709), .Q(queue
		[28]));
	notech_mux2 i_22598(.S(n_56601), .A(queue[28]), .B(n_35549), .Z(n_15923)
		);
	notech_reg queue_reg_29(.CP(n_63480), .D(n_15929), .CD(n_62709), .Q(queue
		[29]));
	notech_mux2 i_22606(.S(n_56601), .A(queue[29]), .B(n_35555), .Z(n_15929)
		);
	notech_reg queue_reg_30(.CP(n_63480), .D(n_15935), .CD(n_62708), .Q(queue
		[30]));
	notech_mux2 i_22614(.S(n_56601), .A(queue[30]), .B(n_35561), .Z(n_15935)
		);
	notech_reg queue_reg_31(.CP(n_63634), .D(n_15941), .CD(n_62708), .Q(queue
		[31]));
	notech_mux2 i_22622(.S(n_56601), .A(queue[31]), .B(n_35567), .Z(n_15941)
		);
	notech_reg queue_reg_32(.CP(n_63548), .D(n_15947), .CD(n_62708), .Q(queue
		[32]));
	notech_mux2 i_22630(.S(n_56608), .A(queue[32]), .B(n_35573), .Z(n_15947)
		);
	notech_reg queue_reg_33(.CP(n_63548), .D(n_15953), .CD(n_62708), .Q(queue
		[33]));
	notech_mux2 i_22638(.S(n_56608), .A(queue[33]), .B(n_35579), .Z(n_15953)
		);
	notech_reg queue_reg_34(.CP(n_63548), .D(n_15959), .CD(n_62708), .Q(queue
		[34]));
	notech_mux2 i_22646(.S(n_56608), .A(queue[34]), .B(n_35585), .Z(n_15959)
		);
	notech_reg queue_reg_35(.CP(n_63548), .D(n_15965), .CD(n_62709), .Q(queue
		[35]));
	notech_mux2 i_22654(.S(n_56608), .A(queue[35]), .B(n_35591), .Z(n_15965)
		);
	notech_reg queue_reg_36(.CP(n_63548), .D(n_15971), .CD(n_62709), .Q(queue
		[36]));
	notech_mux2 i_22662(.S(n_56608), .A(queue[36]), .B(n_35597), .Z(n_15971)
		);
	notech_reg queue_reg_37(.CP(n_63548), .D(n_15977), .CD(n_62709), .Q(queue
		[37]));
	notech_mux2 i_22670(.S(n_56608), .A(queue[37]), .B(n_35603), .Z(n_15977)
		);
	notech_nand3 i_39934531(.A(n_61405), .B(n_60101), .C(queue[20]), .Z(n_1337
		));
	notech_reg queue_reg_38(.CP(n_63548), .D(n_15983), .CD(n_62708), .Q(queue
		[38]));
	notech_mux2 i_22678(.S(n_56608), .A(queue[38]), .B(n_35609), .Z(n_15983)
		);
	notech_reg queue_reg_39(.CP(n_63548), .D(n_15989), .CD(n_62708), .Q(queue
		[39]));
	notech_mux2 i_22686(.S(n_56608), .A(queue[39]), .B(n_35615), .Z(n_15989)
		);
	notech_reg queue_reg_40(.CP(n_63548), .D(n_15995), .CD(n_62703), .Q(queue
		[40]));
	notech_mux2 i_22694(.S(n_56608), .A(queue[40]), .B(n_35621), .Z(n_15995)
		);
	notech_and4 i_1224978(.A(n_2147), .B(n_2146), .C(n_2141), .D(n_2145), .Z
		(squeue_11101075));
	notech_reg queue_reg_41(.CP(n_63548), .D(n_16001), .CD(n_62703), .Q(queue
		[41]));
	notech_mux2 i_22702(.S(n_56608), .A(queue[41]), .B(n_35627), .Z(n_16001)
		);
	notech_nand3 i_38134549(.A(n_59657), .B(n_59928), .C(queue[11]), .Z(n_1334
		));
	notech_reg queue_reg_42(.CP(n_63548), .D(n_16007), .CD(n_62703), .Q(queue
		[42]));
	notech_mux2 i_22710(.S(n_56608), .A(queue[42]), .B(n_35633), .Z(n_16007)
		);
	notech_reg queue_reg_43(.CP(n_63630), .D(n_16013), .CD(n_62703), .Q(queue
		[43]));
	notech_mux2 i_22718(.S(n_56608), .A(queue[43]), .B(n_35639), .Z(n_16013)
		);
	notech_reg queue_reg_44(.CP(n_63630), .D(n_16019), .CD(n_62703), .Q(queue
		[44]));
	notech_mux2 i_22726(.S(n_56608), .A(queue[44]), .B(n_35645), .Z(n_16019)
		);
	notech_reg queue_reg_45(.CP(n_63630), .D(n_16025), .CD(n_62705), .Q(queue
		[45]));
	notech_mux2 i_22734(.S(n_56608), .A(queue[45]), .B(n_35651), .Z(n_16025)
		);
	notech_reg queue_reg_46(.CP(n_63630), .D(n_16031), .CD(n_62705), .Q(queue
		[46]));
	notech_mux2 i_22742(.S(n_56608), .A(queue[46]), .B(n_35657), .Z(n_16031)
		);
	notech_reg queue_reg_47(.CP(n_63630), .D(n_16037), .CD(n_62705), .Q(queue
		[47]));
	notech_mux2 i_22750(.S(n_56608), .A(queue[47]), .B(n_35663), .Z(n_16037)
		);
	notech_reg queue_reg_48(.CP(n_63630), .D(n_16043), .CD(n_62705), .Q(queue
		[48]));
	notech_mux2 i_22758(.S(n_56606), .A(queue[48]), .B(n_35669), .Z(n_16043)
		);
	notech_reg queue_reg_49(.CP(n_63630), .D(n_16049), .CD(n_62705), .Q(queue
		[49]));
	notech_mux2 i_22766(.S(n_56606), .A(queue[49]), .B(n_35675), .Z(n_16049)
		);
	notech_reg queue_reg_50(.CP(n_63630), .D(n_16055), .CD(n_62703), .Q(queue
		[50]));
	notech_mux2 i_22774(.S(n_56606), .A(queue[50]), .B(n_35681), .Z(n_16055)
		);
	notech_reg queue_reg_51(.CP(n_63630), .D(n_16061), .CD(n_62703), .Q(queue
		[51]));
	notech_mux2 i_22782(.S(n_56606), .A(queue[51]), .B(n_35687), .Z(n_16061)
		);
	notech_reg queue_reg_52(.CP(n_63630), .D(n_16067), .CD(n_62703), .Q(queue
		[52]));
	notech_mux2 i_22790(.S(n_56606), .A(queue[52]), .B(n_35693), .Z(n_16067)
		);
	notech_reg queue_reg_53(.CP(n_63630), .D(n_16073), .CD(n_62703), .Q(queue
		[53]));
	notech_mux2 i_22798(.S(n_56606), .A(queue[53]), .B(n_35699), .Z(n_16073)
		);
	notech_reg queue_reg_54(.CP(n_63630), .D(n_16079), .CD(n_62702), .Q(queue
		[54]));
	notech_mux2 i_22806(.S(n_56606), .A(queue[54]), .B(n_35705), .Z(n_16079)
		);
	notech_nand3 i_36834562(.A(n_61409), .B(n_60101), .C(queue[19]), .Z(n_1320
		));
	notech_reg queue_reg_55(.CP(n_63630), .D(n_16085), .CD(n_62702), .Q(queue
		[55]));
	notech_mux2 i_22814(.S(n_56606), .A(queue[55]), .B(n_35711), .Z(n_16085)
		);
	notech_reg queue_reg_56(.CP(n_63630), .D(n_16091), .CD(n_62703), .Q(queue
		[56]));
	notech_mux2 i_22822(.S(n_56606), .A(queue[56]), .B(n_35717), .Z(n_16091)
		);
	notech_reg queue_reg_57(.CP(n_63630), .D(n_16097), .CD(n_62703), .Q(queue
		[57]));
	notech_mux2 i_22830(.S(n_56606), .A(queue[57]), .B(n_35723), .Z(n_16097)
		);
	notech_and4 i_1124977(.A(n_2133), .B(n_2132), .C(n_2127), .D(n_2131), .Z
		(squeue_10101076));
	notech_reg queue_reg_58(.CP(n_63630), .D(n_16103), .CD(n_62703), .Q(queue
		[58]));
	notech_mux2 i_22838(.S(n_56606), .A(queue[58]), .B(n_35729), .Z(n_16103)
		);
	notech_nand3 i_35034580(.A(n_59657), .B(n_59928), .C(queue[10]), .Z(n_1316
		));
	notech_reg queue_reg_59(.CP(n_63630), .D(n_16109), .CD(n_62703), .Q(queue
		[59]));
	notech_mux2 i_22846(.S(n_56606), .A(queue[59]), .B(n_35735), .Z(n_16109)
		);
	notech_reg queue_reg_60(.CP(n_63630), .D(n_16115), .CD(n_62703), .Q(queue
		[60]));
	notech_mux2 i_22854(.S(n_56606), .A(queue[60]), .B(n_35741), .Z(n_16115)
		);
	notech_reg queue_reg_61(.CP(n_63630), .D(n_16121), .CD(n_62705), .Q(queue
		[61]));
	notech_mux2 i_22862(.S(n_56606), .A(queue[61]), .B(n_35747), .Z(n_16121)
		);
	notech_reg queue_reg_62(.CP(n_63678), .D(n_16127), .CD(n_62706), .Q(queue
		[62]));
	notech_mux2 i_22870(.S(n_56606), .A(queue[62]), .B(n_35753), .Z(n_16127)
		);
	notech_reg queue_reg_63(.CP(n_63678), .D(n_16133), .CD(n_62706), .Q(queue
		[63]));
	notech_mux2 i_22878(.S(n_56606), .A(queue[63]), .B(n_35759), .Z(n_16133)
		);
	notech_reg queue_reg_64(.CP(n_63678), .D(n_16139), .CD(n_62706), .Q(queue
		[64]));
	notech_mux2 i_22886(.S(n_56593), .A(queue[64]), .B(n_35765), .Z(n_16139)
		);
	notech_reg queue_reg_65(.CP(n_63678), .D(n_16145), .CD(n_62706), .Q(queue
		[65]));
	notech_mux2 i_22894(.S(n_56593), .A(queue[65]), .B(n_35771), .Z(n_16145)
		);
	notech_reg queue_reg_66(.CP(n_63678), .D(n_16151), .CD(n_62706), .Q(queue
		[66]));
	notech_mux2 i_22902(.S(n_56593), .A(queue[66]), .B(n_35777), .Z(n_16151)
		);
	notech_reg queue_reg_67(.CP(n_63678), .D(n_16157), .CD(n_62706), .Q(queue
		[67]));
	notech_mux2 i_22910(.S(n_56593), .A(queue[67]), .B(n_35783), .Z(n_16157)
		);
	notech_reg queue_reg_68(.CP(n_63678), .D(n_16163), .CD(n_62706), .Q(queue
		[68]));
	notech_mux2 i_22918(.S(n_56593), .A(queue[68]), .B(n_35789), .Z(n_16163)
		);
	notech_reg queue_reg_69(.CP(n_63678), .D(n_16169), .CD(n_62706), .Q(queue
		[69]));
	notech_mux2 i_22926(.S(n_56593), .A(queue[69]), .B(n_35795), .Z(n_16169)
		);
	notech_reg queue_reg_70(.CP(n_63678), .D(n_16175), .CD(n_62706), .Q(queue
		[70]));
	notech_mux2 i_22934(.S(n_56593), .A(queue[70]), .B(n_35801), .Z(n_16175)
		);
	notech_reg queue_reg_71(.CP(n_63678), .D(n_16181), .CD(n_62706), .Q(queue
		[71]));
	notech_mux2 i_22942(.S(n_56593), .A(queue[71]), .B(n_35807), .Z(n_16181)
		);
	notech_nand3 i_33734593(.A(n_61409), .B(n_60101), .C(queue[18]), .Z(n_1293
		));
	notech_reg queue_reg_72(.CP(n_63678), .D(n_16187), .CD(n_62706), .Q(queue
		[72]));
	notech_mux2 i_22950(.S(n_56593), .A(queue[72]), .B(n_35813), .Z(n_16187)
		);
	notech_reg queue_reg_73(.CP(n_63678), .D(n_16193), .CD(n_62705), .Q(queue
		[73]));
	notech_mux2 i_22958(.S(n_56593), .A(queue[73]), .B(n_35819), .Z(n_16193)
		);
	notech_reg queue_reg_74(.CP(n_63678), .D(n_16199), .CD(n_62705), .Q(queue
		[74]));
	notech_mux2 i_22966(.S(n_56593), .A(queue[74]), .B(n_35825), .Z(n_16199)
		);
	notech_and4 i_1024976(.A(n_2119), .B(n_2118), .C(n_2113), .D(n_2117), .Z
		(squeue_9101077));
	notech_reg queue_reg_75(.CP(n_63678), .D(n_16205), .CD(n_62705), .Q(queue
		[75]));
	notech_mux2 i_22974(.S(n_56593), .A(queue[75]), .B(n_35831), .Z(n_16205)
		);
	notech_nand3 i_31934611(.A(n_59657), .B(n_59928), .C(queue[9]), .Z(n_1287
		));
	notech_reg queue_reg_76(.CP(n_63678), .D(n_16211), .CD(n_62705), .Q(queue
		[76]));
	notech_mux2 i_22982(.S(n_56593), .A(queue[76]), .B(n_35837), .Z(n_16211)
		);
	notech_reg queue_reg_77(.CP(n_63678), .D(n_16217), .CD(n_62705), .Q(queue
		[77]));
	notech_mux2 i_22990(.S(n_56593), .A(queue[77]), .B(n_35843), .Z(n_16217)
		);
	notech_reg queue_reg_78(.CP(n_63678), .D(n_16223), .CD(n_62706), .Q(queue
		[78]));
	notech_mux2 i_22998(.S(n_56593), .A(queue[78]), .B(n_35849), .Z(n_16223)
		);
	notech_reg queue_reg_79(.CP(n_63678), .D(n_16229), .CD(n_62706), .Q(queue
		[79]));
	notech_mux2 i_23006(.S(n_56593), .A(queue[79]), .B(n_35855), .Z(n_16229)
		);
	notech_reg queue_reg_80(.CP(n_63678), .D(n_16235), .CD(n_62705), .Q(queue
		[80]));
	notech_mux2 i_23014(.S(n_56591), .A(queue[80]), .B(n_35861), .Z(n_16235)
		);
	notech_reg queue_reg_81(.CP(n_63678), .D(n_16241), .CD(n_62705), .Q(queue
		[81]));
	notech_mux2 i_23022(.S(n_56591), .A(queue[81]), .B(n_35867), .Z(n_16241)
		);
	notech_reg queue_reg_82(.CP(n_63628), .D(n_16247), .CD(n_62705), .Q(queue
		[82]));
	notech_mux2 i_23030(.S(n_56591), .A(queue[82]), .B(n_35873), .Z(n_16247)
		);
	notech_reg queue_reg_83(.CP(n_63628), .D(n_16253), .CD(n_62695), .Q(queue
		[83]));
	notech_mux2 i_23038(.S(n_56591), .A(queue[83]), .B(n_35879), .Z(n_16253)
		);
	notech_reg queue_reg_84(.CP(n_63628), .D(n_16259), .CD(n_62685), .Q(queue
		[84]));
	notech_mux2 i_23046(.S(n_56591), .A(queue[84]), .B(n_35885), .Z(n_16259)
		);
	notech_reg queue_reg_85(.CP(n_63628), .D(n_16265), .CD(n_62685), .Q(queue
		[85]));
	notech_mux2 i_23054(.S(n_56591), .A(queue[85]), .B(n_35891), .Z(n_16265)
		);
	notech_reg queue_reg_86(.CP(n_63628), .D(n_16271), .CD(n_62685), .Q(queue
		[86]));
	notech_mux2 i_23062(.S(n_56591), .A(queue[86]), .B(n_35897), .Z(n_16271)
		);
	notech_reg queue_reg_87(.CP(n_63628), .D(n_16277), .CD(n_62685), .Q(queue
		[87]));
	notech_mux2 i_23070(.S(n_56591), .A(queue[87]), .B(n_35903), .Z(n_16277)
		);
	notech_reg queue_reg_88(.CP(n_63628), .D(n_16283), .CD(n_62685), .Q(queue
		[88]));
	notech_mux2 i_23078(.S(n_56591), .A(queue[88]), .B(n_35909), .Z(n_16283)
		);
	notech_nand3 i_30634624(.A(n_61409), .B(n_60101), .C(queue[17]), .Z(n_1273
		));
	notech_reg queue_reg_89(.CP(n_63628), .D(n_16289), .CD(n_62685), .Q(queue
		[89]));
	notech_mux2 i_23086(.S(n_56591), .A(queue[89]), .B(n_35915), .Z(n_16289)
		);
	notech_reg queue_reg_90(.CP(n_63628), .D(n_16295), .CD(n_62685), .Q(queue
		[90]));
	notech_mux2 i_23094(.S(n_56591), .A(queue[90]), .B(n_35921), .Z(n_16295)
		);
	notech_reg queue_reg_91(.CP(n_63628), .D(n_16301), .CD(n_62685), .Q(queue
		[91]));
	notech_mux2 i_23102(.S(n_56591), .A(queue[91]), .B(n_35927), .Z(n_16301)
		);
	notech_and4 i_924975(.A(n_2105), .B(n_2104), .C(n_2099), .D(n_2103), .Z(squeue_8101078
		));
	notech_reg queue_reg_92(.CP(n_63628), .D(n_16307), .CD(n_62685), .Q(queue
		[92]));
	notech_mux2 i_23110(.S(n_56591), .A(queue[92]), .B(n_35933), .Z(n_16307)
		);
	notech_nand3 i_28834642(.A(n_59657), .B(n_59931), .C(queue[8]), .Z(n_1270
		));
	notech_reg queue_reg_93(.CP(n_63628), .D(n_16313), .CD(n_62685), .Q(queue
		[93]));
	notech_mux2 i_23118(.S(n_56591), .A(queue[93]), .B(n_35939), .Z(n_16313)
		);
	notech_reg queue_reg_94(.CP(n_63632), .D(n_16319), .CD(n_62685), .Q(queue
		[94]));
	notech_mux2 i_23126(.S(n_56591), .A(queue[94]), .B(n_35945), .Z(n_16319)
		);
	notech_reg queue_reg_95(.CP(n_63550), .D(n_16325), .CD(n_62684), .Q(queue
		[95]));
	notech_mux2 i_23134(.S(n_56591), .A(queue[95]), .B(n_35951), .Z(n_16325)
		);
	notech_reg queue_reg_96(.CP(n_63550), .D(n_16331), .CD(n_62684), .Q(queue
		[96]));
	notech_mux2 i_23142(.S(n_56598), .A(queue[96]), .B(n_35957), .Z(n_16331)
		);
	notech_reg queue_reg_97(.CP(n_63550), .D(n_16337), .CD(n_62684), .Q(queue
		[97]));
	notech_mux2 i_23150(.S(n_56598), .A(queue[97]), .B(n_35963), .Z(n_16337)
		);
	notech_reg queue_reg_98(.CP(n_63550), .D(n_16343), .CD(n_62684), .Q(queue
		[98]));
	notech_mux2 i_23158(.S(n_56598), .A(queue[98]), .B(n_35969), .Z(n_16343)
		);
	notech_reg queue_reg_99(.CP(n_63550), .D(n_16349), .CD(n_62684), .Q(queue
		[99]));
	notech_mux2 i_23166(.S(n_56598), .A(queue[99]), .B(n_35975), .Z(n_16349)
		);
	notech_reg queue_reg_100(.CP(n_63550), .D(n_16355), .CD(n_62684), .Q(queue
		[100]));
	notech_mux2 i_23174(.S(n_56598), .A(queue[100]), .B(n_35981), .Z(n_16355
		));
	notech_reg queue_reg_101(.CP(n_63550), .D(n_16361), .CD(n_62685), .Q(queue
		[101]));
	notech_mux2 i_23182(.S(n_56598), .A(queue[101]), .B(n_35987), .Z(n_16361
		));
	notech_reg queue_reg_102(.CP(n_63550), .D(n_16367), .CD(n_62684), .Q(queue
		[102]));
	notech_mux2 i_23190(.S(n_56598), .A(queue[102]), .B(n_35993), .Z(n_16367
		));
	notech_reg queue_reg_103(.CP(n_63550), .D(n_16373), .CD(n_62684), .Q(queue
		[103]));
	notech_mux2 i_23198(.S(n_56598), .A(queue[103]), .B(n_35999), .Z(n_16373
		));
	notech_reg queue_reg_104(.CP(n_63632), .D(n_16379), .CD(n_62684), .Q(queue
		[104]));
	notech_mux2 i_23206(.S(n_56598), .A(queue[104]), .B(n_36005), .Z(n_16379
		));
	notech_reg queue_reg_105(.CP(n_63632), .D(n_16385), .CD(n_62685), .Q(queue
		[105]));
	notech_mux2 i_23214(.S(n_56598), .A(queue[105]), .B(n_36011), .Z(n_16385
		));
	notech_or2 i_27534655(.A(n_59950), .B(n_17323), .Z(n_1257));
	notech_reg queue_reg_106(.CP(n_63632), .D(n_16391), .CD(n_62688), .Q(queue
		[106]));
	notech_mux2 i_23222(.S(n_56598), .A(queue[106]), .B(n_36017), .Z(n_16391
		));
	notech_reg queue_reg_107(.CP(n_63632), .D(n_16397), .CD(n_62688), .Q(queue
		[107]));
	notech_mux2 i_23230(.S(n_56598), .A(queue[107]), .B(n_36023), .Z(n_16397
		));
	notech_reg queue_reg_108(.CP(n_63632), .D(n_16403), .CD(n_62687), .Q(queue
		[108]));
	notech_mux2 i_23238(.S(n_56598), .A(queue[108]), .B(n_36029), .Z(n_16403
		));
	notech_and4 i_724973(.A(n_2091), .B(n_2090), .C(n_2085), .D(n_2089), .Z(squeue_6101079
		));
	notech_reg queue_reg_109(.CP(n_63632), .D(n_16409), .CD(n_62687), .Q(queue
		[109]));
	notech_mux2 i_23246(.S(n_56598), .A(queue[109]), .B(n_36035), .Z(n_16409
		));
	notech_nand3 i_25734673(.A(n_59657), .B(n_59931), .C(queue[6]), .Z(n_1254
		));
	notech_reg queue_reg_110(.CP(n_63632), .D(n_16415), .CD(n_62687), .Q(queue
		[110]));
	notech_mux2 i_23254(.S(n_56598), .A(queue[110]), .B(n_36041), .Z(n_16415
		));
	notech_reg queue_reg_111(.CP(n_63632), .D(n_16421), .CD(n_62688), .Q(queue
		[111]));
	notech_mux2 i_23262(.S(n_56598), .A(queue[111]), .B(n_36047), .Z(n_16421
		));
	notech_reg queue_reg_112(.CP(n_63632), .D(n_16427), .CD(n_62688), .Q(queue
		[112]));
	notech_mux2 i_23270(.S(n_56596), .A(queue[112]), .B(n_36053), .Z(n_16427
		));
	notech_reg queue_reg_113(.CP(n_63632), .D(n_16433), .CD(n_62688), .Q(queue
		[113]));
	notech_mux2 i_23278(.S(n_56596), .A(queue[113]), .B(n_36059), .Z(n_16433
		));
	notech_reg queue_reg_114(.CP(n_63632), .D(n_16439), .CD(n_62688), .Q(queue
		[114]));
	notech_mux2 i_23286(.S(n_56596), .A(queue[114]), .B(n_36065), .Z(n_16439
		));
	notech_reg queue_reg_115(.CP(n_63632), .D(n_16445), .CD(n_62688), .Q(queue
		[115]));
	notech_mux2 i_23294(.S(n_56596), .A(queue[115]), .B(n_36071), .Z(n_16445
		));
	notech_reg queue_reg_116(.CP(n_63632), .D(n_16451), .CD(n_62687), .Q(queue
		[116]));
	notech_mux2 i_23302(.S(n_56596), .A(queue[116]), .B(n_36077), .Z(n_16451
		));
	notech_reg queue_reg_117(.CP(n_63632), .D(n_16457), .CD(n_62687), .Q(queue
		[117]));
	notech_mux2 i_23310(.S(n_56596), .A(queue[117]), .B(n_36083), .Z(n_16457
		));
	notech_reg queue_reg_118(.CP(n_63632), .D(n_16463), .CD(n_62687), .Q(queue
		[118]));
	notech_mux2 i_23318(.S(n_56596), .A(queue[118]), .B(n_36089), .Z(n_16463
		));
	notech_reg queue_reg_119(.CP(n_63632), .D(n_16469), .CD(n_62687), .Q(queue
		[119]));
	notech_mux2 i_23326(.S(n_56596), .A(queue[119]), .B(n_36095), .Z(n_16469
		));
	notech_reg queue_reg_120(.CP(n_63632), .D(n_16475), .CD(n_62687), .Q(queue
		[120]));
	notech_mux2 i_23334(.S(n_56596), .A(queue[120]), .B(n_36101), .Z(n_16475
		));
	notech_reg queue_reg_121(.CP(n_63632), .D(n_16481), .CD(n_62687), .Q(queue
		[121]));
	notech_mux2 i_23342(.S(n_56596), .A(queue[121]), .B(n_36107), .Z(n_16481
		));
	notech_reg queue_reg_122(.CP(n_63550), .D(n_16487), .CD(n_62687), .Q(queue
		[122]));
	notech_mux2 i_23350(.S(n_56596), .A(queue[122]), .B(n_36113), .Z(n_16487
		));
	notech_nand3 i_24434686(.A(queue[14]), .B(n_61409), .C(n_60101), .Z(n_1241
		));
	notech_reg queue_reg_123(.CP(n_63550), .D(n_16493), .CD(n_62687), .Q(queue
		[123]));
	notech_mux2 i_23358(.S(n_56596), .A(queue[123]), .B(n_36119), .Z(n_16493
		));
	notech_reg queue_reg_124(.CP(n_63552), .D(n_16499), .CD(n_62687), .Q(queue
		[124]));
	notech_mux2 i_23366(.S(n_56596), .A(queue[124]), .B(n_36125), .Z(n_16499
		));
	notech_reg queue_reg_125(.CP(n_63552), .D(n_16505), .CD(n_62687), .Q(queue
		[125]));
	notech_mux2 i_23374(.S(n_56596), .A(queue[125]), .B(n_36131), .Z(n_16505
		));
	notech_and4 i_624972(.A(n_2077), .B(n_2076), .C(n_2071), .D(n_2075), .Z(squeue_5101080
		));
	notech_reg queue_reg_126(.CP(n_63552), .D(n_16511), .CD(n_62687), .Q(queue
		[126]));
	notech_mux2 i_23382(.S(n_56596), .A(queue[126]), .B(n_36137), .Z(n_16511
		));
	notech_nand3 i_22634704(.A(n_59657), .B(n_59931), .C(queue[5]), .Z(n_1238
		));
	notech_reg queue_reg_127(.CP(n_63552), .D(n_16517), .CD(n_62682), .Q(queue
		[127]));
	notech_mux2 i_23390(.S(n_56596), .A(queue[127]), .B(n_36143), .Z(n_16517
		));
	notech_reg queue_reg_128(.CP(n_63552), .D(n_16523), .CD(n_62682), .Q(queue
		[128]));
	notech_mux2 i_23398(.S(n_56582), .A(queue[128]), .B(n_17420), .Z(n_16523
		));
	notech_reg queue_reg_129(.CP(n_63552), .D(n_16529), .CD(n_62682), .Q(queue
		[129]));
	notech_mux2 i_23406(.S(n_56582), .A(queue[129]), .B(n_17422), .Z(n_16529
		));
	notech_reg queue_reg_130(.CP(n_63552), .D(n_16535), .CD(n_62681), .Q(queue
		[130]));
	notech_mux2 i_23414(.S(n_56582), .A(queue[130]), .B(n_17424), .Z(n_16535
		));
	notech_reg queue_reg_131(.CP(n_63552), .D(n_16541), .CD(n_62681), .Q(queue
		[131]));
	notech_mux2 i_23422(.S(n_56582), .A(queue[131]), .B(n_17426), .Z(n_16541
		));
	notech_reg queue_reg_132(.CP(n_63552), .D(n_16547), .CD(n_62682), .Q(queue
		[132]));
	notech_mux2 i_23430(.S(n_56582), .A(queue[132]), .B(n_17428), .Z(n_16547
		));
	notech_reg queue_reg_133(.CP(n_63552), .D(n_16553), .CD(n_62682), .Q(queue
		[133]));
	notech_mux2 i_23438(.S(n_56582), .A(queue[133]), .B(n_17430), .Z(n_16553
		));
	notech_reg queue_reg_134(.CP(n_63552), .D(n_16559), .CD(n_62682), .Q(queue
		[134]));
	notech_mux2 i_23446(.S(n_56582), .A(queue[134]), .B(n_17432), .Z(n_16559
		));
	notech_reg queue_reg_135(.CP(n_63552), .D(n_16565), .CD(n_62682), .Q(queue
		[135]));
	notech_mux2 i_23454(.S(n_56582), .A(queue[135]), .B(n_17434), .Z(n_16565
		));
	notech_reg queue_reg_136(.CP(n_63552), .D(n_16571), .CD(n_62682), .Q(queue
		[136]));
	notech_mux2 i_23462(.S(n_56582), .A(queue[136]), .B(n_17436), .Z(n_16571
		));
	notech_reg queue_reg_137(.CP(n_63552), .D(n_16577), .CD(n_62681), .Q(queue
		[137]));
	notech_mux2 i_23470(.S(n_56582), .A(queue[137]), .B(n_17438), .Z(n_16577
		));
	notech_reg queue_reg_138(.CP(n_63552), .D(n_16583), .CD(n_62681), .Q(queue
		[138]));
	notech_mux2 i_23478(.S(n_56582), .A(queue[138]), .B(n_17440), .Z(n_16583
		));
	notech_reg queue_reg_139(.CP(n_63552), .D(n_16589), .CD(n_62681), .Q(queue
		[139]));
	notech_mux2 i_23486(.S(n_56582), .A(queue[139]), .B(n_17442), .Z(n_16589
		));
	notech_nand3 i_21334717(.A(n_61409), .B(n_60101), .C(queue[13]), .Z(n_122560143
		));
	notech_reg queue_reg_140(.CP(n_63552), .D(n_16595), .CD(n_62681), .Q(queue
		[140]));
	notech_mux2 i_23494(.S(n_56582), .A(queue[140]), .B(n_17444), .Z(n_16595
		));
	notech_reg queue_reg_141(.CP(n_63552), .D(n_16601), .CD(n_62681), .Q(queue
		[141]));
	notech_mux2 i_23502(.S(n_56582), .A(queue[141]), .B(n_17446), .Z(n_16601
		));
	notech_reg queue_reg_142(.CP(n_63552), .D(n_16607), .CD(n_62681), .Q(queue
		[142]));
	notech_mux2 i_23510(.S(n_56582), .A(queue[142]), .B(n_17448), .Z(n_16607
		));
	notech_and4 i_524971(.A(n_2063), .B(n_2062), .C(n_2057), .D(n_2061), .Z(squeue_4101081
		));
	notech_reg queue_reg_143(.CP(n_63478), .D(n_16613), .CD(n_62681), .Q(queue
		[143]));
	notech_mux2 i_23518(.S(n_56582), .A(queue[143]), .B(n_17450), .Z(n_16613
		));
	notech_nand3 i_19534735(.A(n_59657), .B(n_59931), .C(queue[4]), .Z(n_122260146
		));
	notech_reg queue_reg_144(.CP(n_63478), .D(n_16619), .CD(n_62681), .Q(queue
		[144]));
	notech_mux2 i_23526(.S(n_56580), .A(queue[144]), .B(n_17452), .Z(n_16619
		));
	notech_reg queue_reg_145(.CP(n_63478), .D(n_16625), .CD(n_62681), .Q(queue
		[145]));
	notech_mux2 i_23534(.S(n_56580), .A(queue[145]), .B(n_17454), .Z(n_16625
		));
	notech_reg queue_reg_146(.CP(n_63478), .D(n_16631), .CD(n_62681), .Q(queue
		[146]));
	notech_mux2 i_23542(.S(n_56580), .A(queue[146]), .B(n_17456), .Z(n_16631
		));
	notech_reg queue_reg_147(.CP(n_63478), .D(n_16637), .CD(n_62681), .Q(queue
		[147]));
	notech_mux2 i_23550(.S(n_56580), .A(queue[147]), .B(n_17458), .Z(n_16637
		));
	notech_reg queue_reg_148(.CP(n_63478), .D(n_16643), .CD(n_62682), .Q(queue
		[148]));
	notech_mux2 i_23558(.S(n_56580), .A(queue[148]), .B(n_17460), .Z(n_16643
		));
	notech_reg queue_reg_149(.CP(n_63478), .D(n_16649), .CD(n_62683), .Q(queue
		[149]));
	notech_mux2 i_23566(.S(n_56580), .A(queue[149]), .B(n_17462), .Z(n_16649
		));
	notech_reg queue_reg_150(.CP(n_63478), .D(n_16655), .CD(n_62683), .Q(queue
		[150]));
	notech_mux2 i_23574(.S(n_56580), .A(queue[150]), .B(n_17464), .Z(n_16655
		));
	notech_reg queue_reg_151(.CP(n_63478), .D(n_16661), .CD(n_62683), .Q(queue
		[151]));
	notech_mux2 i_23582(.S(n_56580), .A(queue[151]), .B(n_17466), .Z(n_16661
		));
	notech_reg queue_reg_152(.CP(n_63478), .D(n_16667), .CD(n_62683), .Q(queue
		[152]));
	notech_mux2 i_23590(.S(n_56580), .A(queue[152]), .B(n_17468), .Z(n_16667
		));
	notech_reg queue_reg_153(.CP(n_63478), .D(n_16673), .CD(n_62683), .Q(queue
		[153]));
	notech_mux2 i_23598(.S(n_56580), .A(queue[153]), .B(n_17470), .Z(n_16673
		));
	notech_reg queue_reg_154(.CP(n_63560), .D(n_16679), .CD(n_62684), .Q(queue
		[154]));
	notech_mux2 i_23606(.S(n_56580), .A(queue[154]), .B(n_17472), .Z(n_16679
		));
	notech_reg queue_reg_155(.CP(clk), .D(n_16685), .CD(n_62684), .Q(queue[
		155]));
	notech_mux2 i_23614(.S(n_56580), .A(queue[155]), .B(n_17474), .Z(n_16685
		));
	notech_reg queue_reg_156(.CP(clk), .D(n_16691), .CD(n_62684), .Q(queue[
		156]));
	notech_mux2 i_23622(.S(n_56580), .A(queue[156]), .B(n_17476), .Z(n_16691
		));
	notech_nand3 i_18234748(.A(n_61409), .B(n_60101), .C(queue[12]), .Z(n_120960159
		));
	notech_reg queue_reg_157(.CP(clk), .D(n_16697), .CD(n_62683), .Q(queue[
		157]));
	notech_mux2 i_23630(.S(n_56580), .A(queue[157]), .B(n_17478), .Z(n_16697
		));
	notech_reg queue_reg_158(.CP(clk), .D(n_16703), .CD(n_62684), .Q(queue[
		158]));
	notech_mux2 i_23638(.S(n_56580), .A(queue[158]), .B(n_17480), .Z(n_16703
		));
	notech_reg queue_reg_159(.CP(n_63490), .D(n_16709), .CD(n_62683), .Q(queue
		[159]));
	notech_mux2 i_23646(.S(n_56580), .A(queue[159]), .B(n_17482), .Z(n_16709
		));
	notech_and4 i_424970(.A(n_2049), .B(n_2048), .C(n_2043), .D(n_2047), .Z(squeue_3101082
		));
	notech_reg queue_reg_160(.CP(n_63490), .D(n_16715), .CD(n_62682), .Q(queue
		[160]));
	notech_mux2 i_23654(.S(n_56587), .A(queue[160]), .B(n_17484), .Z(n_16715
		));
	notech_nand3 i_16434766(.A(n_59657), .B(n_59928), .C(queue[3]), .Z(n_120660162
		));
	notech_reg queue_reg_161(.CP(n_63490), .D(n_16721), .CD(n_62683), .Q(queue
		[161]));
	notech_mux2 i_23662(.S(n_56587), .A(queue[161]), .B(n_17486), .Z(n_16721
		));
	notech_reg queue_reg_162(.CP(n_63490), .D(n_16727), .CD(n_62682), .Q(queue
		[162]));
	notech_mux2 i_23670(.S(n_56587), .A(queue[162]), .B(n_17488), .Z(n_16727
		));
	notech_reg queue_reg_163(.CP(n_63490), .D(n_16733), .CD(n_62682), .Q(queue
		[163]));
	notech_mux2 i_23678(.S(n_56587), .A(queue[163]), .B(n_17490), .Z(n_16733
		));
	notech_reg queue_reg_164(.CP(n_63490), .D(n_16739), .CD(n_62682), .Q(queue
		[164]));
	notech_mux2 i_23686(.S(n_56587), .A(queue[164]), .B(n_17492), .Z(n_16739
		));
	notech_reg queue_reg_165(.CP(n_63490), .D(n_16745), .CD(n_62683), .Q(queue
		[165]));
	notech_mux2 i_23694(.S(n_56587), .A(queue[165]), .B(n_17494), .Z(n_16745
		));
	notech_reg queue_reg_166(.CP(n_63490), .D(n_16751), .CD(n_62683), .Q(queue
		[166]));
	notech_mux2 i_23702(.S(n_56587), .A(queue[166]), .B(n_17496), .Z(n_16751
		));
	notech_reg queue_reg_167(.CP(n_63490), .D(n_16757), .CD(n_62683), .Q(queue
		[167]));
	notech_mux2 i_23710(.S(n_56587), .A(queue[167]), .B(n_17498), .Z(n_16757
		));
	notech_reg queue_reg_168(.CP(n_63490), .D(n_16763), .CD(n_62683), .Q(queue
		[168]));
	notech_mux2 i_23718(.S(n_56587), .A(queue[168]), .B(n_17500), .Z(n_16763
		));
	notech_reg queue_reg_169(.CP(n_63490), .D(n_16769), .CD(n_62683), .Q(queue
		[169]));
	notech_mux2 i_23726(.S(n_56587), .A(queue[169]), .B(n_17502), .Z(n_16769
		));
	notech_reg queue_reg_170(.CP(n_63490), .D(n_16775), .CD(n_62693), .Q(queue
		[170]));
	notech_mux2 i_23734(.S(n_56587), .A(queue[170]), .B(n_17504), .Z(n_16775
		));
	notech_reg queue_reg_171(.CP(n_63490), .D(n_16781), .CD(n_62693), .Q(queue
		[171]));
	notech_mux2 i_23742(.S(n_56587), .A(queue[171]), .B(n_17506), .Z(n_16781
		));
	notech_reg queue_reg_172(.CP(n_63490), .D(n_16787), .CD(n_62693), .Q(queue
		[172]));
	notech_mux2 i_23750(.S(n_56587), .A(queue[172]), .B(n_17508), .Z(n_16787
		));
	notech_reg queue_reg_173(.CP(n_63490), .D(n_16793), .CD(n_62693), .Q(queue
		[173]));
	notech_mux2 i_23758(.S(n_56587), .A(queue[173]), .B(n_17510), .Z(n_16793
		));
	notech_nand3 i_15134779(.A(n_61409), .B(n_60101), .C(queue[11]), .Z(n_119360175
		));
	notech_reg queue_reg_174(.CP(n_63490), .D(n_16799), .CD(n_62693), .Q(queue
		[174]));
	notech_mux2 i_23766(.S(n_56587), .A(queue[174]), .B(n_17512), .Z(n_16799
		));
	notech_reg queue_reg_175(.CP(n_63490), .D(n_16805), .CD(n_62693), .Q(queue
		[175]));
	notech_mux2 i_23774(.S(n_56587), .A(queue[175]), .B(n_17514), .Z(n_16805
		));
	notech_reg queue_reg_176(.CP(n_63490), .D(n_16811), .CD(n_62694), .Q(queue
		[176]));
	notech_mux2 i_23782(.S(n_56585), .A(queue[176]), .B(n_17516), .Z(n_16811
		));
	notech_and4 i_324969(.A(n_2035), .B(n_2034), .C(n_2029), .D(n_2033), .Z(squeue_2101083
		));
	notech_reg queue_reg_177(.CP(n_63490), .D(n_16817), .CD(n_62693), .Q(queue
		[177]));
	notech_mux2 i_23790(.S(n_56585), .A(queue[177]), .B(n_17518), .Z(n_16817
		));
	notech_nand3 i_13334797(.A(n_59657), .B(n_59928), .C(queue[2]), .Z(n_119060178
		));
	notech_reg queue_reg_178(.CP(n_63564), .D(n_16823), .CD(n_62693), .Q(queue
		[178]));
	notech_mux2 i_23798(.S(n_56585), .A(queue[178]), .B(n_17520), .Z(n_16823
		));
	notech_reg queue_reg_179(.CP(n_63488), .D(n_16829), .CD(n_62693), .Q(queue
		[179]));
	notech_mux2 i_23806(.S(n_56585), .A(queue[179]), .B(n_17522), .Z(n_16829
		));
	notech_reg queue_reg_180(.CP(n_63564), .D(n_16835), .CD(n_62693), .Q(queue
		[180]));
	notech_mux2 i_23814(.S(n_56585), .A(queue[180]), .B(n_17524), .Z(n_16835
		));
	notech_reg queue_reg_181(.CP(n_63564), .D(n_16841), .CD(n_62691), .Q(queue
		[181]));
	notech_mux2 i_23822(.S(n_56585), .A(queue[181]), .B(n_17526), .Z(n_16841
		));
	notech_reg queue_reg_182(.CP(n_63564), .D(n_16847), .CD(n_62691), .Q(queue
		[182]));
	notech_mux2 i_23830(.S(n_56585), .A(queue[182]), .B(n_17528), .Z(n_16847
		));
	notech_reg queue_reg_183(.CP(n_63564), .D(n_16853), .CD(n_62691), .Q(queue
		[183]));
	notech_mux2 i_23838(.S(n_56585), .A(queue[183]), .B(n_17530), .Z(n_16853
		));
	notech_reg queue_reg_184(.CP(n_63564), .D(n_16859), .CD(n_62691), .Q(queue
		[184]));
	notech_mux2 i_23846(.S(n_56585), .A(queue[184]), .B(n_17532), .Z(n_16859
		));
	notech_reg queue_reg_185(.CP(n_63564), .D(n_16865), .CD(n_62691), .Q(queue
		[185]));
	notech_mux2 i_23854(.S(n_56585), .A(queue[185]), .B(n_17534), .Z(n_16865
		));
	notech_reg queue_reg_186(.CP(n_63564), .D(n_16871), .CD(n_62693), .Q(queue
		[186]));
	notech_mux2 i_23862(.S(n_56585), .A(queue[186]), .B(n_17536), .Z(n_16871
		));
	notech_reg queue_reg_187(.CP(n_63564), .D(n_16877), .CD(n_62693), .Q(queue
		[187]));
	notech_mux2 i_23870(.S(n_56585), .A(queue[187]), .B(n_17538), .Z(n_16877
		));
	notech_reg queue_reg_188(.CP(n_63564), .D(n_16883), .CD(n_62693), .Q(queue
		[188]));
	notech_mux2 i_23878(.S(n_56585), .A(queue[188]), .B(n_17540), .Z(n_16883
		));
	notech_reg queue_reg_189(.CP(n_63564), .D(n_16889), .CD(n_62691), .Q(queue
		[189]));
	notech_mux2 i_23886(.S(n_56585), .A(queue[189]), .B(n_17542), .Z(n_16889
		));
	notech_reg queue_reg_190(.CP(n_63564), .D(n_16895), .CD(n_62693), .Q(queue
		[190]));
	notech_mux2 i_23894(.S(n_56585), .A(queue[190]), .B(n_17544), .Z(n_16895
		));
	notech_nand3 i_12034810(.A(n_61409), .B(n_60101), .C(queue[10]), .Z(n_1177
		));
	notech_reg queue_reg_191(.CP(n_63564), .D(n_16901), .CD(n_62694), .Q(queue
		[191]));
	notech_mux2 i_23902(.S(n_56585), .A(queue[191]), .B(n_17546), .Z(n_16901
		));
	notech_reg queue_reg_192(.CP(n_63564), .D(n_16907), .CD(n_62695), .Q(queue
		[192]));
	notech_mux2 i_23910(.S(n_56572), .A(queue[192]), .B(n_17548), .Z(n_16907
		));
	notech_reg queue_reg_193(.CP(n_63564), .D(n_16913), .CD(n_62695), .Q(queue
		[193]));
	notech_mux2 i_23918(.S(n_56572), .A(queue[193]), .B(n_17550), .Z(n_16913
		));
	notech_and4 i_224968(.A(n_2021), .B(n_2020), .C(n_2015), .D(n_2019), .Z(squeue_1101084
		));
	notech_reg queue_reg_194(.CP(n_63564), .D(n_16919), .CD(n_62695), .Q(queue
		[194]));
	notech_mux2 i_23926(.S(n_56572), .A(queue[194]), .B(n_17552), .Z(n_16919
		));
	notech_nand3 i_10234828(.A(n_59657), .B(n_59931), .C(queue[1]), .Z(n_1174
		));
	notech_reg queue_reg_195(.CP(n_63564), .D(n_16925), .CD(n_62694), .Q(queue
		[195]));
	notech_mux2 i_23934(.S(n_56572), .A(queue[195]), .B(n_17554), .Z(n_16925
		));
	notech_reg queue_reg_196(.CP(n_63564), .D(n_16931), .CD(n_62695), .Q(queue
		[196]));
	notech_mux2 i_23942(.S(n_56572), .A(queue[196]), .B(n_17556), .Z(n_16931
		));
	notech_reg queue_reg_197(.CP(n_63564), .D(n_16937), .CD(n_62695), .Q(queue
		[197]));
	notech_mux2 i_23950(.S(n_56572), .A(queue[197]), .B(n_17558), .Z(n_16937
		));
	notech_reg queue_reg_198(.CP(n_63488), .D(n_16943), .CD(n_62695), .Q(queue
		[198]));
	notech_mux2 i_23958(.S(n_56572), .A(queue[198]), .B(n_17560), .Z(n_16943
		));
	notech_reg queue_reg_199(.CP(n_63488), .D(n_16949), .CD(n_62695), .Q(queue
		[199]));
	notech_mux2 i_23966(.S(n_56572), .A(queue[199]), .B(n_17562), .Z(n_16949
		));
	notech_reg queue_reg_200(.CP(n_63488), .D(n_16955), .CD(n_62695), .Q(queue
		[200]));
	notech_mux2 i_23974(.S(n_56572), .A(queue[200]), .B(n_17564), .Z(n_16955
		));
	notech_reg queue_reg_201(.CP(n_63488), .D(n_16961), .CD(n_62695), .Q(queue
		[201]));
	notech_mux2 i_23982(.S(n_56572), .A(queue[201]), .B(n_17566), .Z(n_16961
		));
	notech_reg queue_reg_202(.CP(n_63488), .D(n_16967), .CD(n_62694), .Q(queue
		[202]));
	notech_mux2 i_23990(.S(n_56572), .A(queue[202]), .B(n_17568), .Z(n_16967
		));
	notech_reg queue_reg_203(.CP(n_63488), .D(n_16973), .CD(n_62694), .Q(queue
		[203]));
	notech_mux2 i_23998(.S(n_56572), .A(queue[203]), .B(n_17570), .Z(n_16973
		));
	notech_reg queue_reg_204(.CP(clk), .D(n_16979), .CD(n_62694), .Q(queue[
		204]));
	notech_mux2 i_24006(.S(n_56572), .A(queue[204]), .B(n_17572), .Z(n_16979
		));
	notech_reg queue_reg_205(.CP(n_63486), .D(n_16985), .CD(n_62694), .Q(queue
		[205]));
	notech_mux2 i_24014(.S(n_56572), .A(queue[205]), .B(n_17574), .Z(n_16985
		));
	notech_reg queue_reg_206(.CP(n_63560), .D(n_16991), .CD(n_62694), .Q(queue
		[206]));
	notech_mux2 i_24022(.S(n_56572), .A(queue[206]), .B(n_17576), .Z(n_16991
		));
	notech_reg queue_reg_207(.CP(n_63560), .D(n_16997), .CD(n_62694), .Q(queue
		[207]));
	notech_mux2 i_24030(.S(n_56572), .A(queue[207]), .B(n_17578), .Z(n_16997
		));
	notech_nand3 i_8934841(.A(n_61409), .B(n_60101), .C(queue[9]), .Z(n_1161
		));
	notech_reg queue_reg_208(.CP(n_63560), .D(n_17003), .CD(n_62694), .Q(queue
		[208]));
	notech_mux2 i_24038(.S(n_56570), .A(queue[208]), .B(n_17580), .Z(n_17003
		));
	notech_reg queue_reg_209(.CP(n_63560), .D(n_17009), .CD(n_62694), .Q(queue
		[209]));
	notech_mux2 i_24046(.S(n_56570), .A(queue[209]), .B(n_17582), .Z(n_17009
		));
	notech_reg queue_reg_210(.CP(n_63560), .D(n_17015), .CD(n_62694), .Q(queue
		[210]));
	notech_mux2 i_24054(.S(n_56570), .A(queue[210]), .B(n_17584), .Z(n_17015
		));
	notech_and4 i_124967(.A(n_2007), .B(n_2004), .C(n_1993), .D(n_2001), .Z(squeue_0101085
		));
	notech_reg queue_reg_211(.CP(n_63636), .D(n_17021), .CD(n_62694), .Q(queue
		[211]));
	notech_mux2 i_24062(.S(n_56570), .A(queue[211]), .B(n_17586), .Z(n_17021
		));
	notech_nand3 i_6934859(.A(n_59657), .B(n_59931), .C(queue[0]), .Z(n_1158
		));
	notech_reg queue_reg_212(.CP(n_63636), .D(n_17027), .CD(n_62694), .Q(queue
		[212]));
	notech_mux2 i_24070(.S(n_56570), .A(queue[212]), .B(n_17588), .Z(n_17027
		));
	notech_reg queue_reg_213(.CP(n_63636), .D(n_17033), .CD(n_62689), .Q(queue
		[213]));
	notech_mux2 i_24078(.S(n_56570), .A(queue[213]), .B(n_17590), .Z(n_17033
		));
	notech_reg queue_reg_214(.CP(n_63636), .D(n_17039), .CD(n_62689), .Q(queue
		[214]));
	notech_mux2 i_24086(.S(n_56570), .A(queue[214]), .B(n_17592), .Z(n_17039
		));
	notech_reg queue_reg_215(.CP(n_63636), .D(n_17045), .CD(n_62689), .Q(queue
		[215]));
	notech_mux2 i_24094(.S(n_56570), .A(queue[215]), .B(n_17594), .Z(n_17045
		));
	notech_reg queue_reg_216(.CP(n_63636), .D(n_17051), .CD(n_62689), .Q(queue
		[216]));
	notech_mux2 i_24102(.S(n_56570), .A(queue[216]), .B(n_17596), .Z(n_17051
		));
	notech_reg queue_reg_217(.CP(n_63636), .D(n_17057), .CD(n_62689), .Q(queue
		[217]));
	notech_mux2 i_24110(.S(n_56570), .A(queue[217]), .B(n_17598), .Z(n_17057
		));
	notech_reg queue_reg_218(.CP(n_63636), .D(n_17063), .CD(n_62689), .Q(queue
		[218]));
	notech_mux2 i_24118(.S(n_56570), .A(queue[218]), .B(n_17600), .Z(n_17063
		));
	notech_reg queue_reg_219(.CP(n_63636), .D(n_17069), .CD(n_62689), .Q(queue
		[219]));
	notech_mux2 i_24126(.S(n_56570), .A(queue[219]), .B(n_17602), .Z(n_17069
		));
	notech_reg queue_reg_220(.CP(n_63636), .D(n_17075), .CD(n_62689), .Q(queue
		[220]));
	notech_mux2 i_24134(.S(n_56570), .A(queue[220]), .B(n_17604), .Z(n_17075
		));
	notech_reg queue_reg_221(.CP(n_63636), .D(n_17081), .CD(n_62689), .Q(queue
		[221]));
	notech_mux2 i_24142(.S(n_56570), .A(queue[221]), .B(n_17606), .Z(n_17081
		));
	notech_reg queue_reg_222(.CP(n_63636), .D(n_17087), .CD(n_62689), .Q(queue
		[222]));
	notech_mux2 i_24150(.S(n_56570), .A(queue[222]), .B(n_17608), .Z(n_17087
		));
	notech_reg queue_reg_223(.CP(n_63636), .D(n_17093), .CD(n_62689), .Q(queue
		[223]));
	notech_mux2 i_24158(.S(n_56570), .A(queue[223]), .B(n_17610), .Z(n_17093
		));
	notech_reg queue_reg_224(.CP(n_63636), .D(n_17099), .CD(n_62688), .Q(queue
		[224]));
	notech_mux2 i_24166(.S(n_56577), .A(queue[224]), .B(n_17612), .Z(n_17099
		));
	notech_nand3 i_5434872(.A(n_61409), .B(n_60101), .C(queue[8]), .Z(n_1145
		));
	notech_reg queue_reg_225(.CP(n_63636), .D(n_17105), .CD(n_62688), .Q(queue
		[225]));
	notech_mux2 i_24174(.S(n_56577), .A(queue[225]), .B(n_17614), .Z(n_17105
		));
	notech_reg queue_reg_226(.CP(n_63636), .D(n_17111), .CD(n_62688), .Q(queue
		[226]));
	notech_mux2 i_24182(.S(n_56577), .A(queue[226]), .B(n_17616), .Z(n_17111
		));
	notech_reg queue_reg_227(.CP(n_63636), .D(n_17117), .CD(n_62688), .Q(queue
		[227]));
	notech_mux2 i_24190(.S(n_56577), .A(queue[227]), .B(n_17618), .Z(n_17117
		));
	notech_reg queue_reg_228(.CP(n_63636), .D(n_17123), .CD(n_62688), .Q(queue
		[228]));
	notech_mux2 i_24198(.S(n_56577), .A(queue[228]), .B(n_17620), .Z(n_17123
		));
	notech_reg queue_reg_229(.CP(n_63560), .D(n_17129), .CD(n_62689), .Q(queue
		[229]));
	notech_mux2 i_24206(.S(n_56577), .A(queue[229]), .B(n_17622), .Z(n_17129
		));
	notech_nand3 i_45035023(.A(addrshft[3]), .B(n_17678), .C(n_17679), .Z(n_1137
		));
	notech_reg queue_reg_230(.CP(n_63636), .D(n_17135), .CD(n_62689), .Q(queue
		[230]));
	notech_mux2 i_24214(.S(n_56577), .A(queue[230]), .B(n_17624), .Z(n_17135
		));
	notech_nor2 i_3131131(.A(addrshft[0]), .B(addrshft[1]), .Z(n_1134));
	notech_reg queue_reg_231(.CP(n_63562), .D(n_17141), .CD(n_62689), .Q(queue
		[231]));
	notech_mux2 i_24222(.S(n_56577), .A(queue[231]), .B(n_17626), .Z(n_17141
		));
	notech_or2 i_45135022(.A(addrshft[0]), .B(n_17678), .Z(n_113356519));
	notech_reg queue_reg_232(.CP(n_63562), .D(n_17147), .CD(n_62688), .Q(queue
		[232]));
	notech_mux2 i_24230(.S(n_56577), .A(queue[232]), .B(n_17628), .Z(n_17147
		));
	notech_nand3 i_6135438(.A(wptr[0]), .B(n_3070), .C(n_17301), .Z(n_113256518
		));
	notech_reg queue_reg_233(.CP(n_63562), .D(n_17153), .CD(n_62688), .Q(queue
		[233]));
	notech_mux2 i_24238(.S(n_56577), .A(queue[233]), .B(n_17630), .Z(n_17153
		));
	notech_reg queue_reg_234(.CP(n_63562), .D(n_17159), .CD(n_62690), .Q(queue
		[234]));
	notech_mux2 i_24246(.S(n_56577), .A(queue[234]), .B(n_17632), .Z(n_17159
		));
	notech_reg queue_reg_235(.CP(n_63562), .D(n_17165), .CD(n_62691), .Q(queue
		[235]));
	notech_mux2 i_24254(.S(n_56577), .A(queue[235]), .B(n_17634), .Z(n_17165
		));
	notech_ao4 i_3335435(.A(wptr[0]), .B(n_17301), .C(n_113256518), .D(n_17677
		), .Z(n_1129));
	notech_reg queue_reg_236(.CP(n_63562), .D(n_17171), .CD(n_62691), .Q(queue
		[236]));
	notech_mux2 i_24262(.S(n_56577), .A(queue[236]), .B(n_17636), .Z(n_17171
		));
	notech_reg queue_reg_237(.CP(n_63562), .D(n_17177), .CD(n_62691), .Q(queue
		[237]));
	notech_mux2 i_24270(.S(n_56577), .A(queue[237]), .B(n_17638), .Z(n_17177
		));
	notech_reg queue_reg_238(.CP(n_63562), .D(n_17183), .CD(n_62690), .Q(queue
		[238]));
	notech_mux2 i_24278(.S(n_56577), .A(queue[238]), .B(n_17640), .Z(n_17183
		));
	notech_reg queue_reg_239(.CP(n_63562), .D(n_17189), .CD(n_62690), .Q(queue
		[239]));
	notech_mux2 i_24286(.S(n_56577), .A(queue[239]), .B(n_17642), .Z(n_17189
		));
	notech_reg queue_reg_240(.CP(n_63562), .D(n_17195), .CD(n_62691), .Q(queue
		[240]));
	notech_mux2 i_24294(.S(n_56575), .A(queue[240]), .B(n_17644), .Z(n_17195
		));
	notech_reg queue_reg_241(.CP(n_63562), .D(n_17201), .CD(n_62691), .Q(queue
		[241]));
	notech_mux2 i_24302(.S(n_56575), .A(queue[241]), .B(n_17646), .Z(n_17201
		));
	notech_xor2 i_3735431(.A(n_1134), .B(addrshft[2]), .Z(n_1123));
	notech_reg queue_reg_242(.CP(n_63562), .D(n_17207), .CD(n_62691), .Q(queue
		[242]));
	notech_mux2 i_24310(.S(n_56575), .A(queue[242]), .B(n_17648), .Z(n_17207
		));
	notech_reg queue_reg_243(.CP(n_63562), .D(n_17213), .CD(n_62691), .Q(queue
		[243]));
	notech_mux2 i_24318(.S(n_56575), .A(queue[243]), .B(n_17650), .Z(n_17213
		));
	notech_reg queue_reg_244(.CP(n_63562), .D(n_17219), .CD(n_62691), .Q(queue
		[244]));
	notech_mux2 i_24326(.S(n_56575), .A(queue[244]), .B(n_17652), .Z(n_17219
		));
	notech_reg queue_reg_245(.CP(n_63562), .D(n_17225), .CD(n_62690), .Q(queue
		[245]));
	notech_mux2 i_24334(.S(n_56575), .A(queue[245]), .B(n_17654), .Z(n_17225
		));
	notech_reg queue_reg_246(.CP(n_63562), .D(n_17231), .CD(n_62690), .Q(queue
		[246]));
	notech_mux2 i_24342(.S(n_56575), .A(queue[246]), .B(n_17656), .Z(n_17231
		));
	notech_ao4 i_3835430(.A(n_61409), .B(addrshft[3]), .C(addrshft[0]), .D(n_1137
		), .Z(n_1114));
	notech_reg queue_reg_247(.CP(n_63562), .D(n_17237), .CD(n_62690), .Q(queue
		[247]));
	notech_mux2 i_24350(.S(n_56575), .A(queue[247]), .B(n_17658), .Z(n_17237
		));
	notech_reg queue_reg_248(.CP(n_63562), .D(n_17243), .CD(n_62690), .Q(queue
		[248]));
	notech_mux2 i_24358(.S(n_56575), .A(queue[248]), .B(n_17660), .Z(n_17243
		));
	notech_reg queue_reg_249(.CP(n_63562), .D(n_17249), .CD(n_62690), .Q(queue
		[249]));
	notech_mux2 i_24366(.S(n_56575), .A(queue[249]), .B(n_17662), .Z(n_17249
		));
	notech_reg queue_reg_250(.CP(n_63486), .D(n_17255), .CD(n_62690), .Q(queue
		[250]));
	notech_mux2 i_24374(.S(n_56575), .A(queue[250]), .B(n_17664), .Z(n_17255
		));
	notech_reg queue_reg_251(.CP(n_63486), .D(n_17261), .CD(n_62690), .Q(queue
		[251]));
	notech_mux2 i_24382(.S(n_56575), .A(queue[251]), .B(n_17666), .Z(n_17261
		));
	notech_reg queue_reg_252(.CP(n_63486), .D(n_17267), .CD(n_62690), .Q(queue
		[252]));
	notech_mux2 i_24390(.S(n_56575), .A(queue[252]), .B(n_17668), .Z(n_17267
		));
	notech_reg queue_reg_253(.CP(n_63486), .D(n_17273), .CD(n_62690), .Q(queue
		[253]));
	notech_mux2 i_24398(.S(n_56575), .A(queue[253]), .B(n_17670), .Z(n_17273
		));
	notech_reg queue_reg_254(.CP(clk), .D(n_17279), .CD(n_62690), .Q(queue[
		254]));
	notech_mux2 i_24406(.S(n_56575), .A(queue[254]), .B(n_17672), .Z(n_17279
		));
	notech_reg queue_reg_255(.CP(n_63486), .D(n_17285), .CD(n_62690), .Q(queue
		[255]));
	notech_mux2 i_24414(.S(n_56575), .A(queue[255]), .B(n_17674), .Z(n_17285
		));
	notech_inv i_27467(.A(n_14278717), .Z(n_17291));
	notech_inv i_27468(.A(n_8288), .Z(n_17292));
	notech_inv i_27469(.A(n_8293), .Z(n_17293));
	notech_inv i_27470(.A(n_8291), .Z(n_17294));
	notech_inv i_27472(.A(n_51860125), .Z(n_17296));
	notech_inv i_27473(.A(n_309659577), .Z(n_17297));
	notech_inv i_27474(.A(fault_wptr_en), .Z(n_17298));
	notech_inv i_27475(.A(n_35353), .Z(n_17299));
	notech_inv i_27476(.A(wptr[0]), .Z(n_17300));
	notech_inv i_27477(.A(n_61421), .Z(n_17301));
	notech_inv i_27478(.A(\nbus_12116[0] ), .Z(n_17302));
	notech_inv i_27479(.A(n_34952), .Z(n_17303));
	notech_inv i_27480(.A(n_34958), .Z(n_17304));
	notech_inv i_27481(.A(purge), .Z(cacheD[148]));
	notech_inv i_27482(.A(queue[15]), .Z(n_17306));
	notech_inv i_27483(.A(queue[16]), .Z(n_17307));
	notech_inv i_27484(.A(queue[17]), .Z(n_17308));
	notech_inv i_27485(.A(queue[18]), .Z(n_17309));
	notech_inv i_27486(.A(queue[19]), .Z(n_17310));
	notech_inv i_27487(.A(queue[20]), .Z(n_17311));
	notech_inv i_27488(.A(queue[21]), .Z(n_17312));
	notech_inv i_27489(.A(queue[22]), .Z(n_17313));
	notech_inv i_27490(.A(queue[23]), .Z(n_17314));
	notech_inv i_27491(.A(queue[24]), .Z(n_17315));
	notech_inv i_27492(.A(queue[25]), .Z(n_17316));
	notech_inv i_27493(.A(queue[26]), .Z(n_17317));
	notech_inv i_27494(.A(queue[27]), .Z(n_17318));
	notech_inv i_27495(.A(queue[28]), .Z(n_17319));
	notech_inv i_27496(.A(queue[29]), .Z(n_17320));
	notech_inv i_27497(.A(queue[30]), .Z(n_17321));
	notech_inv i_27498(.A(queue[31]), .Z(n_17322));
	notech_inv i_27499(.A(queue[32]), .Z(n_17323));
	notech_inv i_27500(.A(queue[33]), .Z(n_17324));
	notech_inv i_27501(.A(queue[34]), .Z(n_17325));
	notech_inv i_27502(.A(queue[35]), .Z(n_17326));
	notech_inv i_27503(.A(queue[36]), .Z(n_17327));
	notech_inv i_27504(.A(queue[37]), .Z(n_17328));
	notech_inv i_27505(.A(queue[38]), .Z(n_17329));
	notech_inv i_27506(.A(queue[39]), .Z(n_17330));
	notech_inv i_27507(.A(queue[40]), .Z(n_17331));
	notech_inv i_27508(.A(queue[41]), .Z(n_17332));
	notech_inv i_27509(.A(queue[42]), .Z(n_17333));
	notech_inv i_27510(.A(queue[43]), .Z(n_17334));
	notech_inv i_27511(.A(queue[44]), .Z(n_17335));
	notech_inv i_27512(.A(queue[45]), .Z(n_17336));
	notech_inv i_27513(.A(queue[46]), .Z(n_17337));
	notech_inv i_27514(.A(queue[47]), .Z(n_17338));
	notech_inv i_27515(.A(queue[48]), .Z(n_17339));
	notech_inv i_27516(.A(queue[49]), .Z(n_17340));
	notech_inv i_27517(.A(queue[50]), .Z(n_17341));
	notech_inv i_27518(.A(queue[51]), .Z(n_17342));
	notech_inv i_27519(.A(queue[52]), .Z(n_17343));
	notech_inv i_27520(.A(queue[53]), .Z(n_17344));
	notech_inv i_27521(.A(queue[54]), .Z(n_17345));
	notech_inv i_27522(.A(queue[55]), .Z(n_17346));
	notech_inv i_27523(.A(queue[56]), .Z(n_17347));
	notech_inv i_27524(.A(queue[57]), .Z(n_17348));
	notech_inv i_27525(.A(queue[58]), .Z(n_17349));
	notech_inv i_27526(.A(queue[59]), .Z(n_17350));
	notech_inv i_27527(.A(queue[60]), .Z(n_17351));
	notech_inv i_27528(.A(queue[61]), .Z(n_17352));
	notech_inv i_27529(.A(queue[62]), .Z(n_17353));
	notech_inv i_27530(.A(queue[63]), .Z(n_17354));
	notech_inv i_27531(.A(queue[64]), .Z(n_17355));
	notech_inv i_27532(.A(queue[65]), .Z(n_17356));
	notech_inv i_27533(.A(queue[66]), .Z(n_17357));
	notech_inv i_27534(.A(queue[67]), .Z(n_17358));
	notech_inv i_27535(.A(queue[68]), .Z(n_17359));
	notech_inv i_27536(.A(queue[69]), .Z(n_17360));
	notech_inv i_27537(.A(queue[70]), .Z(n_17361));
	notech_inv i_27538(.A(queue[71]), .Z(n_17362));
	notech_inv i_27539(.A(queue[72]), .Z(n_17363));
	notech_inv i_27540(.A(queue[73]), .Z(n_17364));
	notech_inv i_27541(.A(queue[74]), .Z(n_17365));
	notech_inv i_27542(.A(queue[75]), .Z(n_17366));
	notech_inv i_27543(.A(queue[76]), .Z(n_17367));
	notech_inv i_27544(.A(queue[77]), .Z(n_17368));
	notech_inv i_27545(.A(queue[78]), .Z(n_17369));
	notech_inv i_27546(.A(queue[79]), .Z(n_17370));
	notech_inv i_27547(.A(queue[80]), .Z(n_17371));
	notech_inv i_27548(.A(queue[81]), .Z(n_17372));
	notech_inv i_27549(.A(queue[82]), .Z(n_17373));
	notech_inv i_27550(.A(queue[83]), .Z(n_17374));
	notech_inv i_27551(.A(queue[84]), .Z(n_17375));
	notech_inv i_27552(.A(queue[85]), .Z(n_17376));
	notech_inv i_27553(.A(queue[86]), .Z(n_17377));
	notech_inv i_27554(.A(queue[87]), .Z(n_17378));
	notech_inv i_27555(.A(queue[88]), .Z(n_17379));
	notech_inv i_27556(.A(queue[89]), .Z(n_17380));
	notech_inv i_27557(.A(queue[90]), .Z(n_17381));
	notech_inv i_27558(.A(queue[91]), .Z(n_17382));
	notech_inv i_27559(.A(queue[92]), .Z(n_17383));
	notech_inv i_27560(.A(queue[93]), .Z(n_17384));
	notech_inv i_27561(.A(queue[94]), .Z(n_17385));
	notech_inv i_27562(.A(queue[95]), .Z(n_17386));
	notech_inv i_27563(.A(queue[96]), .Z(n_17387));
	notech_inv i_27564(.A(queue[97]), .Z(n_17388));
	notech_inv i_27565(.A(queue[98]), .Z(n_17389));
	notech_inv i_27566(.A(queue[99]), .Z(n_17390));
	notech_inv i_27567(.A(queue[100]), .Z(n_17391));
	notech_inv i_27568(.A(queue[101]), .Z(n_17392));
	notech_inv i_27569(.A(queue[102]), .Z(n_17393));
	notech_inv i_27570(.A(queue[103]), .Z(n_17394));
	notech_inv i_27571(.A(queue[104]), .Z(n_17395));
	notech_inv i_27572(.A(queue[105]), .Z(n_17396));
	notech_inv i_27573(.A(queue[106]), .Z(n_17397));
	notech_inv i_27574(.A(queue[107]), .Z(n_17398));
	notech_inv i_27575(.A(queue[108]), .Z(n_17399));
	notech_inv i_27576(.A(queue[109]), .Z(n_17400));
	notech_inv i_27577(.A(queue[110]), .Z(n_17401));
	notech_inv i_27578(.A(queue[111]), .Z(n_17402));
	notech_inv i_27579(.A(queue[112]), .Z(n_17403));
	notech_inv i_27580(.A(queue[113]), .Z(n_17404));
	notech_inv i_27581(.A(queue[114]), .Z(n_17405));
	notech_inv i_27582(.A(queue[115]), .Z(n_17406));
	notech_inv i_27583(.A(queue[116]), .Z(n_17407));
	notech_inv i_27584(.A(queue[117]), .Z(n_17408));
	notech_inv i_27585(.A(queue[118]), .Z(n_17409));
	notech_inv i_27586(.A(queue[119]), .Z(n_17410));
	notech_inv i_27587(.A(queue[120]), .Z(n_17411));
	notech_inv i_27588(.A(queue[121]), .Z(n_17412));
	notech_inv i_27589(.A(queue[122]), .Z(n_17413));
	notech_inv i_27590(.A(queue[123]), .Z(n_17414));
	notech_inv i_27591(.A(queue[124]), .Z(n_17415));
	notech_inv i_27592(.A(queue[125]), .Z(n_17416));
	notech_inv i_27593(.A(queue[126]), .Z(n_17417));
	notech_inv i_27594(.A(queue[127]), .Z(n_17418));
	notech_inv i_27596(.A(n_36149), .Z(n_17420));
	notech_inv i_27597(.A(queue[128]), .Z(n_17421));
	notech_inv i_27598(.A(n_36155), .Z(n_17422));
	notech_inv i_27599(.A(queue[129]), .Z(n_17423));
	notech_inv i_27600(.A(n_36161), .Z(n_17424));
	notech_inv i_27601(.A(queue[130]), .Z(n_17425));
	notech_inv i_27602(.A(n_36167), .Z(n_17426));
	notech_inv i_27603(.A(queue[131]), .Z(n_17427));
	notech_inv i_27604(.A(n_36173), .Z(n_17428));
	notech_inv i_27605(.A(queue[132]), .Z(n_17429));
	notech_inv i_27606(.A(n_36179), .Z(n_17430));
	notech_inv i_27607(.A(queue[133]), .Z(n_17431));
	notech_inv i_27608(.A(n_36185), .Z(n_17432));
	notech_inv i_27609(.A(queue[134]), .Z(n_17433));
	notech_inv i_27610(.A(n_36191), .Z(n_17434));
	notech_inv i_27611(.A(queue[135]), .Z(n_17435));
	notech_inv i_27612(.A(n_36197), .Z(n_17436));
	notech_inv i_27613(.A(queue[136]), .Z(n_17437));
	notech_inv i_27614(.A(n_36203), .Z(n_17438));
	notech_inv i_27615(.A(queue[137]), .Z(n_17439));
	notech_inv i_27616(.A(n_36209), .Z(n_17440));
	notech_inv i_27617(.A(queue[138]), .Z(n_17441));
	notech_inv i_27618(.A(n_36215), .Z(n_17442));
	notech_inv i_27619(.A(queue[139]), .Z(n_17443));
	notech_inv i_27620(.A(n_36221), .Z(n_17444));
	notech_inv i_27621(.A(queue[140]), .Z(n_17445));
	notech_inv i_27622(.A(n_36227), .Z(n_17446));
	notech_inv i_27623(.A(queue[141]), .Z(n_17447));
	notech_inv i_27624(.A(n_36233), .Z(n_17448));
	notech_inv i_27625(.A(queue[142]), .Z(n_17449));
	notech_inv i_27626(.A(n_36239), .Z(n_17450));
	notech_inv i_27627(.A(queue[143]), .Z(n_17451));
	notech_inv i_27628(.A(n_36245), .Z(n_17452));
	notech_inv i_27629(.A(queue[144]), .Z(n_17453));
	notech_inv i_27630(.A(n_36251), .Z(n_17454));
	notech_inv i_27631(.A(queue[145]), .Z(n_17455));
	notech_inv i_27632(.A(n_36257), .Z(n_17456));
	notech_inv i_27633(.A(queue[146]), .Z(n_17457));
	notech_inv i_27634(.A(n_36263), .Z(n_17458));
	notech_inv i_27635(.A(queue[147]), .Z(n_17459));
	notech_inv i_27636(.A(n_36269), .Z(n_17460));
	notech_inv i_27637(.A(queue[148]), .Z(n_17461));
	notech_inv i_27638(.A(n_36275), .Z(n_17462));
	notech_inv i_27639(.A(queue[149]), .Z(n_17463));
	notech_inv i_27640(.A(n_36281), .Z(n_17464));
	notech_inv i_27641(.A(queue[150]), .Z(n_17465));
	notech_inv i_27642(.A(n_36287), .Z(n_17466));
	notech_inv i_27643(.A(queue[151]), .Z(n_17467));
	notech_inv i_27644(.A(n_36293), .Z(n_17468));
	notech_inv i_27645(.A(queue[152]), .Z(n_17469));
	notech_inv i_27646(.A(n_36299), .Z(n_17470));
	notech_inv i_27647(.A(queue[153]), .Z(n_17471));
	notech_inv i_27648(.A(n_36305), .Z(n_17472));
	notech_inv i_27649(.A(queue[154]), .Z(n_17473));
	notech_inv i_27650(.A(n_36311), .Z(n_17474));
	notech_inv i_27651(.A(queue[155]), .Z(n_17475));
	notech_inv i_27652(.A(n_36317), .Z(n_17476));
	notech_inv i_27653(.A(queue[156]), .Z(n_17477));
	notech_inv i_27654(.A(n_36323), .Z(n_17478));
	notech_inv i_27655(.A(queue[157]), .Z(n_17479));
	notech_inv i_27656(.A(n_36329), .Z(n_17480));
	notech_inv i_27657(.A(queue[158]), .Z(n_17481));
	notech_inv i_27658(.A(n_36335), .Z(n_17482));
	notech_inv i_27659(.A(queue[159]), .Z(n_17483));
	notech_inv i_27660(.A(n_36341), .Z(n_17484));
	notech_inv i_27661(.A(queue[160]), .Z(n_17485));
	notech_inv i_27662(.A(n_36347), .Z(n_17486));
	notech_inv i_27663(.A(queue[161]), .Z(n_17487));
	notech_inv i_27664(.A(n_36353), .Z(n_17488));
	notech_inv i_27665(.A(queue[162]), .Z(n_17489));
	notech_inv i_27666(.A(n_36359), .Z(n_17490));
	notech_inv i_27667(.A(queue[163]), .Z(n_17491));
	notech_inv i_27668(.A(n_36365), .Z(n_17492));
	notech_inv i_27669(.A(queue[164]), .Z(n_17493));
	notech_inv i_27670(.A(n_36371), .Z(n_17494));
	notech_inv i_27671(.A(queue[165]), .Z(n_17495));
	notech_inv i_27672(.A(n_36377), .Z(n_17496));
	notech_inv i_27673(.A(queue[166]), .Z(n_17497));
	notech_inv i_27674(.A(n_36383), .Z(n_17498));
	notech_inv i_27675(.A(queue[167]), .Z(n_17499));
	notech_inv i_27676(.A(n_36389), .Z(n_17500));
	notech_inv i_27677(.A(queue[168]), .Z(n_17501));
	notech_inv i_27678(.A(n_36395), .Z(n_17502));
	notech_inv i_27679(.A(queue[169]), .Z(n_17503));
	notech_inv i_27680(.A(n_36401), .Z(n_17504));
	notech_inv i_27681(.A(queue[170]), .Z(n_17505));
	notech_inv i_27682(.A(n_36407), .Z(n_17506));
	notech_inv i_27683(.A(queue[171]), .Z(n_17507));
	notech_inv i_27684(.A(n_36413), .Z(n_17508));
	notech_inv i_27685(.A(queue[172]), .Z(n_17509));
	notech_inv i_27686(.A(n_36419), .Z(n_17510));
	notech_inv i_27687(.A(queue[173]), .Z(n_17511));
	notech_inv i_27688(.A(n_36425), .Z(n_17512));
	notech_inv i_27689(.A(queue[174]), .Z(n_17513));
	notech_inv i_27690(.A(n_36431), .Z(n_17514));
	notech_inv i_27691(.A(queue[175]), .Z(n_17515));
	notech_inv i_27692(.A(n_36437), .Z(n_17516));
	notech_inv i_27693(.A(queue[176]), .Z(n_17517));
	notech_inv i_27694(.A(n_36443), .Z(n_17518));
	notech_inv i_27695(.A(queue[177]), .Z(n_17519));
	notech_inv i_27696(.A(n_36449), .Z(n_17520));
	notech_inv i_27697(.A(queue[178]), .Z(n_17521));
	notech_inv i_27698(.A(n_36455), .Z(n_17522));
	notech_inv i_27699(.A(queue[179]), .Z(n_17523));
	notech_inv i_27700(.A(n_36461), .Z(n_17524));
	notech_inv i_27701(.A(queue[180]), .Z(n_17525));
	notech_inv i_27702(.A(n_36467), .Z(n_17526));
	notech_inv i_27703(.A(queue[181]), .Z(n_17527));
	notech_inv i_27704(.A(n_36473), .Z(n_17528));
	notech_inv i_27705(.A(queue[182]), .Z(n_17529));
	notech_inv i_27706(.A(n_36479), .Z(n_17530));
	notech_inv i_27707(.A(queue[183]), .Z(n_17531));
	notech_inv i_27708(.A(n_36485), .Z(n_17532));
	notech_inv i_27709(.A(queue[184]), .Z(n_17533));
	notech_inv i_27710(.A(n_36491), .Z(n_17534));
	notech_inv i_27711(.A(queue[185]), .Z(n_17535));
	notech_inv i_27712(.A(n_36497), .Z(n_17536));
	notech_inv i_27713(.A(queue[186]), .Z(n_17537));
	notech_inv i_27714(.A(n_36503), .Z(n_17538));
	notech_inv i_27715(.A(queue[187]), .Z(n_17539));
	notech_inv i_27716(.A(n_36509), .Z(n_17540));
	notech_inv i_27717(.A(queue[188]), .Z(n_17541));
	notech_inv i_27718(.A(n_36515), .Z(n_17542));
	notech_inv i_27719(.A(queue[189]), .Z(n_17543));
	notech_inv i_27720(.A(n_36521), .Z(n_17544));
	notech_inv i_27721(.A(queue[190]), .Z(n_17545));
	notech_inv i_27722(.A(n_36527), .Z(n_17546));
	notech_inv i_27723(.A(queue[191]), .Z(n_17547));
	notech_inv i_27724(.A(n_36533), .Z(n_17548));
	notech_inv i_27725(.A(queue[192]), .Z(n_17549));
	notech_inv i_27726(.A(n_36539), .Z(n_17550));
	notech_inv i_27727(.A(queue[193]), .Z(n_17551));
	notech_inv i_27728(.A(n_36545), .Z(n_17552));
	notech_inv i_27729(.A(queue[194]), .Z(n_17553));
	notech_inv i_27730(.A(n_36551), .Z(n_17554));
	notech_inv i_27731(.A(queue[195]), .Z(n_17555));
	notech_inv i_27732(.A(n_36557), .Z(n_17556));
	notech_inv i_27733(.A(queue[196]), .Z(n_17557));
	notech_inv i_27734(.A(n_36563), .Z(n_17558));
	notech_inv i_27735(.A(queue[197]), .Z(n_17559));
	notech_inv i_27736(.A(n_36569), .Z(n_17560));
	notech_inv i_27737(.A(queue[198]), .Z(n_17561));
	notech_inv i_27738(.A(n_36575), .Z(n_17562));
	notech_inv i_27739(.A(queue[199]), .Z(n_17563));
	notech_inv i_27740(.A(n_36581), .Z(n_17564));
	notech_inv i_27741(.A(queue[200]), .Z(n_17565));
	notech_inv i_27742(.A(n_36587), .Z(n_17566));
	notech_inv i_27743(.A(queue[201]), .Z(n_17567));
	notech_inv i_27744(.A(n_36593), .Z(n_17568));
	notech_inv i_27745(.A(queue[202]), .Z(n_17569));
	notech_inv i_27746(.A(n_36599), .Z(n_17570));
	notech_inv i_27747(.A(queue[203]), .Z(n_17571));
	notech_inv i_27748(.A(n_36605), .Z(n_17572));
	notech_inv i_27749(.A(queue[204]), .Z(n_17573));
	notech_inv i_27750(.A(n_36611), .Z(n_17574));
	notech_inv i_27751(.A(queue[205]), .Z(n_17575));
	notech_inv i_27752(.A(n_36617), .Z(n_17576));
	notech_inv i_27753(.A(queue[206]), .Z(n_17577));
	notech_inv i_27754(.A(n_36623), .Z(n_17578));
	notech_inv i_27755(.A(queue[207]), .Z(n_17579));
	notech_inv i_27756(.A(n_36629), .Z(n_17580));
	notech_inv i_27757(.A(queue[208]), .Z(n_17581));
	notech_inv i_27758(.A(n_36635), .Z(n_17582));
	notech_inv i_27759(.A(queue[209]), .Z(n_17583));
	notech_inv i_27760(.A(n_36641), .Z(n_17584));
	notech_inv i_27761(.A(queue[210]), .Z(n_17585));
	notech_inv i_27762(.A(n_36647), .Z(n_17586));
	notech_inv i_27763(.A(queue[211]), .Z(n_17587));
	notech_inv i_27764(.A(n_36653), .Z(n_17588));
	notech_inv i_27765(.A(queue[212]), .Z(n_17589));
	notech_inv i_27766(.A(n_36659), .Z(n_17590));
	notech_inv i_27767(.A(queue[213]), .Z(n_17591));
	notech_inv i_27768(.A(n_36665), .Z(n_17592));
	notech_inv i_27769(.A(queue[214]), .Z(n_17593));
	notech_inv i_27770(.A(n_36671), .Z(n_17594));
	notech_inv i_27771(.A(queue[215]), .Z(n_17595));
	notech_inv i_27772(.A(n_36677), .Z(n_17596));
	notech_inv i_27773(.A(queue[216]), .Z(n_17597));
	notech_inv i_27774(.A(n_36683), .Z(n_17598));
	notech_inv i_27775(.A(queue[217]), .Z(n_17599));
	notech_inv i_27776(.A(n_36689), .Z(n_17600));
	notech_inv i_27777(.A(queue[218]), .Z(n_17601));
	notech_inv i_27778(.A(n_36695), .Z(n_17602));
	notech_inv i_27779(.A(queue[219]), .Z(n_17603));
	notech_inv i_27780(.A(n_36701), .Z(n_17604));
	notech_inv i_27781(.A(queue[220]), .Z(n_17605));
	notech_inv i_27782(.A(n_36707), .Z(n_17606));
	notech_inv i_27783(.A(queue[221]), .Z(n_17607));
	notech_inv i_27784(.A(n_36713), .Z(n_17608));
	notech_inv i_27785(.A(queue[222]), .Z(n_17609));
	notech_inv i_27786(.A(n_36719), .Z(n_17610));
	notech_inv i_27787(.A(queue[223]), .Z(n_17611));
	notech_inv i_27788(.A(n_36725), .Z(n_17612));
	notech_inv i_27789(.A(queue[224]), .Z(n_17613));
	notech_inv i_27790(.A(n_36731), .Z(n_17614));
	notech_inv i_27791(.A(queue[225]), .Z(n_17615));
	notech_inv i_27792(.A(n_36737), .Z(n_17616));
	notech_inv i_27793(.A(queue[226]), .Z(n_17617));
	notech_inv i_27794(.A(n_36743), .Z(n_17618));
	notech_inv i_27795(.A(queue[227]), .Z(n_17619));
	notech_inv i_27796(.A(n_36749), .Z(n_17620));
	notech_inv i_27797(.A(queue[228]), .Z(n_17621));
	notech_inv i_27798(.A(n_36755), .Z(n_17622));
	notech_inv i_27799(.A(queue[229]), .Z(n_17623));
	notech_inv i_27800(.A(n_36761), .Z(n_17624));
	notech_inv i_27801(.A(queue[230]), .Z(n_17625));
	notech_inv i_27802(.A(n_36767), .Z(n_17626));
	notech_inv i_27803(.A(queue[231]), .Z(n_17627));
	notech_inv i_27804(.A(n_36773), .Z(n_17628));
	notech_inv i_27805(.A(queue[232]), .Z(n_17629));
	notech_inv i_27806(.A(n_36779), .Z(n_17630));
	notech_inv i_27807(.A(queue[233]), .Z(n_17631));
	notech_inv i_27808(.A(n_36785), .Z(n_17632));
	notech_inv i_27809(.A(queue[234]), .Z(n_17633));
	notech_inv i_27810(.A(n_36791), .Z(n_17634));
	notech_inv i_27811(.A(queue[235]), .Z(n_17635));
	notech_inv i_27812(.A(n_36797), .Z(n_17636));
	notech_inv i_27813(.A(queue[236]), .Z(n_17637));
	notech_inv i_27814(.A(n_36803), .Z(n_17638));
	notech_inv i_27815(.A(queue[237]), .Z(n_17639));
	notech_inv i_27816(.A(n_36809), .Z(n_17640));
	notech_inv i_27817(.A(queue[238]), .Z(n_17641));
	notech_inv i_27818(.A(n_36815), .Z(n_17642));
	notech_inv i_27819(.A(queue[239]), .Z(n_17643));
	notech_inv i_27820(.A(n_36821), .Z(n_17644));
	notech_inv i_27821(.A(queue[240]), .Z(n_17645));
	notech_inv i_27822(.A(n_36827), .Z(n_17646));
	notech_inv i_27823(.A(queue[241]), .Z(n_17647));
	notech_inv i_27824(.A(n_36833), .Z(n_17648));
	notech_inv i_27825(.A(queue[242]), .Z(n_17649));
	notech_inv i_27826(.A(n_36839), .Z(n_17650));
	notech_inv i_27827(.A(queue[243]), .Z(n_17651));
	notech_inv i_27828(.A(n_36845), .Z(n_17652));
	notech_inv i_27829(.A(queue[244]), .Z(n_17653));
	notech_inv i_27830(.A(n_36851), .Z(n_17654));
	notech_inv i_27831(.A(queue[245]), .Z(n_17655));
	notech_inv i_27832(.A(n_36857), .Z(n_17656));
	notech_inv i_27833(.A(queue[246]), .Z(n_17657));
	notech_inv i_27834(.A(n_36863), .Z(n_17658));
	notech_inv i_27835(.A(queue[247]), .Z(n_17659));
	notech_inv i_27836(.A(n_36869), .Z(n_17660));
	notech_inv i_27837(.A(queue[248]), .Z(n_17661));
	notech_inv i_27838(.A(n_36875), .Z(n_17662));
	notech_inv i_27839(.A(queue[249]), .Z(n_17663));
	notech_inv i_27840(.A(n_36881), .Z(n_17664));
	notech_inv i_27841(.A(queue[250]), .Z(n_17665));
	notech_inv i_27842(.A(n_36887), .Z(n_17666));
	notech_inv i_27843(.A(queue[251]), .Z(n_17667));
	notech_inv i_27844(.A(n_36893), .Z(n_17668));
	notech_inv i_27845(.A(queue[252]), .Z(n_17669));
	notech_inv i_27846(.A(n_36899), .Z(n_17670));
	notech_inv i_27847(.A(queue[253]), .Z(n_17671));
	notech_inv i_27848(.A(n_36905), .Z(n_17672));
	notech_inv i_27849(.A(queue[254]), .Z(n_17673));
	notech_inv i_27850(.A(n_36911), .Z(n_17674));
	notech_inv i_27851(.A(queue[255]), .Z(n_17675));
	notech_inv i_27853(.A(addrshft[0]), .Z(n_17677));
	notech_inv i_27854(.A(addrshft[1]), .Z(n_17678));
	notech_inv i_27855(.A(addrshft[2]), .Z(n_17679));
	notech_inv i_27856(.A(tagV[0]), .Z(n_17680));
	notech_inv i_27857(.A(tagV[3]), .Z(n_17681));
	notech_inv i_27858(.A(squeue_0101085), .Z(squeue[0]));
	notech_inv i_27859(.A(squeue_1101084), .Z(squeue[1]));
	notech_inv i_27860(.A(squeue_2101083), .Z(squeue[2]));
	notech_inv i_27861(.A(squeue_3101082), .Z(squeue[3]));
	notech_inv i_27862(.A(squeue_4101081), .Z(squeue[4]));
	notech_inv i_27863(.A(squeue_5101080), .Z(squeue[5]));
	notech_inv i_27864(.A(squeue_6101079), .Z(squeue[6]));
	notech_inv i_27865(.A(squeue_8101078), .Z(squeue[8]));
	notech_inv i_27866(.A(squeue_9101077), .Z(squeue[9]));
	notech_inv i_27867(.A(squeue_10101076), .Z(squeue[10]));
	notech_inv i_27868(.A(squeue_11101075), .Z(squeue[11]));
	notech_inv i_27869(.A(squeue_12101074), .Z(squeue[12]));
	notech_inv i_27870(.A(squeue_13101073), .Z(squeue[13]));
	notech_inv i_27871(.A(squeue_15101072), .Z(squeue[15]));
	notech_inv i_27872(.A(squeue_16101071), .Z(squeue[16]));
	notech_inv i_27873(.A(squeue_17101070), .Z(squeue[17]));
	notech_inv i_27874(.A(squeue_18101069), .Z(squeue[18]));
	notech_inv i_27875(.A(squeue_19101068), .Z(squeue[19]));
	notech_inv i_27876(.A(squeue_20101067), .Z(squeue[20]));
	notech_inv i_27877(.A(squeue_21101066), .Z(squeue[21]));
	notech_inv i_27878(.A(squeue_22101065), .Z(squeue[22]));
	notech_inv i_27879(.A(squeue_23101064), .Z(squeue[23]));
	notech_inv i_27880(.A(squeue_24101063), .Z(squeue[24]));
	notech_inv i_27881(.A(squeue_25101062), .Z(squeue[25]));
	notech_inv i_27882(.A(squeue_26101061), .Z(squeue[26]));
	notech_inv i_27883(.A(squeue_27101060), .Z(squeue[27]));
	notech_inv i_27884(.A(squeue_28101059), .Z(squeue[28]));
	notech_inv i_27885(.A(squeue_30101058), .Z(squeue[30]));
	notech_inv i_27886(.A(squeue_31101057), .Z(squeue[31]));
	notech_inv i_27887(.A(squeue_32101056), .Z(squeue[32]));
	notech_inv i_27888(.A(squeue_33101055), .Z(squeue[33]));
	notech_inv i_27889(.A(squeue_34101054), .Z(squeue[34]));
	notech_inv i_27890(.A(squeue_35101053), .Z(squeue[35]));
	notech_inv i_27891(.A(squeue_36101052), .Z(squeue[36]));
	notech_inv i_27892(.A(squeue_38101051), .Z(squeue[38]));
	notech_inv i_27893(.A(squeue_39101050), .Z(squeue[39]));
	notech_inv i_27894(.A(squeue_40101049), .Z(squeue[40]));
	notech_inv i_27895(.A(squeue_41101048), .Z(squeue[41]));
	notech_inv i_27896(.A(squeue_42101047), .Z(squeue[42]));
	notech_inv i_27897(.A(squeue_43101046), .Z(squeue[43]));
	notech_inv i_27898(.A(squeue_44101045), .Z(squeue[44]));
	notech_inv i_27899(.A(squeue_45101044), .Z(squeue[45]));
	notech_inv i_27900(.A(squeue_46101043), .Z(squeue[46]));
	notech_inv i_27901(.A(squeue_47101042), .Z(squeue[47]));
	notech_inv i_27902(.A(squeue_48101041), .Z(squeue[48]));
	notech_inv i_27903(.A(squeue_49101040), .Z(squeue[49]));
	notech_inv i_27904(.A(squeue_50101039), .Z(squeue[50]));
	notech_inv i_27905(.A(squeue_51101038), .Z(squeue[51]));
	notech_inv i_27906(.A(squeue_52101037), .Z(squeue[52]));
	notech_inv i_27907(.A(squeue_53101036), .Z(squeue[53]));
	notech_inv i_27908(.A(squeue_65101035), .Z(squeue[65]));
	notech_inv i_27909(.A(idata[0]), .Z(n_17733));
	notech_inv i_27910(.A(idata[1]), .Z(n_17734));
	notech_inv i_27911(.A(idata[2]), .Z(n_17735));
	notech_inv i_27912(.A(idata[3]), .Z(n_17736));
	notech_inv i_27913(.A(idata[4]), .Z(n_17737));
	notech_inv i_27914(.A(idata[5]), .Z(n_17738));
	notech_inv i_27915(.A(idata[6]), .Z(n_17739));
	notech_inv i_27916(.A(idata[7]), .Z(n_17740));
	notech_inv i_27917(.A(idata[8]), .Z(n_17741));
	notech_inv i_27918(.A(idata[9]), .Z(n_17742));
	notech_inv i_27919(.A(idata[10]), .Z(n_17743));
	notech_inv i_27920(.A(idata[11]), .Z(n_17744));
	notech_inv i_27921(.A(idata[12]), .Z(n_17745));
	notech_inv i_27922(.A(idata[13]), .Z(n_17746));
	notech_inv i_27923(.A(idata[14]), .Z(n_17747));
	notech_inv i_27924(.A(idata[15]), .Z(n_17748));
	notech_inv i_27925(.A(idata[16]), .Z(n_17749));
	notech_inv i_27926(.A(idata[17]), .Z(n_17750));
	notech_inv i_27927(.A(idata[18]), .Z(n_17751));
	notech_inv i_27928(.A(idata[19]), .Z(n_17752));
	notech_inv i_27929(.A(idata[20]), .Z(n_17753));
	notech_inv i_27930(.A(idata[21]), .Z(n_17754));
	notech_inv i_27931(.A(idata[22]), .Z(n_17755));
	notech_inv i_27932(.A(idata[23]), .Z(n_17756));
	notech_inv i_27933(.A(idata[24]), .Z(n_17757));
	notech_inv i_27934(.A(idata[25]), .Z(n_17758));
	notech_inv i_27935(.A(idata[26]), .Z(n_17759));
	notech_inv i_27936(.A(idata[27]), .Z(n_17760));
	notech_inv i_27937(.A(idata[28]), .Z(n_17761));
	notech_inv i_27938(.A(idata[29]), .Z(n_17762));
	notech_inv i_27939(.A(idata[30]), .Z(n_17763));
	notech_inv i_27940(.A(idata[31]), .Z(n_17764));
	notech_inv i_27941(.A(idata[32]), .Z(n_17765));
	notech_inv i_27942(.A(idata[33]), .Z(n_17766));
	notech_inv i_27943(.A(idata[34]), .Z(n_17767));
	notech_inv i_27944(.A(idata[35]), .Z(n_17768));
	notech_inv i_27945(.A(idata[36]), .Z(n_17769));
	notech_inv i_27946(.A(idata[37]), .Z(n_17770));
	notech_inv i_27947(.A(idata[38]), .Z(n_17771));
	notech_inv i_27948(.A(idata[39]), .Z(n_17772));
	notech_inv i_27949(.A(idata[40]), .Z(n_17773));
	notech_inv i_27950(.A(idata[41]), .Z(n_17774));
	notech_inv i_27951(.A(idata[42]), .Z(n_17775));
	notech_inv i_27952(.A(idata[43]), .Z(n_17776));
	notech_inv i_27953(.A(idata[44]), .Z(n_17777));
	notech_inv i_27954(.A(idata[45]), .Z(n_17778));
	notech_inv i_27955(.A(idata[46]), .Z(n_17779));
	notech_inv i_27956(.A(idata[47]), .Z(n_17780));
	notech_inv i_27957(.A(idata[48]), .Z(n_17781));
	notech_inv i_27958(.A(idata[49]), .Z(n_17782));
	notech_inv i_27959(.A(idata[50]), .Z(n_17783));
	notech_inv i_27960(.A(idata[51]), .Z(n_17784));
	notech_inv i_27961(.A(idata[52]), .Z(n_17785));
	notech_inv i_27962(.A(idata[53]), .Z(n_17786));
	notech_inv i_27963(.A(idata[54]), .Z(n_17787));
	notech_inv i_27964(.A(idata[55]), .Z(n_17788));
	notech_inv i_27965(.A(idata[56]), .Z(n_17789));
	notech_inv i_27966(.A(idata[57]), .Z(n_17790));
	notech_inv i_27967(.A(idata[58]), .Z(n_17791));
	notech_inv i_27968(.A(idata[59]), .Z(n_17792));
	notech_inv i_27969(.A(idata[60]), .Z(n_17793));
	notech_inv i_27970(.A(idata[61]), .Z(n_17794));
	notech_inv i_27971(.A(idata[62]), .Z(n_17795));
	notech_inv i_27972(.A(idata[63]), .Z(n_17796));
	notech_inv i_27973(.A(idata[64]), .Z(n_17797));
	notech_inv i_27974(.A(idata[65]), .Z(n_17798));
	notech_inv i_27975(.A(idata[66]), .Z(n_17799));
	notech_inv i_27976(.A(idata[67]), .Z(n_17800));
	notech_inv i_27977(.A(idata[68]), .Z(n_17801));
	notech_inv i_27978(.A(idata[69]), .Z(n_17802));
	notech_inv i_27979(.A(idata[70]), .Z(n_17803));
	notech_inv i_27980(.A(idata[71]), .Z(n_17804));
	notech_inv i_27981(.A(idata[72]), .Z(n_17805));
	notech_inv i_27982(.A(idata[73]), .Z(n_17806));
	notech_inv i_27983(.A(idata[74]), .Z(n_17807));
	notech_inv i_27984(.A(idata[75]), .Z(n_17808));
	notech_inv i_27985(.A(idata[76]), .Z(n_17809));
	notech_inv i_27986(.A(idata[77]), .Z(n_17810));
	notech_inv i_27987(.A(idata[78]), .Z(n_17811));
	notech_inv i_27988(.A(idata[79]), .Z(n_17812));
	notech_inv i_27989(.A(idata[80]), .Z(n_17813));
	notech_inv i_27990(.A(idata[81]), .Z(n_17814));
	notech_inv i_27991(.A(idata[82]), .Z(n_17815));
	notech_inv i_27992(.A(idata[83]), .Z(n_17816));
	notech_inv i_27993(.A(idata[84]), .Z(n_17817));
	notech_inv i_27994(.A(idata[85]), .Z(n_17818));
	notech_inv i_27995(.A(idata[86]), .Z(n_17819));
	notech_inv i_27996(.A(idata[87]), .Z(n_17820));
	notech_inv i_27997(.A(idata[88]), .Z(n_17821));
	notech_inv i_27998(.A(idata[89]), .Z(n_17822));
	notech_inv i_27999(.A(idata[90]), .Z(n_17823));
	notech_inv i_28000(.A(idata[91]), .Z(n_17824));
	notech_inv i_28001(.A(idata[92]), .Z(n_17825));
	notech_inv i_28002(.A(idata[93]), .Z(n_17826));
	notech_inv i_28003(.A(idata[94]), .Z(n_17827));
	notech_inv i_28004(.A(idata[95]), .Z(n_17828));
	notech_inv i_28005(.A(idata[96]), .Z(n_17829));
	notech_inv i_28006(.A(idata[97]), .Z(n_17830));
	notech_inv i_28007(.A(idata[98]), .Z(n_17831));
	notech_inv i_28008(.A(idata[99]), .Z(n_17832));
	notech_inv i_28009(.A(idata[100]), .Z(n_17833));
	notech_inv i_28010(.A(idata[101]), .Z(n_17834));
	notech_inv i_28011(.A(idata[102]), .Z(n_17835));
	notech_inv i_28012(.A(idata[103]), .Z(n_17836));
	notech_inv i_28013(.A(idata[104]), .Z(n_17837));
	notech_inv i_28014(.A(idata[105]), .Z(n_17838));
	notech_inv i_28015(.A(idata[106]), .Z(n_17839));
	notech_inv i_28016(.A(idata[107]), .Z(n_17840));
	notech_inv i_28017(.A(idata[108]), .Z(n_17841));
	notech_inv i_28018(.A(idata[109]), .Z(n_17842));
	notech_inv i_28019(.A(idata[110]), .Z(n_17843));
	notech_inv i_28020(.A(idata[111]), .Z(n_17844));
	notech_inv i_28021(.A(idata[112]), .Z(n_17845));
	notech_inv i_28022(.A(idata[113]), .Z(n_17846));
	notech_inv i_28023(.A(idata[114]), .Z(n_17847));
	notech_inv i_28024(.A(idata[115]), .Z(n_17848));
	notech_inv i_28025(.A(idata[116]), .Z(n_17849));
	notech_inv i_28026(.A(idata[117]), .Z(n_17850));
	notech_inv i_28027(.A(idata[118]), .Z(n_17851));
	notech_inv i_28028(.A(idata[119]), .Z(n_17852));
	notech_inv i_28029(.A(idata[120]), .Z(n_17853));
	notech_inv i_28030(.A(idata[121]), .Z(n_17854));
	notech_inv i_28031(.A(idata[122]), .Z(n_17855));
	notech_inv i_28032(.A(idata[123]), .Z(n_17856));
	notech_inv i_28033(.A(idata[124]), .Z(n_17857));
	notech_inv i_28034(.A(idata[125]), .Z(n_17858));
	notech_inv i_28035(.A(idata[126]), .Z(n_17859));
	notech_inv i_28036(.A(idata[127]), .Z(n_17860));
	notech_inv i_28037(.A(nbus_12105[4]), .Z(n_17861));
	notech_inv i_28038(.A(nbus_12105[5]), .Z(n_17862));
	notech_inv i_28039(.A(valid_len_0101031), .Z(valid_len[0]));
	notech_inv i_28040(.A(valid_len_1101034), .Z(valid_len[1]));
	notech_inv i_28041(.A(valid_len_2101033), .Z(valid_len[2]));
	notech_inv i_28042(.A(valid_len_3101032), .Z(valid_len[3]));
	notech_inv i_28043(.A(valid_len_4101030), .Z(valid_len[4]));
	notech_inv i_28044(.A(\queue_0[27] ), .Z(n_17868));
	notech_inv i_28045(.A(\queue_0[19] ), .Z(n_17869));
	notech_inv i_28046(.A(\queue_0[11] ), .Z(n_17870));
	notech_inv i_28047(.A(\queue_0[3] ), .Z(n_17871));
	notech_inv i_28048(.A(busy_ram), .Z(n_17872));
	notech_inv i_28049(.A(\queue_0[87] ), .Z(n_17873));
	notech_inv i_28050(.A(\queue_0[127] ), .Z(n_17874));
	notech_inv i_28051(.A(\queue_0[126] ), .Z(n_17875));
	notech_inv i_28052(.A(\queue_0[125] ), .Z(n_17876));
	notech_inv i_28053(.A(\queue_0[124] ), .Z(n_17877));
	notech_inv i_28054(.A(\queue_0[123] ), .Z(n_17878));
	notech_inv i_28055(.A(\queue_0[122] ), .Z(n_17879));
	notech_inv i_28056(.A(\queue_0[121] ), .Z(n_17880));
	notech_inv i_28057(.A(\queue_0[120] ), .Z(n_17881));
	notech_inv i_28058(.A(\queue_0[119] ), .Z(n_17882));
	notech_inv i_28059(.A(\queue_0[118] ), .Z(n_17883));
	notech_inv i_28060(.A(\queue_0[117] ), .Z(n_17884));
	notech_inv i_28061(.A(\queue_0[116] ), .Z(n_17885));
	notech_inv i_28062(.A(\queue_0[114] ), .Z(n_17886));
	notech_inv i_28063(.A(\queue_0[113] ), .Z(n_17887));
	notech_inv i_28064(.A(\queue_0[112] ), .Z(n_17888));
	notech_inv i_28065(.A(\queue_0[111] ), .Z(n_17889));
	notech_inv i_28066(.A(\queue_0[110] ), .Z(n_17890));
	notech_inv i_28067(.A(\queue_0[109] ), .Z(n_17891));
	notech_inv i_28068(.A(\queue_0[108] ), .Z(n_17892));
	notech_inv i_28069(.A(\queue_0[107] ), .Z(n_17893));
	notech_inv i_28070(.A(\queue_0[106] ), .Z(n_17894));
	notech_inv i_28071(.A(\queue_0[105] ), .Z(n_17895));
	notech_inv i_28072(.A(\queue_0[104] ), .Z(n_17896));
	notech_inv i_28073(.A(\queue_0[103] ), .Z(n_17897));
	notech_inv i_28074(.A(\queue_0[102] ), .Z(n_17898));
	notech_inv i_28075(.A(\queue_0[101] ), .Z(n_17899));
	notech_inv i_28076(.A(\queue_0[100] ), .Z(n_17900));
	notech_inv i_28077(.A(\queue_0[99] ), .Z(n_17901));
	notech_inv i_28078(.A(\queue_0[98] ), .Z(n_17902));
	notech_inv i_28079(.A(\queue_0[97] ), .Z(n_17903));
	notech_inv i_28080(.A(\queue_0[96] ), .Z(n_17904));
	notech_inv i_28081(.A(\queue_0[95] ), .Z(n_17905));
	notech_inv i_28082(.A(\queue_0[94] ), .Z(n_17906));
	notech_inv i_28083(.A(\queue_0[93] ), .Z(n_17907));
	notech_inv i_28084(.A(\queue_0[92] ), .Z(n_17908));
	notech_inv i_28085(.A(\queue_0[91] ), .Z(n_17909));
	notech_inv i_28086(.A(\queue_0[89] ), .Z(n_17910));
	notech_inv i_28087(.A(\queue_0[88] ), .Z(n_17911));
	notech_inv i_28088(.A(\queue_0[86] ), .Z(n_17912));
	notech_inv i_28089(.A(\queue_0[85] ), .Z(n_17913));
	notech_inv i_28090(.A(\queue_0[84] ), .Z(n_17914));
	notech_inv i_28091(.A(\queue_0[83] ), .Z(n_17915));
	notech_inv i_28092(.A(\queue_0[82] ), .Z(n_17916));
	notech_inv i_28093(.A(\queue_0[81] ), .Z(n_17917));
	notech_inv i_28094(.A(\queue_0[80] ), .Z(n_17918));
	notech_inv i_28095(.A(\queue_0[79] ), .Z(n_17919));
	notech_inv i_28096(.A(\queue_0[78] ), .Z(n_17920));
	notech_inv i_28097(.A(\queue_0[77] ), .Z(n_17921));
	notech_inv i_28098(.A(\queue_0[76] ), .Z(n_17922));
	notech_inv i_28099(.A(\queue_0[75] ), .Z(n_17923));
	notech_inv i_28100(.A(\queue_0[74] ), .Z(n_17924));
	notech_inv i_28101(.A(\queue_0[73] ), .Z(n_17925));
	notech_inv i_28102(.A(\queue_0[72] ), .Z(n_17926));
	notech_inv i_28103(.A(\queue_0[71] ), .Z(n_17927));
	notech_inv i_28104(.A(\queue_0[70] ), .Z(n_17928));
	notech_inv i_28105(.A(\queue_0[69] ), .Z(n_17929));
	notech_inv i_28106(.A(\queue_0[68] ), .Z(n_17930));
	notech_inv i_28107(.A(\queue_0[67] ), .Z(n_17931));
	notech_inv i_28108(.A(\queue_0[66] ), .Z(n_17932));
	notech_inv i_28109(.A(\queue_0[65] ), .Z(n_17933));
	notech_inv i_28110(.A(\queue_0[64] ), .Z(n_17934));
	notech_inv i_28111(.A(\queue_0[63] ), .Z(n_17935));
	notech_inv i_28112(.A(\queue_0[62] ), .Z(n_17936));
	notech_inv i_28113(.A(\queue_0[61] ), .Z(n_17937));
	notech_inv i_28114(.A(\queue_0[60] ), .Z(n_17938));
	notech_inv i_28115(.A(\queue_0[59] ), .Z(n_17939));
	notech_inv i_28116(.A(\queue_0[58] ), .Z(n_17940));
	notech_inv i_28117(.A(\queue_0[57] ), .Z(n_17941));
	notech_inv i_28118(.A(\queue_0[56] ), .Z(n_17942));
	notech_inv i_28119(.A(\queue_0[55] ), .Z(n_17943));
	notech_inv i_28120(.A(\queue_0[54] ), .Z(n_17944));
	notech_inv i_28121(.A(\queue_0[53] ), .Z(n_17945));
	notech_inv i_28122(.A(\queue_0[52] ), .Z(n_17946));
	notech_inv i_28123(.A(\queue_0[51] ), .Z(n_17947));
	notech_inv i_28124(.A(\queue_0[50] ), .Z(n_17948));
	notech_inv i_28125(.A(\queue_0[49] ), .Z(n_17949));
	notech_inv i_28126(.A(\queue_0[48] ), .Z(n_17950));
	notech_inv i_28127(.A(\queue_0[47] ), .Z(n_17951));
	notech_inv i_28128(.A(\queue_0[46] ), .Z(n_17952));
	notech_inv i_28129(.A(\queue_0[45] ), .Z(n_17953));
	notech_inv i_28130(.A(\queue_0[44] ), .Z(n_17954));
	notech_inv i_28131(.A(\queue_0[43] ), .Z(n_17955));
	notech_inv i_28132(.A(\queue_0[42] ), .Z(n_17956));
	notech_inv i_28133(.A(\queue_0[41] ), .Z(n_17957));
	notech_inv i_28134(.A(\queue_0[40] ), .Z(n_17958));
	notech_inv i_28135(.A(\queue_0[39] ), .Z(n_17959));
	notech_inv i_28136(.A(\queue_0[38] ), .Z(n_17960));
	notech_inv i_28137(.A(\queue_0[37] ), .Z(n_17961));
	notech_inv i_28138(.A(\queue_0[36] ), .Z(n_17962));
	notech_inv i_28139(.A(\queue_0[35] ), .Z(n_17963));
	notech_inv i_28140(.A(\queue_0[34] ), .Z(n_17964));
	notech_inv i_28141(.A(\queue_0[33] ), .Z(n_17965));
	notech_inv i_28142(.A(\queue_0[32] ), .Z(n_17966));
	notech_inv i_28143(.A(\queue_0[31] ), .Z(n_17967));
	notech_inv i_28144(.A(\queue_0[30] ), .Z(n_17968));
	notech_inv i_28145(.A(\queue_0[29] ), .Z(n_17969));
	notech_inv i_28146(.A(\queue_0[28] ), .Z(n_17970));
	notech_inv i_28147(.A(\queue_0[26] ), .Z(n_17971));
	notech_inv i_28148(.A(\queue_0[25] ), .Z(n_17972));
	notech_inv i_28149(.A(\queue_0[24] ), .Z(n_17973));
	notech_inv i_28150(.A(\queue_0[23] ), .Z(n_17974));
	notech_inv i_28151(.A(\queue_0[22] ), .Z(n_17975));
	notech_inv i_28152(.A(\queue_0[21] ), .Z(n_17976));
	notech_inv i_28153(.A(\queue_0[20] ), .Z(n_17977));
	notech_inv i_28154(.A(\queue_0[17] ), .Z(n_17978));
	notech_inv i_28155(.A(\queue_0[16] ), .Z(n_17979));
	notech_inv i_28156(.A(\queue_0[15] ), .Z(n_17980));
	notech_inv i_28157(.A(\queue_0[14] ), .Z(n_17981));
	notech_inv i_28158(.A(\queue_0[10] ), .Z(n_17982));
	notech_inv i_28159(.A(\queue_0[9] ), .Z(n_17983));
	notech_inv i_28160(.A(\queue_0[8] ), .Z(n_17984));
	notech_inv i_28161(.A(\queue_0[7] ), .Z(n_17985));
	notech_inv i_28162(.A(\queue_0[6] ), .Z(n_17986));
	notech_inv i_28163(.A(\queue_0[5] ), .Z(n_17987));
	notech_inv i_28164(.A(\queue_0[4] ), .Z(n_17988));
	notech_inv i_28165(.A(\queue_0[1] ), .Z(n_17989));
	notech_inv i_28166(.A(\queue_0[0] ), .Z(n_17990));
	notech_inv i_28167(.A(n_61563), .Z(n_17991));
	notech_inv i_28168(.A(\queue_0[2] ), .Z(n_17992));
	notech_inv i_28169(.A(\queue_0[12] ), .Z(n_17993));
	notech_inv i_28170(.A(\queue_0[13] ), .Z(n_17994));
	notech_inv i_28171(.A(\queue_0[18] ), .Z(n_17995));
	notech_inv i_28172(.A(\queue_0[115] ), .Z(n_17996));
	notech_inv i_28173(.A(\queue_0[90] ), .Z(n_17997));
	AWDP_EQ_228374 i_64346(.O0({n_36941}), .tagA(tagA), .addr({iaddr[31], iaddr
		[30], iaddr[29], iaddr[28], iaddr[27], iaddr[26], iaddr[25], iaddr
		[24], iaddr[23], iaddr[22], iaddr[21], iaddr[20], iaddr[19], iaddr
		[18], iaddr[17], iaddr[16], iaddr[15], iaddr[14]}));
	AWDP_EQ_328640 i_64338(.O0({n_34592}), .addr(iaddr), .addrf(addrf));
	AWDP_ADD_27 i_64328(.O0(nbus_12105), .addrshft(addrshft), .useq_ptr(useq_ptr
		));
	AWDP_INC_10 i_64313(.O0({n_34620, n_34618, n_34616, n_34614, n_34612, n_34610
		, n_34608, n_34606, n_34604, n_34602, n_34600}), .purge_cnt(purge_cnt
		));
	datacache c1(.clk(clk), .A(cacheA), .D({AMBIT_GND, cacheD[148], 
		AMBIT_GND, AMBIT_GND, cacheD[145], cacheD[144], cacheD[143], cacheD
		[142], cacheD[141], cacheD[140], cacheD[139], cacheD[138], cacheD
		[137], cacheD[136], cacheD[135], cacheD[134], cacheD[133], cacheD
		[132], cacheD[131], cacheD[130], cacheD[129], cacheD[128], cacheD
		[127], cacheD[126], cacheD[125], cacheD[124], cacheD[123], cacheD
		[122], cacheD[121], cacheD[120], cacheD[119], cacheD[118], cacheD
		[117], cacheD[116], cacheD[115], cacheD[114], cacheD[113], cacheD
		[112], cacheD[111], cacheD[110], cacheD[109], cacheD[108], cacheD
		[107], cacheD[106], cacheD[105], cacheD[104], cacheD[103], cacheD
		[102], cacheD[101], cacheD[100], cacheD[99], cacheD[98], cacheD[
		97], cacheD[96], cacheD[95], cacheD[94], cacheD[93], cacheD[92],
		 cacheD[91], cacheD[90], cacheD[89], cacheD[88], cacheD[87], cacheD
		[86], cacheD[85], cacheD[84], cacheD[83], cacheD[82], cacheD[81]
		, cacheD[80], cacheD[79], cacheD[78], cacheD[77], cacheD[76], cacheD
		[75], cacheD[74], cacheD[73], cacheD[72], cacheD[71], cacheD[70]
		, cacheD[69], cacheD[68], cacheD[67], cacheD[66], cacheD[65], cacheD
		[64], cacheD[63], cacheD[62], cacheD[61], cacheD[60], cacheD[59]
		, cacheD[58], cacheD[57], cacheD[56], cacheD[55], cacheD[54], cacheD
		[53], cacheD[52], cacheD[51], cacheD[50], cacheD[49], cacheD[48]
		, cacheD[47], cacheD[46], cacheD[45], cacheD[44], cacheD[43], cacheD
		[42], cacheD[41], cacheD[40], cacheD[39], cacheD[38], cacheD[37]
		, cacheD[36], cacheD[35], cacheD[34], cacheD[33], cacheD[32], cacheD
		[31], cacheD[30], cacheD[29], cacheD[28], cacheD[27], cacheD[26]
		, cacheD[25], cacheD[24], cacheD[23], cacheD[22], cacheD[21], cacheD
		[20], cacheD[19], cacheD[18], cacheD[17], cacheD[16], cacheD[15]
		, cacheD[14], cacheD[13], cacheD[12], cacheD[11], cacheD[10], cacheD
		[9], cacheD[8], cacheD[7], cacheD[6], cacheD[5], cacheD[4], cacheD
		[3], cacheD[2], cacheD[1], cacheD[0]}), .Q({tagV[3], tagV[2], tagV
		[1], tagV[0], tagA[17], tagA[16], tagA[15], tagA[14], tagA[13], tagA
		[12], tagA[11], tagA[10], tagA[9], tagA[8], tagA[7], tagA[6], tagA
		[5], tagA[4], tagA[3], tagA[2], tagA[1], tagA[0], \queue_0[127] 
		, \queue_0[126] , \queue_0[125] , \queue_0[124] , \queue_0[123] 
		, \queue_0[122] , \queue_0[121] , \queue_0[120] , \queue_0[119] 
		, \queue_0[118] , \queue_0[117] , \queue_0[116] , \queue_0[115] 
		, \queue_0[114] , \queue_0[113] , \queue_0[112] , \queue_0[111] 
		, \queue_0[110] , \queue_0[109] , \queue_0[108] , \queue_0[107] 
		, \queue_0[106] , \queue_0[105] , \queue_0[104] , \queue_0[103] 
		, \queue_0[102] , \queue_0[101] , \queue_0[100] , \queue_0[99] ,
		 \queue_0[98] , \queue_0[97] , \queue_0[96] , \queue_0[95] , \queue_0[94] 
		, \queue_0[93] , \queue_0[92] , \queue_0[91] , \queue_0[90] , \queue_0[89] 
		, \queue_0[88] , \queue_0[87] , \queue_0[86] , \queue_0[85] , \queue_0[84] 
		, \queue_0[83] , \queue_0[82] , \queue_0[81] , \queue_0[80] , \queue_0[79] 
		, \queue_0[78] , \queue_0[77] , \queue_0[76] , \queue_0[75] , \queue_0[74] 
		, \queue_0[73] , \queue_0[72] , \queue_0[71] , \queue_0[70] , \queue_0[69] 
		, \queue_0[68] , \queue_0[67] , \queue_0[66] , \queue_0[65] , \queue_0[64] 
		, \queue_0[63] , \queue_0[62] , \queue_0[61] , \queue_0[60] , \queue_0[59] 
		, \queue_0[58] , \queue_0[57] , \queue_0[56] , \queue_0[55] , \queue_0[54] 
		, \queue_0[53] , \queue_0[52] , \queue_0[51] , \queue_0[50] , \queue_0[49] 
		, \queue_0[48] , \queue_0[47] , \queue_0[46] , \queue_0[45] , \queue_0[44] 
		, \queue_0[43] , \queue_0[42] , \queue_0[41] , \queue_0[40] , \queue_0[39] 
		, \queue_0[38] , \queue_0[37] , \queue_0[36] , \queue_0[35] , \queue_0[34] 
		, \queue_0[33] , \queue_0[32] , \queue_0[31] , \queue_0[30] , \queue_0[29] 
		, \queue_0[28] , \queue_0[27] , \queue_0[26] , \queue_0[25] , \queue_0[24] 
		, \queue_0[23] , \queue_0[22] , \queue_0[21] , \queue_0[20] , \queue_0[19] 
		, \queue_0[18] , \queue_0[17] , \queue_0[16] , \queue_0[15] , \queue_0[14] 
		, \queue_0[13] , \queue_0[12] , \queue_0[11] , \queue_0[10] , \queue_0[9] 
		, \queue_0[8] , \queue_0[7] , \queue_0[6] , \queue_0[5] , \queue_0[4] 
		, \queue_0[3] , \queue_0[2] , \queue_0[1] , \queue_0[0] }), .WEN
		(codeWEN), .M({AMBIT_VDD, AMBIT_VDD, AMBIT_VDD, AMBIT_VDD, 
		AMBIT_VDD, AMBIT_VDD, AMBIT_VDD, AMBIT_VDD, AMBIT_VDD, AMBIT_VDD
		, AMBIT_VDD, AMBIT_VDD, AMBIT_VDD, AMBIT_VDD, AMBIT_VDD, 
		AMBIT_VDD}));
	AWDP_ADD_9 i_64305(.O0(addr_0), .addr(iaddr));
endmodule
module core(clk, rstn, ivect, int_main, iack, code_addr, code_data, code_req, code_ack
		, code_wreq, code_wack, code_wdata, readio_data, io_add, writeio_data
		, writeio_req, readio_req, writeio_ack, readio_ack, write_req, write_ack
		, write_data, write_sz, read_sz, write_msk, read_req, read_ack, read_data
		, Daddr, busy_ram, ipg_fault, outstanding);

	input clk;
	input rstn;
	input [7:0] ivect;
	input int_main;
	output iack;
	output [31:0] code_addr;
	input [127:0] code_data;
	output code_req;
	input code_ack;
	output code_wreq;
	input code_wack;
	output [31:0] code_wdata;
	input [31:0] readio_data;
	output [31:0] io_add;
	output [31:0] writeio_data;
	output writeio_req;
	output readio_req;
	input writeio_ack;
	input readio_ack;
	output write_req;
	input write_ack;
	output [31:0] write_data;
	output [1:0] write_sz;
	output [1:0] read_sz;
	output [3:0] write_msk;
	output read_req;
	input read_ack;
	input [31:0] read_data;
	output [31:0] Daddr;
	input busy_ram;
	output ipg_fault;
	output outstanding;

	wire [31:0] pc_out;
	wire [3:0] useq_ptr;
	wire [5:0] valid_len;
	wire [31:0] icr2;
	wire [31:0] cr2;
	wire [127:0] queue;
	wire [1:0] int_write_sz;
	wire [31:0] int_Daddr;
	wire [31:0] iwrite_data;
	wire [31:0] int_code_addr;
	wire [31:0] write_data_realign;
	wire [1:0] nbus_14544;
	wire [31:0] Daddr_realign;
	wire [31:0] read_data_realign;



	Dtlb i_Dtlb(.clk(clk), .rstn(rstn), .addr_phys(Daddr_realign), .cr3({\cr3[31] 
		, \cr3[30] , \cr3[29] , \cr3[28] , \cr3[27] , \cr3[26] , \cr3[25] 
		, \cr3[24] , \cr3[23] , \cr3[22] , \cr3[21] , \cr3[20] , \cr3[19] 
		, \cr3[18] , \cr3[17] , \cr3[16] , \cr3[15] , \cr3[14] , \cr3[13] 
		, \cr3[12] , UNCONNECTED_000, UNCONNECTED_001, UNCONNECTED_002, 
		UNCONNECTED_003, UNCONNECTED_004, UNCONNECTED_005, 
		UNCONNECTED_006, UNCONNECTED_007, UNCONNECTED_008, 
		UNCONNECTED_009, UNCONNECTED_010, UNCONNECTED_011}), .cr0({
		UNCONNECTED_012, UNCONNECTED_013, UNCONNECTED_014, 
		UNCONNECTED_015, UNCONNECTED_016, UNCONNECTED_017, 
		UNCONNECTED_018, UNCONNECTED_019, UNCONNECTED_020, 
		UNCONNECTED_021, UNCONNECTED_022, UNCONNECTED_023, 
		UNCONNECTED_024, UNCONNECTED_025, UNCONNECTED_026, \cr0[16] , 
		UNCONNECTED_027, UNCONNECTED_028, UNCONNECTED_029, 
		UNCONNECTED_030, UNCONNECTED_031, UNCONNECTED_032, 
		UNCONNECTED_033, UNCONNECTED_034, UNCONNECTED_035, 
		UNCONNECTED_036, UNCONNECTED_037, UNCONNECTED_038, 
		UNCONNECTED_039, UNCONNECTED_040, UNCONNECTED_041, 
		UNCONNECTED_042}), .data_miss(read_data_realign), .iDaddr(int_Daddr
		), .pg_en(pg_en), .iwrite_data(iwrite_data), .owrite_data(write_data_realign
		), .iread_req(int_read_req), .iread_ack(read_ack_realign), .iwrite_req
		(int_write_req), .iwrite_ack(write_ack_realign), .iwrite_sz(int_write_sz
		), .owrite_sz(nbus_14544), .oread_req(read_req_realign), .oread_ack
		(int_read_ack), .owrite_req(write_req_realign), .owrite_ack(int_write_ack
		), .pg_fault(pg_fault), .wr_fault(wr_fault), .cr2(cr2), .flush_tlb
		(flush_Dtlb), .cs({UNCONNECTED_043, UNCONNECTED_044, 
		UNCONNECTED_045, UNCONNECTED_046, UNCONNECTED_047, 
		UNCONNECTED_048, UNCONNECTED_049, UNCONNECTED_050, 
		UNCONNECTED_051, UNCONNECTED_052, UNCONNECTED_053, 
		UNCONNECTED_054, UNCONNECTED_055, UNCONNECTED_056, 
		UNCONNECTED_057, UNCONNECTED_058, UNCONNECTED_059, 
		UNCONNECTED_060, UNCONNECTED_061, UNCONNECTED_062, 
		UNCONNECTED_063, UNCONNECTED_064, UNCONNECTED_065, 
		UNCONNECTED_066, UNCONNECTED_067, UNCONNECTED_068, 
		UNCONNECTED_069, UNCONNECTED_070, UNCONNECTED_071, 
		UNCONNECTED_072, \cs[1] , \cs[0] }), .pt_fault(pt_fault), .busy_ram
		(busy_ram));
	realign i_realign(.clk(clk), .rstn(rstn), .write_msk_out(write_msk), .addr_in
		(Daddr_realign), .addr_out({Daddr[31], Daddr[30], Daddr[29], Daddr
		[28], Daddr[27], Daddr[26], Daddr[25], Daddr[24], Daddr[23], Daddr
		[22], Daddr[21], Daddr[20], Daddr[19], Daddr[18], Daddr[17], Daddr
		[16], Daddr[15], Daddr[14], Daddr[13], Daddr[12], Daddr[11], Daddr
		[10], Daddr[9], Daddr[8], Daddr[7], Daddr[6], Daddr[5], Daddr[4]
		, Daddr[3], Daddr[2], UNCONNECTED_073, UNCONNECTED_074}), .write_sz_in
		(nbus_14544), .write_req_in(write_req_realign), .write_req_out(write_req
		), .write_ack_in(write_ack), .write_ack_out(write_ack_realign), 
		.read_req_in(read_req_realign), .read_req_out(read_req), .read_ack_in
		(read_ack), .read_ack_out(read_ack_realign), .read_data_in(read_data
		), .read_data_out(read_data_realign), .write_data_in(write_data_realign
		), .write_data_out(write_data));
	Itlb i_Itlb(.clk(clk), .rstn(rstn), .addr_phys({code_addr[31], code_addr
		[30], code_addr[29], code_addr[28], code_addr[27], code_addr[26]
		, code_addr[25], code_addr[24], code_addr[23], code_addr[22], code_addr
		[21], code_addr[20], code_addr[19], code_addr[18], code_addr[17]
		, code_addr[16], code_addr[15], code_addr[14], code_addr[13], code_addr
		[12], code_addr[11], code_addr[10], code_addr[9], code_addr[8], code_addr
		[7], code_addr[6], code_addr[5], code_addr[4], code_addr[3], code_addr
		[2], UNCONNECTED_075, UNCONNECTED_076}), .cr3({\cr3[31] , \cr3[30] 
		, \cr3[29] , \cr3[28] , \cr3[27] , \cr3[26] , \cr3[25] , \cr3[24] 
		, \cr3[23] , \cr3[22] , \cr3[21] , \cr3[20] , \cr3[19] , \cr3[18] 
		, \cr3[17] , \cr3[16] , \cr3[15] , \cr3[14] , \cr3[13] , \cr3[12] 
		, UNCONNECTED_077, UNCONNECTED_078, UNCONNECTED_079, 
		UNCONNECTED_080, UNCONNECTED_081, UNCONNECTED_082, 
		UNCONNECTED_083, UNCONNECTED_084, UNCONNECTED_085, 
		UNCONNECTED_086, UNCONNECTED_087, UNCONNECTED_088}), .data_miss(
		{code_data[31], code_data[30], code_data[29], code_data[28], code_data
		[27], code_data[26], code_data[25], code_data[24], code_data[23]
		, code_data[22], code_data[21], code_data[20], code_data[19], code_data
		[18], code_data[17], code_data[16], code_data[15], code_data[14]
		, code_data[13], code_data[12], UNCONNECTED_089, UNCONNECTED_090
		, UNCONNECTED_091, UNCONNECTED_092, code_data[7], code_data[6], code_data
		[5], code_data[4], code_data[3], code_data[2], code_data[1], code_data
		[0]}), .iDaddr(int_code_addr), .pg_en(pg_en), .owrite_data({
		UNCONNECTED_093, UNCONNECTED_094, UNCONNECTED_095, 
		UNCONNECTED_096, UNCONNECTED_097, UNCONNECTED_098, 
		UNCONNECTED_099, UNCONNECTED_100, UNCONNECTED_101, 
		UNCONNECTED_102, UNCONNECTED_103, UNCONNECTED_104, 
		UNCONNECTED_105, UNCONNECTED_106, UNCONNECTED_107, 
		UNCONNECTED_108, UNCONNECTED_109, UNCONNECTED_110, 
		UNCONNECTED_111, UNCONNECTED_112, UNCONNECTED_113, 
		UNCONNECTED_114, UNCONNECTED_115, UNCONNECTED_116, code_wdata[7]
		, code_wdata[6], code_wdata[5], code_wdata[4], code_wdata[3], code_wdata
		[2], code_wdata[1], code_wdata[0]}), .iread_req(int_code_req), .iread_ack
		(code_ack), .iwrite_ack(code_wack), .oread_req(code_req), .oread_ack
		(int_code_ack), .owrite_req(code_wreq), .pg_fault(n_4695), .cr2(icr2
		), .flush_tlb(flush_Itlb), .busy_ram(busy_ram));
	useq i_useq(.iaddr(int_code_addr), .idata(code_data), .code_req(int_code_req
		), .code_ack(int_code_ack), .clk(clk), .rstn(rstn), .useq_ptr(useq_ptr
		), .squeue(queue), .pc_in(pc_out), .pc_req(pc_req), .pg_fault(n_4695
		), .pc_pg_fault(pc_pg_fault), .valid_len(valid_len), .busy_ram(busy_ram
		));
	cpu i_cpu(.clk(clk), .rstn(rstn), .iack(iack), .int_cpu(int_main), .ivect
		(ivect), .cr0({UNCONNECTED_117, UNCONNECTED_118, UNCONNECTED_119
		, UNCONNECTED_120, UNCONNECTED_121, UNCONNECTED_122, 
		UNCONNECTED_123, UNCONNECTED_124, UNCONNECTED_125, 
		UNCONNECTED_126, UNCONNECTED_127, UNCONNECTED_128, 
		UNCONNECTED_129, UNCONNECTED_130, UNCONNECTED_131, \cr0[16] , 
		UNCONNECTED_132, UNCONNECTED_133, UNCONNECTED_134, 
		UNCONNECTED_135, UNCONNECTED_136, UNCONNECTED_137, 
		UNCONNECTED_138, UNCONNECTED_139, UNCONNECTED_140, 
		UNCONNECTED_141, UNCONNECTED_142, UNCONNECTED_143, 
		UNCONNECTED_144, UNCONNECTED_145, UNCONNECTED_146, 
		UNCONNECTED_147}), .cr2(cr2), .icr2(icr2), .cr3({\cr3[31] , \cr3[30] 
		, \cr3[29] , \cr3[28] , \cr3[27] , \cr3[26] , \cr3[25] , \cr3[24] 
		, \cr3[23] , \cr3[22] , \cr3[21] , \cr3[20] , \cr3[19] , \cr3[18] 
		, \cr3[17] , \cr3[16] , \cr3[15] , \cr3[14] , \cr3[13] , \cr3[12] 
		, UNCONNECTED_148, UNCONNECTED_149, UNCONNECTED_150, 
		UNCONNECTED_151, UNCONNECTED_152, UNCONNECTED_153, 
		UNCONNECTED_154, UNCONNECTED_155, UNCONNECTED_156, 
		UNCONNECTED_157, UNCONNECTED_158, UNCONNECTED_159}), .cs({
		UNCONNECTED_160, UNCONNECTED_161, UNCONNECTED_162, 
		UNCONNECTED_163, UNCONNECTED_164, UNCONNECTED_165, 
		UNCONNECTED_166, UNCONNECTED_167, UNCONNECTED_168, 
		UNCONNECTED_169, UNCONNECTED_170, UNCONNECTED_171, 
		UNCONNECTED_172, UNCONNECTED_173, UNCONNECTED_174, 
		UNCONNECTED_175, UNCONNECTED_176, UNCONNECTED_177, 
		UNCONNECTED_178, UNCONNECTED_179, UNCONNECTED_180, 
		UNCONNECTED_181, UNCONNECTED_182, UNCONNECTED_183, 
		UNCONNECTED_184, UNCONNECTED_185, UNCONNECTED_186, 
		UNCONNECTED_187, UNCONNECTED_188, UNCONNECTED_189, \cs[1] , \cs[0] 
		}), .pg_fault(pg_fault), .ipg_fault(pc_pg_fault), .useq_ptr(useq_ptr
		), .valid_len(valid_len), .queue(queue), .pg_en(pg_en), .pc_out(pc_out
		), .pc_req(pc_req), .read_req(int_read_req), .write_req(int_write_req
		), .read_ack(int_read_ack), .write_ack(int_write_ack), .flush_Itlb
		(flush_Itlb), .flush_Dtlb(flush_Dtlb), .readio_req(readio_req), 
		.writeio_req(writeio_req), .readio_ack(readio_ack), .writeio_ack
		(writeio_ack), .write_data(iwrite_data), .writeio_data(writeio_data
		), .read_data(read_data_realign), .readio_data(readio_data), .write_sz
		(int_write_sz), .io_add({UNCONNECTED_190, UNCONNECTED_191, 
		UNCONNECTED_192, UNCONNECTED_193, UNCONNECTED_194, 
		UNCONNECTED_195, UNCONNECTED_196, UNCONNECTED_197, 
		UNCONNECTED_198, UNCONNECTED_199, UNCONNECTED_200, 
		UNCONNECTED_201, UNCONNECTED_202, UNCONNECTED_203, 
		UNCONNECTED_204, UNCONNECTED_205, io_add[15], io_add[14], io_add
		[13], io_add[12], io_add[11], io_add[10], io_add[9], io_add[8], io_add
		[7], io_add[6], io_add[5], io_add[4], io_add[3], io_add[2], io_add
		[1], io_add[0]}), .Daddr(int_Daddr), .pt_fault(pt_fault), .wr_fault
		(wr_fault));
endmodule
module v586(m00_AXI_RSTN, m00_AXI_CLK, m00_AXI_AWADDR, m00_AXI_AWVALID, m00_AXI_AWREADY
		, m00_AXI_AWBURST, m00_AXI_AWLEN, m00_AXI_AWSIZE, m00_AXI_ARADDR
		, m00_AXI_ARVALID, m00_AXI_ARREADY, m00_AXI_ARBURST, m00_AXI_ARLEN
		, m00_AXI_ARSIZE, m00_AXI_WDATA, m00_AXI_WVALID, m00_AXI_WREADY,
		 m00_AXI_WSTRB, m00_AXI_WLAST, m00_AXI_RDATA, m00_AXI_RVALID, m00_AXI_RREADY
		, m00_AXI_RLAST, m00_AXI_BVALID, m00_AXI_BREADY, m01_AXI_AWADDR,
		 m01_AXI_AWVALID, m01_AXI_AWREADY, m01_AXI_AWBURST, m01_AXI_AWLEN
		, m01_AXI_AWSIZE, m01_AXI_ARADDR, m01_AXI_ARVALID, m01_AXI_ARREADY
		, m01_AXI_ARBURST, m01_AXI_ARLEN, m01_AXI_ARSIZE, m01_AXI_WDATA,
		 m01_AXI_WVALID, m01_AXI_WREADY, m01_AXI_WSTRB, m01_AXI_WLAST, m01_AXI_RDATA
		, m01_AXI_RVALID, m01_AXI_RREADY, m01_AXI_RLAST, m01_AXI_BVALID,
		 m01_AXI_BREADY, int_pic, iack, ivect, debug);

	input m00_AXI_RSTN;
	input m00_AXI_CLK;
	output [31:0] m00_AXI_AWADDR;
	output m00_AXI_AWVALID;
	input m00_AXI_AWREADY;
	output [1:0] m00_AXI_AWBURST;
	output [7:0] m00_AXI_AWLEN;
	output [2:0] m00_AXI_AWSIZE;
	output [31:0] m00_AXI_ARADDR;
	output m00_AXI_ARVALID;
	input m00_AXI_ARREADY;
	output [1:0] m00_AXI_ARBURST;
	output [7:0] m00_AXI_ARLEN;
	output [2:0] m00_AXI_ARSIZE;
	output [31:0] m00_AXI_WDATA;
	output m00_AXI_WVALID;
	input m00_AXI_WREADY;
	output [3:0] m00_AXI_WSTRB;
	output m00_AXI_WLAST;
	input [31:0] m00_AXI_RDATA;
	input m00_AXI_RVALID;
	output m00_AXI_RREADY;
	input m00_AXI_RLAST;
	input m00_AXI_BVALID;
	output m00_AXI_BREADY;
	output [31:0] m01_AXI_AWADDR;
	output m01_AXI_AWVALID;
	input m01_AXI_AWREADY;
	output [1:0] m01_AXI_AWBURST;
	output [7:0] m01_AXI_AWLEN;
	output [2:0] m01_AXI_AWSIZE;
	output [31:0] m01_AXI_ARADDR;
	output m01_AXI_ARVALID;
	input m01_AXI_ARREADY;
	output [1:0] m01_AXI_ARBURST;
	output [7:0] m01_AXI_ARLEN;
	output [2:0] m01_AXI_ARSIZE;
	output [31:0] m01_AXI_WDATA;
	output m01_AXI_WVALID;
	input m01_AXI_WREADY;
	output [3:0] m01_AXI_WSTRB;
	output m01_AXI_WLAST;
	input [31:0] m01_AXI_RDATA;
	input m01_AXI_RVALID;
	output m01_AXI_RREADY;
	input m01_AXI_RLAST;
	input m01_AXI_BVALID;
	output m01_AXI_BREADY;
	input int_pic;
	output iack;
	input [7:0] ivect;
	output [4:0] debug;

	wire [3:0] write_msk;
	wire [31:0] writeio_data;
	wire [31:0] readio_data;
	wire [31:0] read_data;
	wire [31:0] write_data;
	wire [127:0] code_data;

	assign m00_AXI_BREADY = 1'b1;
	assign m01_AXI_AWBURST[1] = 1'b0;
	assign m01_AXI_AWBURST[0] = 1'b1;
	assign m01_AXI_AWLEN[7] = 1'b0;
	assign m01_AXI_AWLEN[6] = 1'b0;
	assign m01_AXI_AWLEN[5] = 1'b0;
	assign m01_AXI_AWLEN[4] = 1'b0;
	assign m01_AXI_AWLEN[3] = 1'b0;
	assign m01_AXI_AWLEN[2] = 1'b0;
	assign m01_AXI_AWLEN[1] = 1'b0;
	assign m01_AXI_AWLEN[0] = 1'b0;
	assign m01_AXI_AWSIZE[2] = 1'b0;
	assign m01_AXI_AWSIZE[1] = 1'b1;
	assign m01_AXI_AWSIZE[0] = 1'b0;
	assign m01_AXI_ARBURST[1] = 1'b0;
	assign m01_AXI_ARBURST[0] = 1'b1;
	assign m01_AXI_ARLEN[7] = 1'b0;
	assign m01_AXI_ARLEN[6] = 1'b0;
	assign m01_AXI_ARLEN[5] = 1'b0;
	assign m01_AXI_ARLEN[4] = 1'b0;
	assign m01_AXI_ARLEN[3] = 1'b0;
	assign m01_AXI_ARLEN[2] = 1'b0;
	assign m01_AXI_ARLEN[1] = 1'b0;
	assign m01_AXI_ARLEN[0] = 1'b0;
	assign m01_AXI_ARSIZE[2] = 1'b0;
	assign m01_AXI_ARSIZE[1] = 1'b1;
	assign m01_AXI_ARSIZE[0] = 1'b0;
	assign m01_AXI_WSTRB[3] = 1'b0;
	assign m01_AXI_WSTRB[2] = 1'b0;
	assign m01_AXI_WSTRB[1] = 1'b0;
	assign m01_AXI_WSTRB[0] = 1'b1;


	notech_inv i_15112(.A(n_63278), .Z(n_63280));
	notech_inv i_15111(.A(n_63278), .Z(n_63279));
	notech_inv i_15110(.A(m00_AXI_CLK), .Z(n_63278));
	biu32_axi ubiu(.rstn(m00_AXI_RSTN), .clk(n_63279), .write_req(write_req)
		, .write_ack(write_ack), .write_data(write_data), .write_msk(write_msk
		), .read_req(read_req), .read_ack(read_ack), .read_data(read_data
		), .Daddr({\Daddr[31] , \Daddr[30] , \Daddr[29] , \Daddr[28] , \Daddr[27] 
		, \Daddr[26] , \Daddr[25] , \Daddr[24] , \Daddr[23] , \Daddr[22] 
		, \Daddr[21] , \Daddr[20] , \Daddr[19] , \Daddr[18] , \Daddr[17] 
		, \Daddr[16] , \Daddr[15] , \Daddr[14] , \Daddr[13] , \Daddr[12] 
		, \Daddr[11] , \Daddr[10] , \Daddr[9] , \Daddr[8] , \Daddr[7] , \Daddr[6] 
		, \Daddr[5] , \Daddr[4] , \Daddr[3] , \Daddr[2] , 
		UNCONNECTED_000, UNCONNECTED_001}), .code_req(code_req), .code_ack
		(code_ack), .code_data(code_data), .code_addr({\code_addr[31] , \code_addr[30] 
		, \code_addr[29] , \code_addr[28] , \code_addr[27] , \code_addr[26] 
		, \code_addr[25] , \code_addr[24] , \code_addr[23] , \code_addr[22] 
		, \code_addr[21] , \code_addr[20] , \code_addr[19] , \code_addr[18] 
		, \code_addr[17] , \code_addr[16] , \code_addr[15] , \code_addr[14] 
		, \code_addr[13] , \code_addr[12] , \code_addr[11] , \code_addr[10] 
		, \code_addr[9] , \code_addr[8] , \code_addr[7] , \code_addr[6] 
		, \code_addr[5] , \code_addr[4] , \code_addr[3] , \code_addr[2] 
		, UNCONNECTED_002, UNCONNECTED_003}), .code_wreq(code_wreq), .code_wack
		(code_wack), .code_wdata({UNCONNECTED_004, UNCONNECTED_005, 
		UNCONNECTED_006, UNCONNECTED_007, UNCONNECTED_008, 
		UNCONNECTED_009, UNCONNECTED_010, UNCONNECTED_011, 
		UNCONNECTED_012, UNCONNECTED_013, UNCONNECTED_014, 
		UNCONNECTED_015, UNCONNECTED_016, UNCONNECTED_017, 
		UNCONNECTED_018, UNCONNECTED_019, UNCONNECTED_020, 
		UNCONNECTED_021, UNCONNECTED_022, UNCONNECTED_023, 
		UNCONNECTED_024, UNCONNECTED_025, UNCONNECTED_026, 
		UNCONNECTED_027, \code_wdata[7] , \code_wdata[6] , \code_wdata[5] 
		, \code_wdata[4] , \code_wdata[3] , \code_wdata[2] , \code_wdata[1] 
		, \code_wdata[0] }), .readio_req(readio_req), .writeio_req(writeio_req
		), .readio_ack(readio_ack), .writeio_ack(writeio_ack), .writeio_data
		(writeio_data), .readio_data(readio_data), .io_add({
		UNCONNECTED_028, UNCONNECTED_029, UNCONNECTED_030, 
		UNCONNECTED_031, UNCONNECTED_032, UNCONNECTED_033, 
		UNCONNECTED_034, UNCONNECTED_035, UNCONNECTED_036, 
		UNCONNECTED_037, UNCONNECTED_038, UNCONNECTED_039, 
		UNCONNECTED_040, UNCONNECTED_041, UNCONNECTED_042, 
		UNCONNECTED_043, \io_add[15] , \io_add[14] , \io_add[13] , \io_add[12] 
		, \io_add[11] , \io_add[10] , \io_add[9] , \io_add[8] , \io_add[7] 
		, \io_add[6] , \io_add[5] , \io_add[4] , \io_add[3] , \io_add[2] 
		, \io_add[1] , \io_add[0] }), .axi_AW(m00_AXI_AWADDR), .axi_AWVALID
		(m00_AXI_AWVALID), .axi_AWREADY(m00_AXI_AWREADY), .axi_AWBURST(m00_AXI_AWBURST
		), .axi_AWLEN(m00_AXI_AWLEN), .axi_AWSIZE(m00_AXI_AWSIZE), .axi_W
		(m00_AXI_WDATA), .axi_WVALID(m00_AXI_WVALID), .axi_WREADY(m00_AXI_WREADY
		), .axi_WSTRB(m00_AXI_WSTRB), .axi_WLAST(m00_AXI_WLAST), .axi_AR
		(m00_AXI_ARADDR), .axi_ARVALID(m00_AXI_ARVALID), .axi_ARREADY(m00_AXI_ARREADY
		), .axi_ARBURST(m00_AXI_ARBURST), .axi_ARLEN(m00_AXI_ARLEN), .axi_ARSIZE
		(m00_AXI_ARSIZE), .axi_R(m00_AXI_RDATA), .axi_RVALID(m00_AXI_RVALID
		), .axi_RREADY(m00_AXI_RREADY), .axi_RLAST(m00_AXI_RLAST), .axi_io_AW
		(m01_AXI_AWADDR), .axi_io_AWVALID(m01_AXI_AWVALID), .axi_io_AWREADY
		(m01_AXI_AWREADY), .axi_io_W(m01_AXI_WDATA), .axi_io_WVALID(m01_AXI_WVALID
		), .axi_io_WREADY(m01_AXI_WREADY), .axi_io_WLAST(m01_AXI_WLAST),
		 .axi_io_AR(m01_AXI_ARADDR), .axi_io_ARVALID(m01_AXI_ARVALID), .axi_io_ARREADY
		(m01_AXI_ARREADY), .axi_io_R(m01_AXI_RDATA), .axi_io_RVALID(m01_AXI_RVALID
		), .axi_io_RREADY(m01_AXI_RREADY), .busy(busy_ram));
	core ucore(.clk(n_63280), .rstn(m00_AXI_RSTN), .ivect(ivect), .int_main(int_pic
		), .iack(iack), .code_addr({\code_addr[31] , \code_addr[30] , \code_addr[29] 
		, \code_addr[28] , \code_addr[27] , \code_addr[26] , \code_addr[25] 
		, \code_addr[24] , \code_addr[23] , \code_addr[22] , \code_addr[21] 
		, \code_addr[20] , \code_addr[19] , \code_addr[18] , \code_addr[17] 
		, \code_addr[16] , \code_addr[15] , \code_addr[14] , \code_addr[13] 
		, \code_addr[12] , \code_addr[11] , \code_addr[10] , \code_addr[9] 
		, \code_addr[8] , \code_addr[7] , \code_addr[6] , \code_addr[5] 
		, \code_addr[4] , \code_addr[3] , \code_addr[2] , 
		UNCONNECTED_044, UNCONNECTED_045}), .code_data(code_data), .code_req
		(code_req), .code_ack(code_ack), .code_wreq(code_wreq), .code_wack
		(code_wack), .code_wdata({UNCONNECTED_046, UNCONNECTED_047, 
		UNCONNECTED_048, UNCONNECTED_049, UNCONNECTED_050, 
		UNCONNECTED_051, UNCONNECTED_052, UNCONNECTED_053, 
		UNCONNECTED_054, UNCONNECTED_055, UNCONNECTED_056, 
		UNCONNECTED_057, UNCONNECTED_058, UNCONNECTED_059, 
		UNCONNECTED_060, UNCONNECTED_061, UNCONNECTED_062, 
		UNCONNECTED_063, UNCONNECTED_064, UNCONNECTED_065, 
		UNCONNECTED_066, UNCONNECTED_067, UNCONNECTED_068, 
		UNCONNECTED_069, \code_wdata[7] , \code_wdata[6] , \code_wdata[5] 
		, \code_wdata[4] , \code_wdata[3] , \code_wdata[2] , \code_wdata[1] 
		, \code_wdata[0] }), .readio_data(readio_data), .io_add({
		UNCONNECTED_070, UNCONNECTED_071, UNCONNECTED_072, 
		UNCONNECTED_073, UNCONNECTED_074, UNCONNECTED_075, 
		UNCONNECTED_076, UNCONNECTED_077, UNCONNECTED_078, 
		UNCONNECTED_079, UNCONNECTED_080, UNCONNECTED_081, 
		UNCONNECTED_082, UNCONNECTED_083, UNCONNECTED_084, 
		UNCONNECTED_085, \io_add[15] , \io_add[14] , \io_add[13] , \io_add[12] 
		, \io_add[11] , \io_add[10] , \io_add[9] , \io_add[8] , \io_add[7] 
		, \io_add[6] , \io_add[5] , \io_add[4] , \io_add[3] , \io_add[2] 
		, \io_add[1] , \io_add[0] }), .writeio_data(writeio_data), .writeio_req
		(writeio_req), .readio_req(readio_req), .writeio_ack(writeio_ack
		), .readio_ack(readio_ack), .write_req(write_req), .write_ack(write_ack
		), .write_data(write_data), .write_msk(write_msk), .read_req(read_req
		), .read_ack(read_ack), .read_data(read_data), .Daddr({\Daddr[31] 
		, \Daddr[30] , \Daddr[29] , \Daddr[28] , \Daddr[27] , \Daddr[26] 
		, \Daddr[25] , \Daddr[24] , \Daddr[23] , \Daddr[22] , \Daddr[21] 
		, \Daddr[20] , \Daddr[19] , \Daddr[18] , \Daddr[17] , \Daddr[16] 
		, \Daddr[15] , \Daddr[14] , \Daddr[13] , \Daddr[12] , \Daddr[11] 
		, \Daddr[10] , \Daddr[9] , \Daddr[8] , \Daddr[7] , \Daddr[6] , \Daddr[5] 
		, \Daddr[4] , \Daddr[3] , \Daddr[2] , UNCONNECTED_086, 
		UNCONNECTED_087}), .busy_ram(busy_ram));
endmodule
